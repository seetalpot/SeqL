
module b17 ( datai_31_, datai_30_, datai_29_, datai_28_, datai_27_, datai_26_,
datai_25_, datai_24_, datai_23_, datai_22_, datai_21_, datai_20_,
datai_19_, datai_18_, datai_17_, datai_16_, datai_15_, datai_14_,
datai_13_, datai_12_, datai_11_, datai_10_, datai_9_, datai_8_,
datai_7_, datai_6_, datai_5_, datai_4_, datai_3_, datai_2_, datai_1_,
datai_0_, hold, na, bs16, ready1, ready2, buf1_reg_0_, buf1_reg_1_,
buf1_reg_2_, buf1_reg_3_, buf1_reg_4_, buf1_reg_5_, buf1_reg_6_,
buf1_reg_7_, buf1_reg_8_, buf1_reg_9_, buf1_reg_10_, buf1_reg_11_,
buf1_reg_12_, buf1_reg_13_, buf1_reg_14_, buf1_reg_15_, buf1_reg_16_,
buf1_reg_17_, buf1_reg_18_, buf1_reg_19_, buf1_reg_20_, buf1_reg_21_,
buf1_reg_22_, buf1_reg_23_, buf1_reg_24_, buf1_reg_25_, buf1_reg_26_,
buf1_reg_27_, buf1_reg_28_, buf1_reg_29_, buf1_reg_30_, buf1_reg_31_,
buf2_reg_0_, buf2_reg_1_, buf2_reg_2_, buf2_reg_3_, buf2_reg_4_,
buf2_reg_5_, buf2_reg_6_, buf2_reg_7_, buf2_reg_8_, buf2_reg_9_,
buf2_reg_10_, buf2_reg_11_, buf2_reg_12_, buf2_reg_13_, buf2_reg_14_,
buf2_reg_15_, buf2_reg_16_, buf2_reg_17_, buf2_reg_18_, buf2_reg_19_,
buf2_reg_20_, buf2_reg_21_, buf2_reg_22_, buf2_reg_23_, buf2_reg_24_,
buf2_reg_25_, buf2_reg_26_, buf2_reg_27_, buf2_reg_28_, buf2_reg_29_,
buf2_reg_30_, buf2_reg_31_, ready12_reg, ready21_reg, ready22_reg,
ready11_reg, p3_be_n_reg_3_, p3_be_n_reg_2_, p3_be_n_reg_1_,
p3_be_n_reg_0_, p3_address_reg_29_, p3_address_reg_28_,
p3_address_reg_27_, p3_address_reg_26_, p3_address_reg_25_,
p3_address_reg_24_, p3_address_reg_23_, p3_address_reg_22_,
p3_address_reg_21_, p3_address_reg_20_, p3_address_reg_19_,
p3_address_reg_18_, p3_address_reg_17_, p3_address_reg_16_,
p3_address_reg_15_, p3_address_reg_14_, p3_address_reg_13_,
p3_address_reg_12_, p3_address_reg_11_, p3_address_reg_10_,
p3_address_reg_9_, p3_address_reg_8_, p3_address_reg_7_,
p3_address_reg_6_, p3_address_reg_5_, p3_address_reg_4_,
p3_address_reg_3_, p3_address_reg_2_, p3_address_reg_1_,
p3_address_reg_0_, p3_state_reg_2_, p3_state_reg_1_, p3_state_reg_0_,
p3_datawidth_reg_0_, p3_datawidth_reg_1_, p3_datawidth_reg_2_,
p3_datawidth_reg_3_, p3_datawidth_reg_4_, p3_datawidth_reg_5_,
p3_datawidth_reg_6_, p3_datawidth_reg_7_, p3_datawidth_reg_8_,
p3_datawidth_reg_9_, p3_datawidth_reg_10_, p3_datawidth_reg_11_,
p3_datawidth_reg_12_, p3_datawidth_reg_13_, p3_datawidth_reg_14_,
p3_datawidth_reg_15_, p3_datawidth_reg_16_, p3_datawidth_reg_17_,
p3_datawidth_reg_18_, p3_datawidth_reg_19_, p3_datawidth_reg_20_,
p3_datawidth_reg_21_, p3_datawidth_reg_22_, p3_datawidth_reg_23_,
p3_datawidth_reg_24_, p3_datawidth_reg_25_, p3_datawidth_reg_26_,
p3_datawidth_reg_27_, p3_datawidth_reg_28_, p3_datawidth_reg_29_,
p3_datawidth_reg_30_, p3_datawidth_reg_31_, p3_state2_reg_3_,
p3_state2_reg_2_, p3_state2_reg_1_, p3_state2_reg_0_,
p3_instqueue_reg_15__7_, p3_instqueue_reg_15__6_,
p3_instqueue_reg_15__5_, p3_instqueue_reg_15__4_,
p3_instqueue_reg_15__3_, p3_instqueue_reg_15__2_,
p3_instqueue_reg_15__1_, p3_instqueue_reg_15__0_,
p3_instqueue_reg_14__7_, p3_instqueue_reg_14__6_,
p3_instqueue_reg_14__5_, p3_instqueue_reg_14__4_,
p3_instqueue_reg_14__3_, p3_instqueue_reg_14__2_,
p3_instqueue_reg_14__1_, p3_instqueue_reg_14__0_,
p3_instqueue_reg_13__7_, p3_instqueue_reg_13__6_,
p3_instqueue_reg_13__5_, p3_instqueue_reg_13__4_,
p3_instqueue_reg_13__3_, p3_instqueue_reg_13__2_,
p3_instqueue_reg_13__1_, p3_instqueue_reg_13__0_,
p3_instqueue_reg_12__7_, p3_instqueue_reg_12__6_,
p3_instqueue_reg_12__5_, p3_instqueue_reg_12__4_,
p3_instqueue_reg_12__3_, p3_instqueue_reg_12__2_,
p3_instqueue_reg_12__1_, p3_instqueue_reg_12__0_,
p3_instqueue_reg_11__7_, p3_instqueue_reg_11__6_,
p3_instqueue_reg_11__5_, p3_instqueue_reg_11__4_,
p3_instqueue_reg_11__3_, p3_instqueue_reg_11__2_,
p3_instqueue_reg_11__1_, p3_instqueue_reg_11__0_,
p3_instqueue_reg_10__7_, p3_instqueue_reg_10__6_,
p3_instqueue_reg_10__5_, p3_instqueue_reg_10__4_,
p3_instqueue_reg_10__3_, p3_instqueue_reg_10__2_,
p3_instqueue_reg_10__1_, p3_instqueue_reg_10__0_,
p3_instqueue_reg_9__7_, p3_instqueue_reg_9__6_, p3_instqueue_reg_9__5_,
p3_instqueue_reg_9__4_, p3_instqueue_reg_9__3_, p3_instqueue_reg_9__2_,
p3_instqueue_reg_9__1_, p3_instqueue_reg_9__0_, p3_instqueue_reg_8__7_,
p3_instqueue_reg_8__6_, p3_instqueue_reg_8__5_, p3_instqueue_reg_8__4_,
p3_instqueue_reg_8__3_, p3_instqueue_reg_8__2_, p3_instqueue_reg_8__1_,
p3_instqueue_reg_8__0_, p3_instqueue_reg_7__7_, p3_instqueue_reg_7__6_,
p3_instqueue_reg_7__5_, p3_instqueue_reg_7__4_, p3_instqueue_reg_7__3_,
p3_instqueue_reg_7__2_, p3_instqueue_reg_7__1_, p3_instqueue_reg_7__0_,
p3_instqueue_reg_6__7_, p3_instqueue_reg_6__6_, p3_instqueue_reg_6__5_,
p3_instqueue_reg_6__4_, p3_instqueue_reg_6__3_, p3_instqueue_reg_6__2_,
p3_instqueue_reg_6__1_, p3_instqueue_reg_6__0_, p3_instqueue_reg_5__7_,
p3_instqueue_reg_5__6_, p3_instqueue_reg_5__5_, p3_instqueue_reg_5__4_,
p3_instqueue_reg_5__3_, p3_instqueue_reg_5__2_, p3_instqueue_reg_5__1_,
p3_instqueue_reg_5__0_, p3_instqueue_reg_4__7_, p3_instqueue_reg_4__6_,
p3_instqueue_reg_4__5_, p3_instqueue_reg_4__4_, p3_instqueue_reg_4__3_,
p3_instqueue_reg_4__2_, p3_instqueue_reg_4__1_, p3_instqueue_reg_4__0_,
p3_instqueue_reg_3__7_, p3_instqueue_reg_3__6_, p3_instqueue_reg_3__5_,
p3_instqueue_reg_3__4_, p3_instqueue_reg_3__3_, p3_instqueue_reg_3__2_,
p3_instqueue_reg_3__1_, p3_instqueue_reg_3__0_, p3_instqueue_reg_2__7_,
p3_instqueue_reg_2__6_, p3_instqueue_reg_2__5_, p3_instqueue_reg_2__4_,
p3_instqueue_reg_2__3_, p3_instqueue_reg_2__2_, p3_instqueue_reg_2__1_,
p3_instqueue_reg_2__0_, p3_instqueue_reg_1__7_, p3_instqueue_reg_1__6_,
p3_instqueue_reg_1__5_, p3_instqueue_reg_1__4_, p3_instqueue_reg_1__3_,
p3_instqueue_reg_1__2_, p3_instqueue_reg_1__1_, p3_instqueue_reg_1__0_,
p3_instqueue_reg_0__7_, p3_instqueue_reg_0__6_, p3_instqueue_reg_0__5_,
p3_instqueue_reg_0__4_, p3_instqueue_reg_0__3_, p3_instqueue_reg_0__2_,
p3_instqueue_reg_0__1_, p3_instqueue_reg_0__0_,
p3_instqueuerd_addr_reg_4_, p3_instqueuerd_addr_reg_3_,
p3_instqueuerd_addr_reg_2_, p3_instqueuerd_addr_reg_1_,
p3_instqueuerd_addr_reg_0_, p3_instqueuewr_addr_reg_4_,
p3_instqueuewr_addr_reg_3_, p3_instqueuewr_addr_reg_2_,
p3_instqueuewr_addr_reg_1_, p3_instqueuewr_addr_reg_0_,
p3_instaddrpointer_reg_0_, p3_instaddrpointer_reg_1_,
p3_instaddrpointer_reg_2_, p3_instaddrpointer_reg_3_,
p3_instaddrpointer_reg_4_, p3_instaddrpointer_reg_5_,
p3_instaddrpointer_reg_6_, p3_instaddrpointer_reg_7_,
p3_instaddrpointer_reg_8_, p3_instaddrpointer_reg_9_,
p3_instaddrpointer_reg_10_, p3_instaddrpointer_reg_11_,
p3_instaddrpointer_reg_12_, p3_instaddrpointer_reg_13_,
p3_instaddrpointer_reg_14_, p3_instaddrpointer_reg_15_,
p3_instaddrpointer_reg_16_, p3_instaddrpointer_reg_17_,
p3_instaddrpointer_reg_18_, p3_instaddrpointer_reg_19_,
p3_instaddrpointer_reg_20_, p3_instaddrpointer_reg_21_,
p3_instaddrpointer_reg_22_, p3_instaddrpointer_reg_23_,
p3_instaddrpointer_reg_24_, p3_instaddrpointer_reg_25_,
p3_instaddrpointer_reg_26_, p3_instaddrpointer_reg_27_,
p3_instaddrpointer_reg_28_, p3_instaddrpointer_reg_29_,
p3_instaddrpointer_reg_30_, p3_instaddrpointer_reg_31_,
p3_phyaddrpointer_reg_0_, p3_phyaddrpointer_reg_1_,
p3_phyaddrpointer_reg_2_, p3_phyaddrpointer_reg_3_,
p3_phyaddrpointer_reg_4_, p3_phyaddrpointer_reg_5_,
p3_phyaddrpointer_reg_6_, p3_phyaddrpointer_reg_7_,
p3_phyaddrpointer_reg_8_, p3_phyaddrpointer_reg_9_,
p3_phyaddrpointer_reg_10_, p3_phyaddrpointer_reg_11_,
p3_phyaddrpointer_reg_12_, p3_phyaddrpointer_reg_13_,
p3_phyaddrpointer_reg_14_, p3_phyaddrpointer_reg_15_,
p3_phyaddrpointer_reg_16_, p3_phyaddrpointer_reg_17_,
p3_phyaddrpointer_reg_18_, p3_phyaddrpointer_reg_19_,
p3_phyaddrpointer_reg_20_, p3_phyaddrpointer_reg_21_,
p3_phyaddrpointer_reg_22_, p3_phyaddrpointer_reg_23_,
p3_phyaddrpointer_reg_24_, p3_phyaddrpointer_reg_25_,
p3_phyaddrpointer_reg_26_, p3_phyaddrpointer_reg_27_,
p3_phyaddrpointer_reg_28_, p3_phyaddrpointer_reg_29_,
p3_phyaddrpointer_reg_30_, p3_phyaddrpointer_reg_31_, p3_lword_reg_15_,
p3_lword_reg_14_, p3_lword_reg_13_, p3_lword_reg_12_, p3_lword_reg_11_,
p3_lword_reg_10_, p3_lword_reg_9_, p3_lword_reg_8_, p3_lword_reg_7_,
p3_lword_reg_6_, p3_lword_reg_5_, p3_lword_reg_4_, p3_lword_reg_3_,
p3_lword_reg_2_, p3_lword_reg_1_, p3_lword_reg_0_, p3_uword_reg_14_,
p3_uword_reg_13_, p3_uword_reg_12_, p3_uword_reg_11_, p3_uword_reg_10_,
p3_uword_reg_9_, p3_uword_reg_8_, p3_uword_reg_7_, p3_uword_reg_6_,
p3_uword_reg_5_, p3_uword_reg_4_, p3_uword_reg_3_, p3_uword_reg_2_,
p3_uword_reg_1_, p3_uword_reg_0_, p3_datao_reg_0_, p3_datao_reg_1_,
p3_datao_reg_2_, p3_datao_reg_3_, p3_datao_reg_4_, p3_datao_reg_5_,
p3_datao_reg_6_, p3_datao_reg_7_, p3_datao_reg_8_, p3_datao_reg_9_,
p3_datao_reg_10_, p3_datao_reg_11_, p3_datao_reg_12_, p3_datao_reg_13_,
p3_datao_reg_14_, p3_datao_reg_15_, p3_datao_reg_16_, p3_datao_reg_17_,
p3_datao_reg_18_, p3_datao_reg_19_, p3_datao_reg_20_, p3_datao_reg_21_,
p3_datao_reg_22_, p3_datao_reg_23_, p3_datao_reg_24_, p3_datao_reg_25_,
p3_datao_reg_26_, p3_datao_reg_27_, p3_datao_reg_28_, p3_datao_reg_29_,
p3_datao_reg_30_, p3_datao_reg_31_, p3_eax_reg_0_, p3_eax_reg_1_,
p3_eax_reg_2_, p3_eax_reg_3_, p3_eax_reg_4_, p3_eax_reg_5_,
p3_eax_reg_6_, p3_eax_reg_7_, p3_eax_reg_8_, p3_eax_reg_9_,
p3_eax_reg_10_, p3_eax_reg_11_, p3_eax_reg_12_, p3_eax_reg_13_,
p3_eax_reg_14_, p3_eax_reg_15_, p3_eax_reg_16_, p3_eax_reg_17_,
p3_eax_reg_18_, p3_eax_reg_19_, p3_eax_reg_20_, p3_eax_reg_21_,
p3_eax_reg_22_, p3_eax_reg_23_, p3_eax_reg_24_, p3_eax_reg_25_,
p3_eax_reg_26_, p3_eax_reg_27_, p3_eax_reg_28_, p3_eax_reg_29_,
p3_eax_reg_30_, p3_eax_reg_31_, p3_ebx_reg_0_, p3_ebx_reg_1_,
p3_ebx_reg_2_, p3_ebx_reg_3_, p3_ebx_reg_4_, p3_ebx_reg_5_,
p3_ebx_reg_6_, p3_ebx_reg_7_, p3_ebx_reg_8_, p3_ebx_reg_9_,
p3_ebx_reg_10_, p3_ebx_reg_11_, p3_ebx_reg_12_, p3_ebx_reg_13_,
p3_ebx_reg_14_, p3_ebx_reg_15_, p3_ebx_reg_16_, p3_ebx_reg_17_,
p3_ebx_reg_18_, p3_ebx_reg_19_, p3_ebx_reg_20_, p3_ebx_reg_21_,
p3_ebx_reg_22_, p3_ebx_reg_23_, p3_ebx_reg_24_, p3_ebx_reg_25_,
p3_ebx_reg_26_, p3_ebx_reg_27_, p3_ebx_reg_28_, p3_ebx_reg_29_,
p3_ebx_reg_30_, p3_ebx_reg_31_, p3_reip_reg_0_, p3_reip_reg_1_,
p3_reip_reg_2_, p3_reip_reg_3_, p3_reip_reg_4_, p3_reip_reg_5_,
p3_reip_reg_6_, p3_reip_reg_7_, p3_reip_reg_8_, p3_reip_reg_9_,
p3_reip_reg_10_, p3_reip_reg_11_, p3_reip_reg_12_, p3_reip_reg_13_,
p3_reip_reg_14_, p3_reip_reg_15_, p3_reip_reg_16_, p3_reip_reg_17_,
p3_reip_reg_18_, p3_reip_reg_19_, p3_reip_reg_20_, p3_reip_reg_21_,
p3_reip_reg_22_, p3_reip_reg_23_, p3_reip_reg_24_, p3_reip_reg_25_,
p3_reip_reg_26_, p3_reip_reg_27_, p3_reip_reg_28_, p3_reip_reg_29_,
p3_reip_reg_30_, p3_reip_reg_31_, p3_byteenable_reg_3_,
p3_byteenable_reg_2_, p3_byteenable_reg_1_, p3_byteenable_reg_0_,
p3_w_r_n_reg, p3_flush_reg, p3_more_reg, p3_statebs16_reg,
p3_requestpending_reg, p3_d_c_n_reg, p3_m_io_n_reg, p3_codefetch_reg,
p3_ads_n_reg, p3_readrequest_reg, p3_memoryfetch_reg, p2_be_n_reg_3_,
p2_be_n_reg_2_, p2_be_n_reg_1_, p2_be_n_reg_0_, p2_address_reg_29_,
p2_address_reg_28_, p2_address_reg_27_, p2_address_reg_26_,
p2_address_reg_25_, p2_address_reg_24_, p2_address_reg_23_,
p2_address_reg_22_, p2_address_reg_21_, p2_address_reg_20_,
p2_address_reg_19_, p2_address_reg_18_, p2_address_reg_17_,
p2_address_reg_16_, p2_address_reg_15_, p2_address_reg_14_,
p2_address_reg_13_, p2_address_reg_12_, p2_address_reg_11_,
p2_address_reg_10_, p2_address_reg_9_, p2_address_reg_8_,
p2_address_reg_7_, p2_address_reg_6_, p2_address_reg_5_,
p2_address_reg_4_, p2_address_reg_3_, p2_address_reg_2_,
p2_address_reg_1_, p2_address_reg_0_, p2_state_reg_2_, p2_state_reg_1_,
p2_state_reg_0_, p2_datawidth_reg_0_, p2_datawidth_reg_1_,
p2_datawidth_reg_2_, p2_datawidth_reg_3_, p2_datawidth_reg_4_,
p2_datawidth_reg_5_, p2_datawidth_reg_6_, p2_datawidth_reg_7_,
p2_datawidth_reg_8_, p2_datawidth_reg_9_, p2_datawidth_reg_10_,
p2_datawidth_reg_11_, p2_datawidth_reg_12_, p2_datawidth_reg_13_,
p2_datawidth_reg_14_, p2_datawidth_reg_15_, p2_datawidth_reg_16_,
p2_datawidth_reg_17_, p2_datawidth_reg_18_, p2_datawidth_reg_19_,
p2_datawidth_reg_20_, p2_datawidth_reg_21_, p2_datawidth_reg_22_,
p2_datawidth_reg_23_, p2_datawidth_reg_24_, p2_datawidth_reg_25_,
p2_datawidth_reg_26_, p2_datawidth_reg_27_, p2_datawidth_reg_28_,
p2_datawidth_reg_29_, p2_datawidth_reg_30_, p2_datawidth_reg_31_,
p2_state2_reg_3_, p2_state2_reg_2_, p2_state2_reg_1_, p2_state2_reg_0_,
p2_instqueue_reg_15__7_, p2_instqueue_reg_15__6_,
p2_instqueue_reg_15__5_, p2_instqueue_reg_15__4_,
p2_instqueue_reg_15__3_, p2_instqueue_reg_15__2_,
p2_instqueue_reg_15__1_, p2_instqueue_reg_15__0_,
p2_instqueue_reg_14__7_, p2_instqueue_reg_14__6_,
p2_instqueue_reg_14__5_, p2_instqueue_reg_14__4_,
p2_instqueue_reg_14__3_, p2_instqueue_reg_14__2_,
p2_instqueue_reg_14__1_, p2_instqueue_reg_14__0_,
p2_instqueue_reg_13__7_, p2_instqueue_reg_13__6_,
p2_instqueue_reg_13__5_, p2_instqueue_reg_13__4_,
p2_instqueue_reg_13__3_, p2_instqueue_reg_13__2_,
p2_instqueue_reg_13__1_, p2_instqueue_reg_13__0_,
p2_instqueue_reg_12__7_, p2_instqueue_reg_12__6_,
p2_instqueue_reg_12__5_, p2_instqueue_reg_12__4_,
p2_instqueue_reg_12__3_, p2_instqueue_reg_12__2_,
p2_instqueue_reg_12__1_, p2_instqueue_reg_12__0_,
p2_instqueue_reg_11__7_, p2_instqueue_reg_11__6_,
p2_instqueue_reg_11__5_, p2_instqueue_reg_11__4_,
p2_instqueue_reg_11__3_, p2_instqueue_reg_11__2_,
p2_instqueue_reg_11__1_, p2_instqueue_reg_11__0_,
p2_instqueue_reg_10__7_, p2_instqueue_reg_10__6_,
p2_instqueue_reg_10__5_, p2_instqueue_reg_10__4_,
p2_instqueue_reg_10__3_, p2_instqueue_reg_10__2_,
p2_instqueue_reg_10__1_, p2_instqueue_reg_10__0_,
p2_instqueue_reg_9__7_, p2_instqueue_reg_9__6_, p2_instqueue_reg_9__5_,
p2_instqueue_reg_9__4_, p2_instqueue_reg_9__3_, p2_instqueue_reg_9__2_,
p2_instqueue_reg_9__1_, p2_instqueue_reg_9__0_, p2_instqueue_reg_8__7_,
p2_instqueue_reg_8__6_, p2_instqueue_reg_8__5_, p2_instqueue_reg_8__4_,
p2_instqueue_reg_8__3_, p2_instqueue_reg_8__2_, p2_instqueue_reg_8__1_,
p2_instqueue_reg_8__0_, p2_instqueue_reg_7__7_, p2_instqueue_reg_7__6_,
p2_instqueue_reg_7__5_, p2_instqueue_reg_7__4_, p2_instqueue_reg_7__3_,
p2_instqueue_reg_7__2_, p2_instqueue_reg_7__1_, p2_instqueue_reg_7__0_,
p2_instqueue_reg_6__7_, p2_instqueue_reg_6__6_, p2_instqueue_reg_6__5_,
p2_instqueue_reg_6__4_, p2_instqueue_reg_6__3_, p2_instqueue_reg_6__2_,
p2_instqueue_reg_6__1_, p2_instqueue_reg_6__0_, p2_instqueue_reg_5__7_,
p2_instqueue_reg_5__6_, p2_instqueue_reg_5__5_, p2_instqueue_reg_5__4_,
p2_instqueue_reg_5__3_, p2_instqueue_reg_5__2_, p2_instqueue_reg_5__1_,
p2_instqueue_reg_5__0_, p2_instqueue_reg_4__7_, p2_instqueue_reg_4__6_,
p2_instqueue_reg_4__5_, p2_instqueue_reg_4__4_, p2_instqueue_reg_4__3_,
p2_instqueue_reg_4__2_, p2_instqueue_reg_4__1_, p2_instqueue_reg_4__0_,
p2_instqueue_reg_3__7_, p2_instqueue_reg_3__6_, p2_instqueue_reg_3__5_,
p2_instqueue_reg_3__4_, p2_instqueue_reg_3__3_, p2_instqueue_reg_3__2_,
p2_instqueue_reg_3__1_, p2_instqueue_reg_3__0_, p2_instqueue_reg_2__7_,
p2_instqueue_reg_2__6_, p2_instqueue_reg_2__5_, p2_instqueue_reg_2__4_,
p2_instqueue_reg_2__3_, p2_instqueue_reg_2__2_, p2_instqueue_reg_2__1_,
p2_instqueue_reg_2__0_, p2_instqueue_reg_1__7_, p2_instqueue_reg_1__6_,
p2_instqueue_reg_1__5_, p2_instqueue_reg_1__4_, p2_instqueue_reg_1__3_,
p2_instqueue_reg_1__2_, p2_instqueue_reg_1__1_, p2_instqueue_reg_1__0_,
p2_instqueue_reg_0__7_, p2_instqueue_reg_0__6_, p2_instqueue_reg_0__5_,
p2_instqueue_reg_0__4_, p2_instqueue_reg_0__3_, p2_instqueue_reg_0__2_,
p2_instqueue_reg_0__1_, p2_instqueue_reg_0__0_,
p2_instqueuerd_addr_reg_4_, p2_instqueuerd_addr_reg_3_,
p2_instqueuerd_addr_reg_2_, p2_instqueuerd_addr_reg_1_,
p2_instqueuerd_addr_reg_0_, p2_instqueuewr_addr_reg_4_,
p2_instqueuewr_addr_reg_3_, p2_instqueuewr_addr_reg_2_,
p2_instqueuewr_addr_reg_1_, p2_instqueuewr_addr_reg_0_,
p2_instaddrpointer_reg_0_, p2_instaddrpointer_reg_1_,
p2_instaddrpointer_reg_2_, p2_instaddrpointer_reg_3_,
p2_instaddrpointer_reg_4_, p2_instaddrpointer_reg_5_,
p2_instaddrpointer_reg_6_, p2_instaddrpointer_reg_7_,
p2_instaddrpointer_reg_8_, p2_instaddrpointer_reg_9_,
p2_instaddrpointer_reg_10_, p2_instaddrpointer_reg_11_,
p2_instaddrpointer_reg_12_, p2_instaddrpointer_reg_13_,
p2_instaddrpointer_reg_14_, p2_instaddrpointer_reg_15_,
p2_instaddrpointer_reg_16_, p2_instaddrpointer_reg_17_,
p2_instaddrpointer_reg_18_, p2_instaddrpointer_reg_19_,
p2_instaddrpointer_reg_20_, p2_instaddrpointer_reg_21_,
p2_instaddrpointer_reg_22_, p2_instaddrpointer_reg_23_,
p2_instaddrpointer_reg_24_, p2_instaddrpointer_reg_25_,
p2_instaddrpointer_reg_26_, p2_instaddrpointer_reg_27_,
p2_instaddrpointer_reg_28_, p2_instaddrpointer_reg_29_,
p2_instaddrpointer_reg_30_, p2_instaddrpointer_reg_31_,
p2_phyaddrpointer_reg_0_, p2_phyaddrpointer_reg_1_,
p2_phyaddrpointer_reg_2_, p2_phyaddrpointer_reg_3_,
p2_phyaddrpointer_reg_4_, p2_phyaddrpointer_reg_5_,
p2_phyaddrpointer_reg_6_, p2_phyaddrpointer_reg_7_,
p2_phyaddrpointer_reg_8_, p2_phyaddrpointer_reg_9_,
p2_phyaddrpointer_reg_10_, p2_phyaddrpointer_reg_11_,
p2_phyaddrpointer_reg_12_, p2_phyaddrpointer_reg_13_,
p2_phyaddrpointer_reg_14_, p2_phyaddrpointer_reg_15_,
p2_phyaddrpointer_reg_16_, p2_phyaddrpointer_reg_17_,
p2_phyaddrpointer_reg_18_, p2_phyaddrpointer_reg_19_,
p2_phyaddrpointer_reg_20_, p2_phyaddrpointer_reg_21_,
p2_phyaddrpointer_reg_22_, p2_phyaddrpointer_reg_23_,
p2_phyaddrpointer_reg_24_, p2_phyaddrpointer_reg_25_,
p2_phyaddrpointer_reg_26_, p2_phyaddrpointer_reg_27_,
p2_phyaddrpointer_reg_28_, p2_phyaddrpointer_reg_29_,
p2_phyaddrpointer_reg_30_, p2_phyaddrpointer_reg_31_, p2_lword_reg_15_,
p2_lword_reg_14_, p2_lword_reg_13_, p2_lword_reg_12_, p2_lword_reg_11_,
p2_lword_reg_10_, p2_lword_reg_9_, p2_lword_reg_8_, p2_lword_reg_7_,
p2_lword_reg_6_, p2_lword_reg_5_, p2_lword_reg_4_, p2_lword_reg_3_,
p2_lword_reg_2_, p2_lword_reg_1_, p2_lword_reg_0_, p2_uword_reg_14_,
p2_uword_reg_13_, p2_uword_reg_12_, p2_uword_reg_11_, p2_uword_reg_10_,
p2_uword_reg_9_, p2_uword_reg_8_, p2_uword_reg_7_, p2_uword_reg_6_,
p2_uword_reg_5_, p2_uword_reg_4_, p2_uword_reg_3_, p2_uword_reg_2_,
p2_uword_reg_1_, p2_uword_reg_0_, p2_datao_reg_0_, p2_datao_reg_1_,
p2_datao_reg_2_, p2_datao_reg_3_, p2_datao_reg_4_, p2_datao_reg_5_,
p2_datao_reg_6_, p2_datao_reg_7_, p2_datao_reg_8_, p2_datao_reg_9_,
p2_datao_reg_10_, p2_datao_reg_11_, p2_datao_reg_12_, p2_datao_reg_13_,
p2_datao_reg_14_, p2_datao_reg_15_, p2_datao_reg_16_, p2_datao_reg_17_,
p2_datao_reg_18_, p2_datao_reg_19_, p2_datao_reg_20_, p2_datao_reg_21_,
p2_datao_reg_22_, p2_datao_reg_23_, p2_datao_reg_24_, p2_datao_reg_25_,
p2_datao_reg_26_, p2_datao_reg_27_, p2_datao_reg_28_, p2_datao_reg_29_,
p2_datao_reg_30_, p2_datao_reg_31_, p2_eax_reg_0_, p2_eax_reg_1_,
p2_eax_reg_2_, p2_eax_reg_3_, p2_eax_reg_4_, p2_eax_reg_5_,
p2_eax_reg_6_, p2_eax_reg_7_, p2_eax_reg_8_, p2_eax_reg_9_,
p2_eax_reg_10_, p2_eax_reg_11_, p2_eax_reg_12_, p2_eax_reg_13_,
p2_eax_reg_14_, p2_eax_reg_15_, p2_eax_reg_16_, p2_eax_reg_17_,
p2_eax_reg_18_, p2_eax_reg_19_, p2_eax_reg_20_, p2_eax_reg_21_,
p2_eax_reg_22_, p2_eax_reg_23_, p2_eax_reg_24_, p2_eax_reg_25_,
p2_eax_reg_26_, p2_eax_reg_27_, p2_eax_reg_28_, p2_eax_reg_29_,
p2_eax_reg_30_, p2_eax_reg_31_, p2_ebx_reg_0_, p2_ebx_reg_1_,
p2_ebx_reg_2_, p2_ebx_reg_3_, p2_ebx_reg_4_, p2_ebx_reg_5_,
p2_ebx_reg_6_, p2_ebx_reg_7_, p2_ebx_reg_8_, p2_ebx_reg_9_,
p2_ebx_reg_10_, p2_ebx_reg_11_, p2_ebx_reg_12_, p2_ebx_reg_13_,
p2_ebx_reg_14_, p2_ebx_reg_15_, p2_ebx_reg_16_, p2_ebx_reg_17_,
p2_ebx_reg_18_, p2_ebx_reg_19_, p2_ebx_reg_20_, p2_ebx_reg_21_,
p2_ebx_reg_22_, p2_ebx_reg_23_, p2_ebx_reg_24_, p2_ebx_reg_25_,
p2_ebx_reg_26_, p2_ebx_reg_27_, p2_ebx_reg_28_, p2_ebx_reg_29_,
p2_ebx_reg_30_, p2_ebx_reg_31_, p2_reip_reg_0_, p2_reip_reg_1_,
p2_reip_reg_2_, p2_reip_reg_3_, p2_reip_reg_4_, p2_reip_reg_5_,
p2_reip_reg_6_, p2_reip_reg_7_, p2_reip_reg_8_, p2_reip_reg_9_,
p2_reip_reg_10_, p2_reip_reg_11_, p2_reip_reg_12_, p2_reip_reg_13_,
p2_reip_reg_14_, p2_reip_reg_15_, p2_reip_reg_16_, p2_reip_reg_17_,
p2_reip_reg_18_, p2_reip_reg_19_, p2_reip_reg_20_, p2_reip_reg_21_,
p2_reip_reg_22_, p2_reip_reg_23_, p2_reip_reg_24_, p2_reip_reg_25_,
p2_reip_reg_26_, p2_reip_reg_27_, p2_reip_reg_28_, p2_reip_reg_29_,
p2_reip_reg_30_, p2_reip_reg_31_, p2_byteenable_reg_3_,
p2_byteenable_reg_2_, p2_byteenable_reg_1_, p2_byteenable_reg_0_,
p2_w_r_n_reg, p2_flush_reg, p2_more_reg, p2_statebs16_reg,
p2_requestpending_reg, p2_d_c_n_reg, p2_m_io_n_reg, p2_codefetch_reg,
p2_ads_n_reg, p2_readrequest_reg, p2_memoryfetch_reg, p1_be_n_reg_3_,
p1_be_n_reg_2_, p1_be_n_reg_1_, p1_be_n_reg_0_, p1_state_reg_2_,
p1_state_reg_1_, p1_state_reg_0_, p1_datawidth_reg_0_,
p1_datawidth_reg_1_, p1_datawidth_reg_2_, p1_datawidth_reg_3_,
p1_datawidth_reg_4_, p1_datawidth_reg_5_, p1_datawidth_reg_6_,
p1_datawidth_reg_7_, p1_datawidth_reg_8_, p1_datawidth_reg_9_,
p1_datawidth_reg_10_, p1_datawidth_reg_11_, p1_datawidth_reg_12_,
p1_datawidth_reg_13_, p1_datawidth_reg_14_, p1_datawidth_reg_15_,
p1_datawidth_reg_16_, p1_datawidth_reg_17_, p1_datawidth_reg_18_,
p1_datawidth_reg_19_, p1_datawidth_reg_20_, p1_datawidth_reg_21_,
p1_datawidth_reg_22_, p1_datawidth_reg_23_, p1_datawidth_reg_24_,
p1_datawidth_reg_25_, p1_datawidth_reg_26_, p1_datawidth_reg_27_,
p1_datawidth_reg_28_, p1_datawidth_reg_29_, p1_datawidth_reg_30_,
p1_datawidth_reg_31_, p1_state2_reg_3_, p1_state2_reg_2_,
p1_state2_reg_1_, p1_state2_reg_0_, p1_instqueue_reg_15__7_,
p1_instqueue_reg_15__6_, p1_instqueue_reg_15__5_,
p1_instqueue_reg_15__4_, p1_instqueue_reg_15__3_,
p1_instqueue_reg_15__2_, p1_instqueue_reg_15__1_,
p1_instqueue_reg_15__0_, p1_instqueue_reg_14__7_,
p1_instqueue_reg_14__6_, p1_instqueue_reg_14__5_,
p1_instqueue_reg_14__4_, p1_instqueue_reg_14__3_,
p1_instqueue_reg_14__2_, p1_instqueue_reg_14__1_,
p1_instqueue_reg_14__0_, p1_instqueue_reg_13__7_,
p1_instqueue_reg_13__6_, p1_instqueue_reg_13__5_,
p1_instqueue_reg_13__4_, p1_instqueue_reg_13__3_,
p1_instqueue_reg_13__2_, p1_instqueue_reg_13__1_,
p1_instqueue_reg_13__0_, p1_instqueue_reg_12__7_,
p1_instqueue_reg_12__6_, p1_instqueue_reg_12__5_,
p1_instqueue_reg_12__4_, p1_instqueue_reg_12__3_,
p1_instqueue_reg_12__2_, p1_instqueue_reg_12__1_,
p1_instqueue_reg_12__0_, p1_instqueue_reg_11__7_,
p1_instqueue_reg_11__6_, p1_instqueue_reg_11__5_,
p1_instqueue_reg_11__4_, p1_instqueue_reg_11__3_,
p1_instqueue_reg_11__2_, p1_instqueue_reg_11__1_,
p1_instqueue_reg_11__0_, p1_instqueue_reg_10__7_,
p1_instqueue_reg_10__6_, p1_instqueue_reg_10__5_,
p1_instqueue_reg_10__4_, p1_instqueue_reg_10__3_,
p1_instqueue_reg_10__2_, p1_instqueue_reg_10__1_,
p1_instqueue_reg_10__0_, p1_instqueue_reg_9__7_,
p1_instqueue_reg_9__6_, p1_instqueue_reg_9__5_, p1_instqueue_reg_9__4_,
p1_instqueue_reg_9__3_, p1_instqueue_reg_9__2_, p1_instqueue_reg_9__1_,
p1_instqueue_reg_9__0_, p1_instqueue_reg_8__7_, p1_instqueue_reg_8__6_,
p1_instqueue_reg_8__5_, p1_instqueue_reg_8__4_, p1_instqueue_reg_8__3_,
p1_instqueue_reg_8__2_, p1_instqueue_reg_8__1_, p1_instqueue_reg_8__0_,
p1_instqueue_reg_7__7_, p1_instqueue_reg_7__6_, p1_instqueue_reg_7__5_,
p1_instqueue_reg_7__4_, p1_instqueue_reg_7__3_, p1_instqueue_reg_7__2_,
p1_instqueue_reg_7__1_, p1_instqueue_reg_7__0_, p1_instqueue_reg_6__7_,
p1_instqueue_reg_6__6_, p1_instqueue_reg_6__5_, p1_instqueue_reg_6__4_,
p1_instqueue_reg_6__3_, p1_instqueue_reg_6__2_, p1_instqueue_reg_6__1_,
p1_instqueue_reg_6__0_, p1_instqueue_reg_5__7_, p1_instqueue_reg_5__6_,
p1_instqueue_reg_5__5_, p1_instqueue_reg_5__4_, p1_instqueue_reg_5__3_,
p1_instqueue_reg_5__2_, p1_instqueue_reg_5__1_, p1_instqueue_reg_5__0_,
p1_instqueue_reg_4__7_, p1_instqueue_reg_4__6_, p1_instqueue_reg_4__5_,
p1_instqueue_reg_4__4_, p1_instqueue_reg_4__3_, p1_instqueue_reg_4__2_,
p1_instqueue_reg_4__1_, p1_instqueue_reg_4__0_, p1_instqueue_reg_3__7_,
p1_instqueue_reg_3__6_, p1_instqueue_reg_3__5_, p1_instqueue_reg_3__4_,
p1_instqueue_reg_3__3_, p1_instqueue_reg_3__2_, p1_instqueue_reg_3__1_,
p1_instqueue_reg_3__0_, p1_instqueue_reg_2__7_, p1_instqueue_reg_2__6_,
p1_instqueue_reg_2__5_, p1_instqueue_reg_2__4_, p1_instqueue_reg_2__3_,
p1_instqueue_reg_2__2_, p1_instqueue_reg_2__1_, p1_instqueue_reg_2__0_,
p1_instqueue_reg_1__7_, p1_instqueue_reg_1__6_, p1_instqueue_reg_1__5_,
p1_instqueue_reg_1__4_, p1_instqueue_reg_1__3_, p1_instqueue_reg_1__2_,
p1_instqueue_reg_1__1_, p1_instqueue_reg_1__0_, p1_instqueue_reg_0__7_,
p1_instqueue_reg_0__6_, p1_instqueue_reg_0__5_, p1_instqueue_reg_0__4_,
p1_instqueue_reg_0__3_, p1_instqueue_reg_0__2_, p1_instqueue_reg_0__1_,
p1_instqueue_reg_0__0_, p1_instqueuerd_addr_reg_4_,
p1_instqueuerd_addr_reg_3_, p1_instqueuerd_addr_reg_2_,
p1_instqueuerd_addr_reg_1_, p1_instqueuerd_addr_reg_0_,
p1_instqueuewr_addr_reg_4_, p1_instqueuewr_addr_reg_3_,
p1_instqueuewr_addr_reg_2_, p1_instqueuewr_addr_reg_1_,
p1_instqueuewr_addr_reg_0_, p1_instaddrpointer_reg_0_,
p1_instaddrpointer_reg_1_, p1_instaddrpointer_reg_2_,
p1_instaddrpointer_reg_3_, p1_instaddrpointer_reg_4_,
p1_instaddrpointer_reg_5_, p1_instaddrpointer_reg_6_,
p1_instaddrpointer_reg_7_, p1_instaddrpointer_reg_8_,
p1_instaddrpointer_reg_9_, p1_instaddrpointer_reg_10_,
p1_instaddrpointer_reg_11_, p1_instaddrpointer_reg_12_,
p1_instaddrpointer_reg_13_, p1_instaddrpointer_reg_14_,
p1_instaddrpointer_reg_15_, p1_instaddrpointer_reg_16_,
p1_instaddrpointer_reg_17_, p1_instaddrpointer_reg_18_,
p1_instaddrpointer_reg_19_, p1_instaddrpointer_reg_20_,
p1_instaddrpointer_reg_21_, p1_instaddrpointer_reg_22_,
p1_instaddrpointer_reg_23_, p1_instaddrpointer_reg_24_,
p1_instaddrpointer_reg_25_, p1_instaddrpointer_reg_26_,
p1_instaddrpointer_reg_27_, p1_instaddrpointer_reg_28_,
p1_instaddrpointer_reg_29_, p1_instaddrpointer_reg_30_,
p1_instaddrpointer_reg_31_, p1_phyaddrpointer_reg_0_,
p1_phyaddrpointer_reg_1_, p1_phyaddrpointer_reg_2_,
p1_phyaddrpointer_reg_3_, p1_phyaddrpointer_reg_4_,
p1_phyaddrpointer_reg_5_, p1_phyaddrpointer_reg_6_,
p1_phyaddrpointer_reg_7_, p1_phyaddrpointer_reg_8_,
p1_phyaddrpointer_reg_9_, p1_phyaddrpointer_reg_10_,
p1_phyaddrpointer_reg_11_, p1_phyaddrpointer_reg_12_,
p1_phyaddrpointer_reg_13_, p1_phyaddrpointer_reg_14_,
p1_phyaddrpointer_reg_15_, p1_phyaddrpointer_reg_16_,
p1_phyaddrpointer_reg_17_, p1_phyaddrpointer_reg_18_,
p1_phyaddrpointer_reg_19_, p1_phyaddrpointer_reg_20_,
p1_phyaddrpointer_reg_21_, p1_phyaddrpointer_reg_22_,
p1_phyaddrpointer_reg_23_, p1_phyaddrpointer_reg_24_,
p1_phyaddrpointer_reg_25_, p1_phyaddrpointer_reg_26_,
p1_phyaddrpointer_reg_27_, p1_phyaddrpointer_reg_28_,
p1_phyaddrpointer_reg_29_, p1_phyaddrpointer_reg_30_,
p1_phyaddrpointer_reg_31_, p1_lword_reg_15_, p1_lword_reg_14_,
p1_lword_reg_13_, p1_lword_reg_12_, p1_lword_reg_11_, p1_lword_reg_10_,
p1_lword_reg_9_, p1_lword_reg_8_, p1_lword_reg_7_, p1_lword_reg_6_,
p1_lword_reg_5_, p1_lword_reg_4_, p1_lword_reg_3_, p1_lword_reg_2_,
p1_lword_reg_1_, p1_lword_reg_0_, p1_uword_reg_14_, p1_uword_reg_13_,
p1_uword_reg_12_, p1_uword_reg_11_, p1_uword_reg_10_, p1_uword_reg_9_,
p1_uword_reg_8_, p1_uword_reg_7_, p1_uword_reg_6_, p1_uword_reg_5_,
p1_uword_reg_4_, p1_uword_reg_3_, p1_uword_reg_2_, p1_uword_reg_1_,
p1_uword_reg_0_, p1_datao_reg_0_, p1_datao_reg_1_, p1_datao_reg_2_,
p1_datao_reg_3_, p1_datao_reg_4_, p1_datao_reg_5_, p1_datao_reg_6_,
p1_datao_reg_7_, p1_datao_reg_8_, p1_datao_reg_9_, p1_datao_reg_10_,
p1_datao_reg_11_, p1_datao_reg_12_, p1_datao_reg_13_, p1_datao_reg_14_,
p1_datao_reg_15_, p1_datao_reg_16_, p1_datao_reg_17_, p1_datao_reg_18_,
p1_datao_reg_19_, p1_datao_reg_20_, p1_datao_reg_21_, p1_datao_reg_22_,
p1_datao_reg_23_, p1_datao_reg_24_, p1_datao_reg_25_, p1_datao_reg_26_,
p1_datao_reg_27_, p1_datao_reg_28_, p1_datao_reg_29_, p1_datao_reg_30_,
p1_datao_reg_31_, p1_eax_reg_0_, p1_eax_reg_1_, p1_eax_reg_2_,
p1_eax_reg_3_, p1_eax_reg_4_, p1_eax_reg_5_, p1_eax_reg_6_,
p1_eax_reg_7_, p1_eax_reg_8_, p1_eax_reg_9_, p1_eax_reg_10_,
p1_eax_reg_11_, p1_eax_reg_12_, p1_eax_reg_13_, p1_eax_reg_14_,
p1_eax_reg_15_, p1_eax_reg_16_, p1_eax_reg_17_, p1_eax_reg_18_,
p1_eax_reg_19_, p1_eax_reg_20_, p1_eax_reg_21_, p1_eax_reg_22_,
p1_eax_reg_23_, p1_eax_reg_24_, p1_eax_reg_25_, p1_eax_reg_26_,
p1_eax_reg_27_, p1_eax_reg_28_, p1_eax_reg_29_, p1_eax_reg_30_,
p1_eax_reg_31_, p1_ebx_reg_0_, p1_ebx_reg_1_, p1_ebx_reg_2_,
p1_ebx_reg_3_, p1_ebx_reg_4_, p1_ebx_reg_5_, p1_ebx_reg_6_,
p1_ebx_reg_7_, p1_ebx_reg_8_, p1_ebx_reg_9_, p1_ebx_reg_10_,
p1_ebx_reg_11_, p1_ebx_reg_12_, p1_ebx_reg_13_, p1_ebx_reg_14_,
p1_ebx_reg_15_, p1_ebx_reg_16_, p1_ebx_reg_17_, p1_ebx_reg_18_,
p1_ebx_reg_19_, p1_ebx_reg_20_, p1_ebx_reg_21_, p1_ebx_reg_22_,
p1_ebx_reg_23_, p1_ebx_reg_24_, p1_ebx_reg_25_, p1_ebx_reg_26_,
p1_ebx_reg_27_, p1_ebx_reg_28_, p1_ebx_reg_29_, p1_ebx_reg_30_,
p1_ebx_reg_31_, p1_reip_reg_0_, p1_reip_reg_1_, p1_reip_reg_2_,
p1_reip_reg_3_, p1_reip_reg_4_, p1_reip_reg_5_, p1_reip_reg_6_,
p1_reip_reg_7_, p1_reip_reg_8_, p1_reip_reg_9_, p1_reip_reg_10_,
p1_reip_reg_11_, p1_reip_reg_12_, p1_reip_reg_13_, p1_reip_reg_14_,
p1_reip_reg_15_, p1_reip_reg_16_, p1_reip_reg_17_, p1_reip_reg_18_,
p1_reip_reg_19_, p1_reip_reg_20_, p1_reip_reg_21_, p1_reip_reg_22_,
p1_reip_reg_23_, p1_reip_reg_24_, p1_reip_reg_25_, p1_reip_reg_26_,
p1_reip_reg_27_, p1_reip_reg_28_, p1_reip_reg_29_, p1_reip_reg_30_,
p1_reip_reg_31_, p1_byteenable_reg_3_, p1_byteenable_reg_2_,
p1_byteenable_reg_1_, p1_byteenable_reg_0_, p1_w_r_n_reg, p1_flush_reg,
p1_more_reg, p1_statebs16_reg, p1_requestpending_reg, p1_d_c_n_reg,
p1_m_io_n_reg, p1_codefetch_reg, p1_ads_n_reg, p1_readrequest_reg,
p1_memoryfetch_reg, p1_address_reg_29_, p1_address_reg_28_,
p1_address_reg_27_, p1_address_reg_26_, p1_address_reg_25_,
p1_address_reg_24_, p1_address_reg_23_, p1_address_reg_22_,
p1_address_reg_21_, p1_address_reg_20_, p1_address_reg_19_,
p1_address_reg_18_, p1_address_reg_17_, p1_address_reg_16_,
p1_address_reg_15_, p1_address_reg_14_, p1_address_reg_13_,
p1_address_reg_12_, p1_address_reg_11_, p1_address_reg_10_,
p1_address_reg_9_, p1_address_reg_8_, p1_address_reg_7_,
p1_address_reg_6_, p1_address_reg_5_, p1_address_reg_4_,
p1_address_reg_3_, p1_address_reg_2_, p1_address_reg_1_,
p1_address_reg_0_, u355, u356, u357, u358, u359, u360, u361, u362,
u363, u364, u366, u367, u368, u369, u370, u371, u372, u373, u374, u375,
u347, u348, u349, u350, u351, u352, u353, u354, u365, u376, u247, u246,
u245, u244, u243, u242, u241, u240, u239, u238, u237, u236, u235, u234,
u233, u232, u231, u230, u229, u228, u227, u226, u225, u224, u223, u222,
u221, u220, u219, u218, u217, u216, u251, u252, u253, u254, u255, u256,
u257, u258, u259, u260, u261, u262, u263, u264, u265, u266, u267, u268,
u269, u270, u271, u272, u273, u274, u275, u276, u277, u278, u279, u280,
u281, u282, u212, u215, u213, u214, p3_u3274, p3_u3275, p3_u3276,
p3_u3277, p3_u3061, p3_u3060, p3_u3059, p3_u3058, p3_u3057, p3_u3056,
p3_u3055, p3_u3054, p3_u3053, p3_u3052, p3_u3051, p3_u3050, p3_u3049,
p3_u3048, p3_u3047, p3_u3046, p3_u3045, p3_u3044, p3_u3043, p3_u3042,
p3_u3041, p3_u3040, p3_u3039, p3_u3038, p3_u3037, p3_u3036, p3_u3035,
p3_u3034, p3_u3033, p3_u3032, p3_u3031, p3_u3030, p3_u3029, p3_u3280,
p3_u3281, p3_u3028, p3_u3027, p3_u3026, p3_u3025, p3_u3024, p3_u3023,
p3_u3022, p3_u3021, p3_u3020, p3_u3019, p3_u3018, p3_u3017, p3_u3016,
p3_u3015, p3_u3014, p3_u3013, p3_u3012, p3_u3011, p3_u3010, p3_u3009,
p3_u3008, p3_u3007, p3_u3006, p3_u3005, p3_u3004, p3_u3003, p3_u3002,
p3_u3001, p3_u3000, p3_u2999, p3_u3282, p3_u2998, p3_u2997, p3_u2996,
p3_u2995, p3_u2994, p3_u2993, p3_u2992, p3_u2991, p3_u2990, p3_u2989,
p3_u2988, p3_u2987, p3_u2986, p3_u2985, p3_u2984, p3_u2983, p3_u2982,
p3_u2981, p3_u2980, p3_u2979, p3_u2978, p3_u2977, p3_u2976, p3_u2975,
p3_u2974, p3_u2973, p3_u2972, p3_u2971, p3_u2970, p3_u2969, p3_u2968,
p3_u2967, p3_u2966, p3_u2965, p3_u2964, p3_u2963, p3_u2962, p3_u2961,
p3_u2960, p3_u2959, p3_u2958, p3_u2957, p3_u2956, p3_u2955, p3_u2954,
p3_u2953, p3_u2952, p3_u2951, p3_u2950, p3_u2949, p3_u2948, p3_u2947,
p3_u2946, p3_u2945, p3_u2944, p3_u2943, p3_u2942, p3_u2941, p3_u2940,
p3_u2939, p3_u2938, p3_u2937, p3_u2936, p3_u2935, p3_u2934, p3_u2933,
p3_u2932, p3_u2931, p3_u2930, p3_u2929, p3_u2928, p3_u2927, p3_u2926,
p3_u2925, p3_u2924, p3_u2923, p3_u2922, p3_u2921, p3_u2920, p3_u2919,
p3_u2918, p3_u2917, p3_u2916, p3_u2915, p3_u2914, p3_u2913, p3_u2912,
p3_u2911, p3_u2910, p3_u2909, p3_u2908, p3_u2907, p3_u2906, p3_u2905,
p3_u2904, p3_u2903, p3_u2902, p3_u2901, p3_u2900, p3_u2899, p3_u2898,
p3_u2897, p3_u2896, p3_u2895, p3_u2894, p3_u2893, p3_u2892, p3_u2891,
p3_u2890, p3_u2889, p3_u2888, p3_u2887, p3_u2886, p3_u2885, p3_u2884,
p3_u2883, p3_u2882, p3_u2881, p3_u2880, p3_u2879, p3_u2878, p3_u2877,
p3_u2876, p3_u2875, p3_u2874, p3_u2873, p3_u2872, p3_u2871, p3_u2870,
p3_u2869, p3_u2868, p3_u3284, p3_u3285, p3_u3288, p3_u3289, p3_u3290,
p3_u2867, p3_u2866, p3_u2865, p3_u2864, p3_u2863, p3_u2862, p3_u2861,
p3_u2860, p3_u2859, p3_u2858, p3_u2857, p3_u2856, p3_u2855, p3_u2854,
p3_u2853, p3_u2852, p3_u2851, p3_u2850, p3_u2849, p3_u2848, p3_u2847,
p3_u2846, p3_u2845, p3_u2844, p3_u2843, p3_u2842, p3_u2841, p3_u2840,
p3_u2839, p3_u2838, p3_u2837, p3_u2836, p3_u2835, p3_u2834, p3_u2833,
p3_u2832, p3_u2831, p3_u2830, p3_u2829, p3_u2828, p3_u2827, p3_u2826,
p3_u2825, p3_u2824, p3_u2823, p3_u2822, p3_u2821, p3_u2820, p3_u2819,
p3_u2818, p3_u2817, p3_u2816, p3_u2815, p3_u2814, p3_u2813, p3_u2812,
p3_u2811, p3_u2810, p3_u2809, p3_u2808, p3_u2807, p3_u2806, p3_u2805,
p3_u2804, p3_u2803, p3_u2802, p3_u2801, p3_u2800, p3_u2799, p3_u2798,
p3_u2797, p3_u2796, p3_u2795, p3_u2794, p3_u2793, p3_u2792, p3_u2791,
p3_u2790, p3_u2789, p3_u2788, p3_u2787, p3_u2786, p3_u2785, p3_u2784,
p3_u2783, p3_u2782, p3_u2781, p3_u2780, p3_u2779, p3_u2778, p3_u2777,
p3_u2776, p3_u2775, p3_u2774, p3_u2773, p3_u2772, p3_u2771, p3_u2770,
p3_u2769, p3_u2768, p3_u2767, p3_u2766, p3_u2765, p3_u2764, p3_u2763,
p3_u2762, p3_u2761, p3_u2760, p3_u2759, p3_u2758, p3_u2757, p3_u2756,
p3_u2755, p3_u2754, p3_u2753, p3_u2752, p3_u2751, p3_u2750, p3_u2749,
p3_u2748, p3_u2747, p3_u2746, p3_u2745, p3_u2744, p3_u2743, p3_u2742,
p3_u2741, p3_u2740, p3_u2739, p3_u2738, p3_u2737, p3_u2736, p3_u2735,
p3_u2734, p3_u2733, p3_u2732, p3_u2731, p3_u2730, p3_u2729, p3_u2728,
p3_u2727, p3_u2726, p3_u2725, p3_u2724, p3_u2723, p3_u2722, p3_u2721,
p3_u2720, p3_u2719, p3_u2718, p3_u2717, p3_u2716, p3_u2715, p3_u2714,
p3_u2713, p3_u2712, p3_u2711, p3_u2710, p3_u2709, p3_u2708, p3_u2707,
p3_u2706, p3_u2705, p3_u2704, p3_u2703, p3_u2702, p3_u2701, p3_u2700,
p3_u2699, p3_u2698, p3_u2697, p3_u2696, p3_u2695, p3_u2694, p3_u2693,
p3_u2692, p3_u2691, p3_u2690, p3_u2689, p3_u2688, p3_u2687, p3_u2686,
p3_u2685, p3_u2684, p3_u2683, p3_u2682, p3_u2681, p3_u2680, p3_u2679,
p3_u2678, p3_u2677, p3_u2676, p3_u2675, p3_u2674, p3_u2673, p3_u2672,
p3_u2671, p3_u2670, p3_u2669, p3_u2668, p3_u2667, p3_u2666, p3_u2665,
p3_u2664, p3_u2663, p3_u2662, p3_u2661, p3_u2660, p3_u2659, p3_u2658,
p3_u2657, p3_u2656, p3_u2655, p3_u2654, p3_u2653, p3_u2652, p3_u2651,
p3_u2650, p3_u2649, p3_u2648, p3_u2647, p3_u2646, p3_u2645, p3_u2644,
p3_u2643, p3_u2642, p3_u2641, p3_u2640, p3_u2639, p3_u3292, p3_u2638,
p3_u3293, p3_u3294, p3_u2637, p3_u3295, p3_u2636, p3_u3296, p3_u2635,
p3_u3297, p3_u2634, p3_u2633, p3_u3298, p3_u3299, p2_u3585, p2_u3586,
p2_u3587, p2_u3588, p2_u3241, p2_u3240, p2_u3239, p2_u3238, p2_u3237,
p2_u3236, p2_u3235, p2_u3234, p2_u3233, p2_u3232, p2_u3231, p2_u3230,
p2_u3229, p2_u3228, p2_u3227, p2_u3226, p2_u3225, p2_u3224, p2_u3223,
p2_u3222, p2_u3221, p2_u3220, p2_u3219, p2_u3218, p2_u3217, p2_u3216,
p2_u3215, p2_u3214, p2_u3213, p2_u3212, p2_u3211, p2_u3210, p2_u3209,
p2_u3591, p2_u3592, p2_u3208, p2_u3207, p2_u3206, p2_u3205, p2_u3204,
p2_u3203, p2_u3202, p2_u3201, p2_u3200, p2_u3199, p2_u3198, p2_u3197,
p2_u3196, p2_u3195, p2_u3194, p2_u3193, p2_u3192, p2_u3191, p2_u3190,
p2_u3189, p2_u3188, p2_u3187, p2_u3186, p2_u3185, p2_u3184, p2_u3183,
p2_u3182, p2_u3181, p2_u3180, p2_u3179, p2_u3593, p2_u3178, p2_u3177,
p2_u3176, p2_u3175, p2_u3174, p2_u3173, p2_u3172, p2_u3171, p2_u3170,
p2_u3169, p2_u3168, p2_u3167, p2_u3166, p2_u3165, p2_u3164, p2_u3163,
p2_u3162, p2_u3161, p2_u3160, p2_u3159, p2_u3158, p2_u3157, p2_u3156,
p2_u3155, p2_u3154, p2_u3153, p2_u3152, p2_u3151, p2_u3150, p2_u3149,
p2_u3148, p2_u3147, p2_u3146, p2_u3145, p2_u3144, p2_u3143, p2_u3142,
p2_u3141, p2_u3140, p2_u3139, p2_u3138, p2_u3137, p2_u3136, p2_u3135,
p2_u3134, p2_u3133, p2_u3132, p2_u3131, p2_u3130, p2_u3129, p2_u3128,
p2_u3127, p2_u3126, p2_u3125, p2_u3124, p2_u3123, p2_u3122, p2_u3121,
p2_u3120, p2_u3119, p2_u3118, p2_u3117, p2_u3116, p2_u3115, p2_u3114,
p2_u3113, p2_u3112, p2_u3111, p2_u3110, p2_u3109, p2_u3108, p2_u3107,
p2_u3106, p2_u3105, p2_u3104, p2_u3103, p2_u3102, p2_u3101, p2_u3100,
p2_u3099, p2_u3098, p2_u3097, p2_u3096, p2_u3095, p2_u3094, p2_u3093,
p2_u3092, p2_u3091, p2_u3090, p2_u3089, p2_u3088, p2_u3087, p2_u3086,
p2_u3085, p2_u3084, p2_u3083, p2_u3082, p2_u3081, p2_u3080, p2_u3079,
p2_u3078, p2_u3077, p2_u3076, p2_u3075, p2_u3074, p2_u3073, p2_u3072,
p2_u3071, p2_u3070, p2_u3069, p2_u3068, p2_u3067, p2_u3066, p2_u3065,
p2_u3064, p2_u3063, p2_u3062, p2_u3061, p2_u3060, p2_u3059, p2_u3058,
p2_u3057, p2_u3056, p2_u3055, p2_u3054, p2_u3053, p2_u3052, p2_u3051,
p2_u3050, p2_u3049, p2_u3048, p2_u3595, p2_u3596, p2_u3599, p2_u3600,
p2_u3601, p2_u3047, p2_u3602, p2_u3603, p2_u3604, p2_u3605, p2_u3046,
p2_u3045, p2_u3044, p2_u3043, p2_u3042, p2_u3041, p2_u3040, p2_u3039,
p2_u3038, p2_u3037, p2_u3036, p2_u3035, p2_u3034, p2_u3033, p2_u3032,
p2_u3031, p2_u3030, p2_u3029, p2_u3028, p2_u3027, p2_u3026, p2_u3025,
p2_u3024, p2_u3023, p2_u3022, p2_u3021, p2_u3020, p2_u3019, p2_u3018,
p2_u3017, p2_u3016, p2_u3015, p2_u3014, p2_u3013, p2_u3012, p2_u3011,
p2_u3010, p2_u3009, p2_u3008, p2_u3007, p2_u3006, p2_u3005, p2_u3004,
p2_u3003, p2_u3002, p2_u3001, p2_u3000, p2_u2999, p2_u2998, p2_u2997,
p2_u2996, p2_u2995, p2_u2994, p2_u2993, p2_u2992, p2_u2991, p2_u2990,
p2_u2989, p2_u2988, p2_u2987, p2_u2986, p2_u2985, p2_u2984, p2_u2983,
p2_u2982, p2_u2981, p2_u2980, p2_u2979, p2_u2978, p2_u2977, p2_u2976,
p2_u2975, p2_u2974, p2_u2973, p2_u2972, p2_u2971, p2_u2970, p2_u2969,
p2_u2968, p2_u2967, p2_u2966, p2_u2965, p2_u2964, p2_u2963, p2_u2962,
p2_u2961, p2_u2960, p2_u2959, p2_u2958, p2_u2957, p2_u2956, p2_u2955,
p2_u2954, p2_u2953, p2_u2952, p2_u2951, p2_u2950, p2_u2949, p2_u2948,
p2_u2947, p2_u2946, p2_u2945, p2_u2944, p2_u2943, p2_u2942, p2_u2941,
p2_u2940, p2_u2939, p2_u2938, p2_u2937, p2_u2936, p2_u2935, p2_u2934,
p2_u2933, p2_u2932, p2_u2931, p2_u2930, p2_u2929, p2_u2928, p2_u2927,
p2_u2926, p2_u2925, p2_u2924, p2_u2923, p2_u2922, p2_u2921, p2_u2920,
p2_u2919, p2_u2918, p2_u2917, p2_u2916, p2_u2915, p2_u2914, p2_u2913,
p2_u2912, p2_u2911, p2_u2910, p2_u2909, p2_u2908, p2_u2907, p2_u2906,
p2_u2905, p2_u2904, p2_u2903, p2_u2902, p2_u2901, p2_u2900, p2_u2899,
p2_u2898, p2_u2897, p2_u2896, p2_u2895, p2_u2894, p2_u2893, p2_u2892,
p2_u2891, p2_u2890, p2_u2889, p2_u2888, p2_u2887, p2_u2886, p2_u2885,
p2_u2884, p2_u2883, p2_u2882, p2_u2881, p2_u2880, p2_u2879, p2_u2878,
p2_u2877, p2_u2876, p2_u2875, p2_u2874, p2_u2873, p2_u2872, p2_u2871,
p2_u2870, p2_u2869, p2_u2868, p2_u2867, p2_u2866, p2_u2865, p2_u2864,
p2_u2863, p2_u2862, p2_u2861, p2_u2860, p2_u2859, p2_u2858, p2_u2857,
p2_u2856, p2_u2855, p2_u2854, p2_u2853, p2_u2852, p2_u2851, p2_u2850,
p2_u2849, p2_u2848, p2_u2847, p2_u2846, p2_u2845, p2_u2844, p2_u2843,
p2_u2842, p2_u2841, p2_u2840, p2_u2839, p2_u2838, p2_u2837, p2_u2836,
p2_u2835, p2_u2834, p2_u2833, p2_u2832, p2_u2831, p2_u2830, p2_u2829,
p2_u2828, p2_u2827, p2_u2826, p2_u2825, p2_u2824, p2_u2823, p2_u2822,
p2_u2821, p2_u2820, p2_u3608, p2_u2819, p2_u3609, p2_u2818, p2_u3610,
p2_u2817, p2_u3611, p2_u2816, p2_u2815, p2_u3612, p2_u2814, p1_u3458,
p1_u3459, p1_u3460, p1_u3461, p1_u3226, p1_u3225, p1_u3224, p1_u3223,
p1_u3222, p1_u3221, p1_u3220, p1_u3219, p1_u3218, p1_u3217, p1_u3216,
p1_u3215, p1_u3214, p1_u3213, p1_u3212, p1_u3211, p1_u3210, p1_u3209,
p1_u3208, p1_u3207, p1_u3206, p1_u3205, p1_u3204, p1_u3203, p1_u3202,
p1_u3201, p1_u3200, p1_u3199, p1_u3198, p1_u3197, p1_u3196, p1_u3195,
p1_u3194, p1_u3464, p1_u3465, p1_u3193, p1_u3192, p1_u3191, p1_u3190,
p1_u3189, p1_u3188, p1_u3187, p1_u3186, p1_u3185, p1_u3184, p1_u3183,
p1_u3182, p1_u3181, p1_u3180, p1_u3179, p1_u3178, p1_u3177, p1_u3176,
p1_u3175, p1_u3174, p1_u3173, p1_u3172, p1_u3171, p1_u3170, p1_u3169,
p1_u3168, p1_u3167, p1_u3166, p1_u3165, p1_u3164, p1_u3466, p1_u3163,
p1_u3162, p1_u3161, p1_u3160, p1_u3159, p1_u3158, p1_u3157, p1_u3156,
p1_u3155, p1_u3154, p1_u3153, p1_u3152, p1_u3151, p1_u3150, p1_u3149,
p1_u3148, p1_u3147, p1_u3146, p1_u3145, p1_u3144, p1_u3143, p1_u3142,
p1_u3141, p1_u3140, p1_u3139, p1_u3138, p1_u3137, p1_u3136, p1_u3135,
p1_u3134, p1_u3133, p1_u3132, p1_u3131, p1_u3130, p1_u3129, p1_u3128,
p1_u3127, p1_u3126, p1_u3125, p1_u3124, p1_u3123, p1_u3122, p1_u3121,
p1_u3120, p1_u3119, p1_u3118, p1_u3117, p1_u3116, p1_u3115, p1_u3114,
p1_u3113, p1_u3112, p1_u3111, p1_u3110, p1_u3109, p1_u3108, p1_u3107,
p1_u3106, p1_u3105, p1_u3104, p1_u3103, p1_u3102, p1_u3101, p1_u3100,
p1_u3099, p1_u3098, p1_u3097, p1_u3096, p1_u3095, p1_u3094, p1_u3093,
p1_u3092, p1_u3091, p1_u3090, p1_u3089, p1_u3088, p1_u3087, p1_u3086,
p1_u3085, p1_u3084, p1_u3083, p1_u3082, p1_u3081, p1_u3080, p1_u3079,
p1_u3078, p1_u3077, p1_u3076, p1_u3075, p1_u3074, p1_u3073, p1_u3072,
p1_u3071, p1_u3070, p1_u3069, p1_u3068, p1_u3067, p1_u3066, p1_u3065,
p1_u3064, p1_u3063, p1_u3062, p1_u3061, p1_u3060, p1_u3059, p1_u3058,
p1_u3057, p1_u3056, p1_u3055, p1_u3054, p1_u3053, p1_u3052, p1_u3051,
p1_u3050, p1_u3049, p1_u3048, p1_u3047, p1_u3046, p1_u3045, p1_u3044,
p1_u3043, p1_u3042, p1_u3041, p1_u3040, p1_u3039, p1_u3038, p1_u3037,
p1_u3036, p1_u3035, p1_u3034, p1_u3033, p1_u3468, p1_u3469, p1_u3472,
p1_u3473, p1_u3474, p1_u3032, p1_u3475, p1_u3476, p1_u3477, p1_u3478,
p1_u3031, p1_u3030, p1_u3029, p1_u3028, p1_u3027, p1_u3026, p1_u3025,
p1_u3024, p1_u3023, p1_u3022, p1_u3021, p1_u3020, p1_u3019, p1_u3018,
p1_u3017, p1_u3016, p1_u3015, p1_u3014, p1_u3013, p1_u3012, p1_u3011,
p1_u3010, p1_u3009, p1_u3008, p1_u3007, p1_u3006, p1_u3005, p1_u3004,
p1_u3003, p1_u3002, p1_u3001, p1_u3000, p1_u2999, p1_u2998, p1_u2997,
p1_u2996, p1_u2995, p1_u2994, p1_u2993, p1_u2992, p1_u2991, p1_u2990,
p1_u2989, p1_u2988, p1_u2987, p1_u2986, p1_u2985, p1_u2984, p1_u2983,
p1_u2982, p1_u2981, p1_u2980, p1_u2979, p1_u2978, p1_u2977, p1_u2976,
p1_u2975, p1_u2974, p1_u2973, p1_u2972, p1_u2971, p1_u2970, p1_u2969,
p1_u2968, p1_u2967, p1_u2966, p1_u2965, p1_u2964, p1_u2963, p1_u2962,
p1_u2961, p1_u2960, p1_u2959, p1_u2958, p1_u2957, p1_u2956, p1_u2955,
p1_u2954, p1_u2953, p1_u2952, p1_u2951, p1_u2950, p1_u2949, p1_u2948,
p1_u2947, p1_u2946, p1_u2945, p1_u2944, p1_u2943, p1_u2942, p1_u2941,
p1_u2940, p1_u2939, p1_u2938, p1_u2937, p1_u2936, p1_u2935, p1_u2934,
p1_u2933, p1_u2932, p1_u2931, p1_u2930, p1_u2929, p1_u2928, p1_u2927,
p1_u2926, p1_u2925, p1_u2924, p1_u2923, p1_u2922, p1_u2921, p1_u2920,
p1_u2919, p1_u2918, p1_u2917, p1_u2916, p1_u2915, p1_u2914, p1_u2913,
p1_u2912, p1_u2911, p1_u2910, p1_u2909, p1_u2908, p1_u2907, p1_u2906,
p1_u2905, p1_u2904, p1_u2903, p1_u2902, p1_u2901, p1_u2900, p1_u2899,
p1_u2898, p1_u2897, p1_u2896, p1_u2895, p1_u2894, p1_u2893, p1_u2892,
p1_u2891, p1_u2890, p1_u2889, p1_u2888, p1_u2887, p1_u2886, p1_u2885,
p1_u2884, p1_u2883, p1_u2882, p1_u2881, p1_u2880, p1_u2879, p1_u2878,
p1_u2877, p1_u2876, p1_u2875, p1_u2874, p1_u2873, p1_u2872, p1_u2871,
p1_u2870, p1_u2869, p1_u2868, p1_u2867, p1_u2866, p1_u2865, p1_u2864,
p1_u2863, p1_u2862, p1_u2861, p1_u2860, p1_u2859, p1_u2858, p1_u2857,
p1_u2856, p1_u2855, p1_u2854, p1_u2853, p1_u2852, p1_u2851, p1_u2850,
p1_u2849, p1_u2848, p1_u2847, p1_u2846, p1_u2845, p1_u2844, p1_u2843,
p1_u2842, p1_u2841, p1_u2840, p1_u2839, p1_u2838, p1_u2837, p1_u2836,
p1_u2835, p1_u2834, p1_u2833, p1_u2832, p1_u2831, p1_u2830, p1_u2829,
p1_u2828, p1_u2827, p1_u2826, p1_u2825, p1_u2824, p1_u2823, p1_u2822,
p1_u2821, p1_u2820, p1_u2819, p1_u2818, p1_u2817, p1_u2816, p1_u2815,
p1_u2814, p1_u2813, p1_u2812, p1_u2811, p1_u2810, p1_u2809, p1_u2808,
p1_u3481, p1_u2807, p1_u3482, p1_u3483, p1_u2806, p1_u3484, p1_u2805,
p1_u3485, p1_u2804, p1_u3486, p1_u2803, p1_u2802, p1_u3487, p1_u2801
);
input datai_31_, datai_30_, datai_29_, datai_28_, datai_27_, datai_26_,
datai_25_, datai_24_, datai_23_, datai_22_, datai_21_, datai_20_,
datai_19_, datai_18_, datai_17_, datai_16_, datai_15_, datai_14_,
datai_13_, datai_12_, datai_11_, datai_10_, datai_9_, datai_8_,
datai_7_, datai_6_, datai_5_, datai_4_, datai_3_, datai_2_, datai_1_,
datai_0_, hold, na, bs16, ready1, ready2, buf1_reg_0_, buf1_reg_1_,
buf1_reg_2_, buf1_reg_3_, buf1_reg_4_, buf1_reg_5_, buf1_reg_6_,
buf1_reg_7_, buf1_reg_8_, buf1_reg_9_, buf1_reg_10_, buf1_reg_11_,
buf1_reg_12_, buf1_reg_13_, buf1_reg_14_, buf1_reg_15_, buf1_reg_16_,
buf1_reg_17_, buf1_reg_18_, buf1_reg_19_, buf1_reg_20_, buf1_reg_21_,
buf1_reg_22_, buf1_reg_23_, buf1_reg_24_, buf1_reg_25_, buf1_reg_26_,
buf1_reg_27_, buf1_reg_28_, buf1_reg_29_, buf1_reg_30_, buf1_reg_31_,
buf2_reg_0_, buf2_reg_1_, buf2_reg_2_, buf2_reg_3_, buf2_reg_4_,
buf2_reg_5_, buf2_reg_6_, buf2_reg_7_, buf2_reg_8_, buf2_reg_9_,
buf2_reg_10_, buf2_reg_11_, buf2_reg_12_, buf2_reg_13_, buf2_reg_14_,
buf2_reg_15_, buf2_reg_16_, buf2_reg_17_, buf2_reg_18_, buf2_reg_19_,
buf2_reg_20_, buf2_reg_21_, buf2_reg_22_, buf2_reg_23_, buf2_reg_24_,
buf2_reg_25_, buf2_reg_26_, buf2_reg_27_, buf2_reg_28_, buf2_reg_29_,
buf2_reg_30_, buf2_reg_31_, ready12_reg, ready21_reg, ready22_reg,
ready11_reg, p3_be_n_reg_3_, p3_be_n_reg_2_, p3_be_n_reg_1_,
p3_be_n_reg_0_, p3_address_reg_29_, p3_address_reg_28_,
p3_address_reg_27_, p3_address_reg_26_, p3_address_reg_25_,
p3_address_reg_24_, p3_address_reg_23_, p3_address_reg_22_,
p3_address_reg_21_, p3_address_reg_20_, p3_address_reg_19_,
p3_address_reg_18_, p3_address_reg_17_, p3_address_reg_16_,
p3_address_reg_15_, p3_address_reg_14_, p3_address_reg_13_,
p3_address_reg_12_, p3_address_reg_11_, p3_address_reg_10_,
p3_address_reg_9_, p3_address_reg_8_, p3_address_reg_7_,
p3_address_reg_6_, p3_address_reg_5_, p3_address_reg_4_,
p3_address_reg_3_, p3_address_reg_2_, p3_address_reg_1_,
p3_address_reg_0_, p3_state_reg_2_, p3_state_reg_1_, p3_state_reg_0_,
p3_datawidth_reg_0_, p3_datawidth_reg_1_, p3_datawidth_reg_2_,
p3_datawidth_reg_3_, p3_datawidth_reg_4_, p3_datawidth_reg_5_,
p3_datawidth_reg_6_, p3_datawidth_reg_7_, p3_datawidth_reg_8_,
p3_datawidth_reg_9_, p3_datawidth_reg_10_, p3_datawidth_reg_11_,
p3_datawidth_reg_12_, p3_datawidth_reg_13_, p3_datawidth_reg_14_,
p3_datawidth_reg_15_, p3_datawidth_reg_16_, p3_datawidth_reg_17_,
p3_datawidth_reg_18_, p3_datawidth_reg_19_, p3_datawidth_reg_20_,
p3_datawidth_reg_21_, p3_datawidth_reg_22_, p3_datawidth_reg_23_,
p3_datawidth_reg_24_, p3_datawidth_reg_25_, p3_datawidth_reg_26_,
p3_datawidth_reg_27_, p3_datawidth_reg_28_, p3_datawidth_reg_29_,
p3_datawidth_reg_30_, p3_datawidth_reg_31_, p3_state2_reg_3_,
p3_state2_reg_2_, p3_state2_reg_1_, p3_state2_reg_0_,
p3_instqueue_reg_15__7_, p3_instqueue_reg_15__6_,
p3_instqueue_reg_15__5_, p3_instqueue_reg_15__4_,
p3_instqueue_reg_15__3_, p3_instqueue_reg_15__2_,
p3_instqueue_reg_15__1_, p3_instqueue_reg_15__0_,
p3_instqueue_reg_14__7_, p3_instqueue_reg_14__6_,
p3_instqueue_reg_14__5_, p3_instqueue_reg_14__4_,
p3_instqueue_reg_14__3_, p3_instqueue_reg_14__2_,
p3_instqueue_reg_14__1_, p3_instqueue_reg_14__0_,
p3_instqueue_reg_13__7_, p3_instqueue_reg_13__6_,
p3_instqueue_reg_13__5_, p3_instqueue_reg_13__4_,
p3_instqueue_reg_13__3_, p3_instqueue_reg_13__2_,
p3_instqueue_reg_13__1_, p3_instqueue_reg_13__0_,
p3_instqueue_reg_12__7_, p3_instqueue_reg_12__6_,
p3_instqueue_reg_12__5_, p3_instqueue_reg_12__4_,
p3_instqueue_reg_12__3_, p3_instqueue_reg_12__2_,
p3_instqueue_reg_12__1_, p3_instqueue_reg_12__0_,
p3_instqueue_reg_11__7_, p3_instqueue_reg_11__6_,
p3_instqueue_reg_11__5_, p3_instqueue_reg_11__4_,
p3_instqueue_reg_11__3_, p3_instqueue_reg_11__2_,
p3_instqueue_reg_11__1_, p3_instqueue_reg_11__0_,
p3_instqueue_reg_10__7_, p3_instqueue_reg_10__6_,
p3_instqueue_reg_10__5_, p3_instqueue_reg_10__4_,
p3_instqueue_reg_10__3_, p3_instqueue_reg_10__2_,
p3_instqueue_reg_10__1_, p3_instqueue_reg_10__0_,
p3_instqueue_reg_9__7_, p3_instqueue_reg_9__6_,
p3_instqueue_reg_9__5_, p3_instqueue_reg_9__4_,
p3_instqueue_reg_9__3_, p3_instqueue_reg_9__2_,
p3_instqueue_reg_9__1_, p3_instqueue_reg_9__0_,
p3_instqueue_reg_8__7_, p3_instqueue_reg_8__6_,
p3_instqueue_reg_8__5_, p3_instqueue_reg_8__4_,
p3_instqueue_reg_8__3_, p3_instqueue_reg_8__2_,
p3_instqueue_reg_8__1_, p3_instqueue_reg_8__0_,
p3_instqueue_reg_7__7_, p3_instqueue_reg_7__6_,
p3_instqueue_reg_7__5_, p3_instqueue_reg_7__4_,
p3_instqueue_reg_7__3_, p3_instqueue_reg_7__2_,
p3_instqueue_reg_7__1_, p3_instqueue_reg_7__0_,
p3_instqueue_reg_6__7_, p3_instqueue_reg_6__6_,
p3_instqueue_reg_6__5_, p3_instqueue_reg_6__4_,
p3_instqueue_reg_6__3_, p3_instqueue_reg_6__2_,
p3_instqueue_reg_6__1_, p3_instqueue_reg_6__0_,
p3_instqueue_reg_5__7_, p3_instqueue_reg_5__6_,
p3_instqueue_reg_5__5_, p3_instqueue_reg_5__4_,
p3_instqueue_reg_5__3_, p3_instqueue_reg_5__2_,
p3_instqueue_reg_5__1_, p3_instqueue_reg_5__0_,
p3_instqueue_reg_4__7_, p3_instqueue_reg_4__6_,
p3_instqueue_reg_4__5_, p3_instqueue_reg_4__4_,
p3_instqueue_reg_4__3_, p3_instqueue_reg_4__2_,
p3_instqueue_reg_4__1_, p3_instqueue_reg_4__0_,
p3_instqueue_reg_3__7_, p3_instqueue_reg_3__6_,
p3_instqueue_reg_3__5_, p3_instqueue_reg_3__4_,
p3_instqueue_reg_3__3_, p3_instqueue_reg_3__2_,
p3_instqueue_reg_3__1_, p3_instqueue_reg_3__0_,
p3_instqueue_reg_2__7_, p3_instqueue_reg_2__6_,
p3_instqueue_reg_2__5_, p3_instqueue_reg_2__4_,
p3_instqueue_reg_2__3_, p3_instqueue_reg_2__2_,
p3_instqueue_reg_2__1_, p3_instqueue_reg_2__0_,
p3_instqueue_reg_1__7_, p3_instqueue_reg_1__6_,
p3_instqueue_reg_1__5_, p3_instqueue_reg_1__4_,
p3_instqueue_reg_1__3_, p3_instqueue_reg_1__2_,
p3_instqueue_reg_1__1_, p3_instqueue_reg_1__0_,
p3_instqueue_reg_0__7_, p3_instqueue_reg_0__6_,
p3_instqueue_reg_0__5_, p3_instqueue_reg_0__4_,
p3_instqueue_reg_0__3_, p3_instqueue_reg_0__2_,
p3_instqueue_reg_0__1_, p3_instqueue_reg_0__0_,
p3_instqueuerd_addr_reg_4_, p3_instqueuerd_addr_reg_3_,
p3_instqueuerd_addr_reg_2_, p3_instqueuerd_addr_reg_1_,
p3_instqueuerd_addr_reg_0_, p3_instqueuewr_addr_reg_4_,
p3_instqueuewr_addr_reg_3_, p3_instqueuewr_addr_reg_2_,
p3_instqueuewr_addr_reg_1_, p3_instqueuewr_addr_reg_0_,
p3_instaddrpointer_reg_0_, p3_instaddrpointer_reg_1_,
p3_instaddrpointer_reg_2_, p3_instaddrpointer_reg_3_,
p3_instaddrpointer_reg_4_, p3_instaddrpointer_reg_5_,
p3_instaddrpointer_reg_6_, p3_instaddrpointer_reg_7_,
p3_instaddrpointer_reg_8_, p3_instaddrpointer_reg_9_,
p3_instaddrpointer_reg_10_, p3_instaddrpointer_reg_11_,
p3_instaddrpointer_reg_12_, p3_instaddrpointer_reg_13_,
p3_instaddrpointer_reg_14_, p3_instaddrpointer_reg_15_,
p3_instaddrpointer_reg_16_, p3_instaddrpointer_reg_17_,
p3_instaddrpointer_reg_18_, p3_instaddrpointer_reg_19_,
p3_instaddrpointer_reg_20_, p3_instaddrpointer_reg_21_,
p3_instaddrpointer_reg_22_, p3_instaddrpointer_reg_23_,
p3_instaddrpointer_reg_24_, p3_instaddrpointer_reg_25_,
p3_instaddrpointer_reg_26_, p3_instaddrpointer_reg_27_,
p3_instaddrpointer_reg_28_, p3_instaddrpointer_reg_29_,
p3_instaddrpointer_reg_30_, p3_instaddrpointer_reg_31_,
p3_phyaddrpointer_reg_0_, p3_phyaddrpointer_reg_1_,
p3_phyaddrpointer_reg_2_, p3_phyaddrpointer_reg_3_,
p3_phyaddrpointer_reg_4_, p3_phyaddrpointer_reg_5_,
p3_phyaddrpointer_reg_6_, p3_phyaddrpointer_reg_7_,
p3_phyaddrpointer_reg_8_, p3_phyaddrpointer_reg_9_,
p3_phyaddrpointer_reg_10_, p3_phyaddrpointer_reg_11_,
p3_phyaddrpointer_reg_12_, p3_phyaddrpointer_reg_13_,
p3_phyaddrpointer_reg_14_, p3_phyaddrpointer_reg_15_,
p3_phyaddrpointer_reg_16_, p3_phyaddrpointer_reg_17_,
p3_phyaddrpointer_reg_18_, p3_phyaddrpointer_reg_19_,
p3_phyaddrpointer_reg_20_, p3_phyaddrpointer_reg_21_,
p3_phyaddrpointer_reg_22_, p3_phyaddrpointer_reg_23_,
p3_phyaddrpointer_reg_24_, p3_phyaddrpointer_reg_25_,
p3_phyaddrpointer_reg_26_, p3_phyaddrpointer_reg_27_,
p3_phyaddrpointer_reg_28_, p3_phyaddrpointer_reg_29_,
p3_phyaddrpointer_reg_30_, p3_phyaddrpointer_reg_31_,
p3_lword_reg_15_, p3_lword_reg_14_, p3_lword_reg_13_,
p3_lword_reg_12_, p3_lword_reg_11_, p3_lword_reg_10_, p3_lword_reg_9_,
p3_lword_reg_8_, p3_lword_reg_7_, p3_lword_reg_6_, p3_lword_reg_5_,
p3_lword_reg_4_, p3_lword_reg_3_, p3_lword_reg_2_, p3_lword_reg_1_,
p3_lword_reg_0_, p3_uword_reg_14_, p3_uword_reg_13_, p3_uword_reg_12_,
p3_uword_reg_11_, p3_uword_reg_10_, p3_uword_reg_9_, p3_uword_reg_8_,
p3_uword_reg_7_, p3_uword_reg_6_, p3_uword_reg_5_, p3_uword_reg_4_,
p3_uword_reg_3_, p3_uword_reg_2_, p3_uword_reg_1_, p3_uword_reg_0_,
p3_datao_reg_0_, p3_datao_reg_1_, p3_datao_reg_2_, p3_datao_reg_3_,
p3_datao_reg_4_, p3_datao_reg_5_, p3_datao_reg_6_, p3_datao_reg_7_,
p3_datao_reg_8_, p3_datao_reg_9_, p3_datao_reg_10_, p3_datao_reg_11_,
p3_datao_reg_12_, p3_datao_reg_13_, p3_datao_reg_14_,
p3_datao_reg_15_, p3_datao_reg_16_, p3_datao_reg_17_,
p3_datao_reg_18_, p3_datao_reg_19_, p3_datao_reg_20_,
p3_datao_reg_21_, p3_datao_reg_22_, p3_datao_reg_23_,
p3_datao_reg_24_, p3_datao_reg_25_, p3_datao_reg_26_,
p3_datao_reg_27_, p3_datao_reg_28_, p3_datao_reg_29_,
p3_datao_reg_30_, p3_datao_reg_31_, p3_eax_reg_0_, p3_eax_reg_1_,
p3_eax_reg_2_, p3_eax_reg_3_, p3_eax_reg_4_, p3_eax_reg_5_,
p3_eax_reg_6_, p3_eax_reg_7_, p3_eax_reg_8_, p3_eax_reg_9_,
p3_eax_reg_10_, p3_eax_reg_11_, p3_eax_reg_12_, p3_eax_reg_13_,
p3_eax_reg_14_, p3_eax_reg_15_, p3_eax_reg_16_, p3_eax_reg_17_,
p3_eax_reg_18_, p3_eax_reg_19_, p3_eax_reg_20_, p3_eax_reg_21_,
p3_eax_reg_22_, p3_eax_reg_23_, p3_eax_reg_24_, p3_eax_reg_25_,
p3_eax_reg_26_, p3_eax_reg_27_, p3_eax_reg_28_, p3_eax_reg_29_,
p3_eax_reg_30_, p3_eax_reg_31_, p3_ebx_reg_0_, p3_ebx_reg_1_,
p3_ebx_reg_2_, p3_ebx_reg_3_, p3_ebx_reg_4_, p3_ebx_reg_5_,
p3_ebx_reg_6_, p3_ebx_reg_7_, p3_ebx_reg_8_, p3_ebx_reg_9_,
p3_ebx_reg_10_, p3_ebx_reg_11_, p3_ebx_reg_12_, p3_ebx_reg_13_,
p3_ebx_reg_14_, p3_ebx_reg_15_, p3_ebx_reg_16_, p3_ebx_reg_17_,
p3_ebx_reg_18_, p3_ebx_reg_19_, p3_ebx_reg_20_, p3_ebx_reg_21_,
p3_ebx_reg_22_, p3_ebx_reg_23_, p3_ebx_reg_24_, p3_ebx_reg_25_,
p3_ebx_reg_26_, p3_ebx_reg_27_, p3_ebx_reg_28_, p3_ebx_reg_29_,
p3_ebx_reg_30_, p3_ebx_reg_31_, p3_reip_reg_0_, p3_reip_reg_1_,
p3_reip_reg_2_, p3_reip_reg_3_, p3_reip_reg_4_, p3_reip_reg_5_,
p3_reip_reg_6_, p3_reip_reg_7_, p3_reip_reg_8_, p3_reip_reg_9_,
p3_reip_reg_10_, p3_reip_reg_11_, p3_reip_reg_12_, p3_reip_reg_13_,
p3_reip_reg_14_, p3_reip_reg_15_, p3_reip_reg_16_, p3_reip_reg_17_,
p3_reip_reg_18_, p3_reip_reg_19_, p3_reip_reg_20_, p3_reip_reg_21_,
p3_reip_reg_22_, p3_reip_reg_23_, p3_reip_reg_24_, p3_reip_reg_25_,
p3_reip_reg_26_, p3_reip_reg_27_, p3_reip_reg_28_, p3_reip_reg_29_,
p3_reip_reg_30_, p3_reip_reg_31_, p3_byteenable_reg_3_,
p3_byteenable_reg_2_, p3_byteenable_reg_1_, p3_byteenable_reg_0_,
p3_w_r_n_reg, p3_flush_reg, p3_more_reg, p3_statebs16_reg,
p3_requestpending_reg, p3_d_c_n_reg, p3_m_io_n_reg, p3_codefetch_reg,
p3_ads_n_reg, p3_readrequest_reg, p3_memoryfetch_reg, p2_be_n_reg_3_,
p2_be_n_reg_2_, p2_be_n_reg_1_, p2_be_n_reg_0_, p2_address_reg_29_,
p2_address_reg_28_, p2_address_reg_27_, p2_address_reg_26_,
p2_address_reg_25_, p2_address_reg_24_, p2_address_reg_23_,
p2_address_reg_22_, p2_address_reg_21_, p2_address_reg_20_,
p2_address_reg_19_, p2_address_reg_18_, p2_address_reg_17_,
p2_address_reg_16_, p2_address_reg_15_, p2_address_reg_14_,
p2_address_reg_13_, p2_address_reg_12_, p2_address_reg_11_,
p2_address_reg_10_, p2_address_reg_9_, p2_address_reg_8_,
p2_address_reg_7_, p2_address_reg_6_, p2_address_reg_5_,
p2_address_reg_4_, p2_address_reg_3_, p2_address_reg_2_,
p2_address_reg_1_, p2_address_reg_0_, p2_state_reg_2_,
p2_state_reg_1_, p2_state_reg_0_, p2_datawidth_reg_0_,
p2_datawidth_reg_1_, p2_datawidth_reg_2_, p2_datawidth_reg_3_,
p2_datawidth_reg_4_, p2_datawidth_reg_5_, p2_datawidth_reg_6_,
p2_datawidth_reg_7_, p2_datawidth_reg_8_, p2_datawidth_reg_9_,
p2_datawidth_reg_10_, p2_datawidth_reg_11_, p2_datawidth_reg_12_,
p2_datawidth_reg_13_, p2_datawidth_reg_14_, p2_datawidth_reg_15_,
p2_datawidth_reg_16_, p2_datawidth_reg_17_, p2_datawidth_reg_18_,
p2_datawidth_reg_19_, p2_datawidth_reg_20_, p2_datawidth_reg_21_,
p2_datawidth_reg_22_, p2_datawidth_reg_23_, p2_datawidth_reg_24_,
p2_datawidth_reg_25_, p2_datawidth_reg_26_, p2_datawidth_reg_27_,
p2_datawidth_reg_28_, p2_datawidth_reg_29_, p2_datawidth_reg_30_,
p2_datawidth_reg_31_, p2_state2_reg_3_, p2_state2_reg_2_,
p2_state2_reg_1_, p2_state2_reg_0_, p2_instqueue_reg_15__7_,
p2_instqueue_reg_15__6_, p2_instqueue_reg_15__5_,
p2_instqueue_reg_15__4_, p2_instqueue_reg_15__3_,
p2_instqueue_reg_15__2_, p2_instqueue_reg_15__1_,
p2_instqueue_reg_15__0_, p2_instqueue_reg_14__7_,
p2_instqueue_reg_14__6_, p2_instqueue_reg_14__5_,
p2_instqueue_reg_14__4_, p2_instqueue_reg_14__3_,
p2_instqueue_reg_14__2_, p2_instqueue_reg_14__1_,
p2_instqueue_reg_14__0_, p2_instqueue_reg_13__7_,
p2_instqueue_reg_13__6_, p2_instqueue_reg_13__5_,
p2_instqueue_reg_13__4_, p2_instqueue_reg_13__3_,
p2_instqueue_reg_13__2_, p2_instqueue_reg_13__1_,
p2_instqueue_reg_13__0_, p2_instqueue_reg_12__7_,
p2_instqueue_reg_12__6_, p2_instqueue_reg_12__5_,
p2_instqueue_reg_12__4_, p2_instqueue_reg_12__3_,
p2_instqueue_reg_12__2_, p2_instqueue_reg_12__1_,
p2_instqueue_reg_12__0_, p2_instqueue_reg_11__7_,
p2_instqueue_reg_11__6_, p2_instqueue_reg_11__5_,
p2_instqueue_reg_11__4_, p2_instqueue_reg_11__3_,
p2_instqueue_reg_11__2_, p2_instqueue_reg_11__1_,
p2_instqueue_reg_11__0_, p2_instqueue_reg_10__7_,
p2_instqueue_reg_10__6_, p2_instqueue_reg_10__5_,
p2_instqueue_reg_10__4_, p2_instqueue_reg_10__3_,
p2_instqueue_reg_10__2_, p2_instqueue_reg_10__1_,
p2_instqueue_reg_10__0_, p2_instqueue_reg_9__7_,
p2_instqueue_reg_9__6_, p2_instqueue_reg_9__5_,
p2_instqueue_reg_9__4_, p2_instqueue_reg_9__3_,
p2_instqueue_reg_9__2_, p2_instqueue_reg_9__1_,
p2_instqueue_reg_9__0_, p2_instqueue_reg_8__7_,
p2_instqueue_reg_8__6_, p2_instqueue_reg_8__5_,
p2_instqueue_reg_8__4_, p2_instqueue_reg_8__3_,
p2_instqueue_reg_8__2_, p2_instqueue_reg_8__1_,
p2_instqueue_reg_8__0_, p2_instqueue_reg_7__7_,
p2_instqueue_reg_7__6_, p2_instqueue_reg_7__5_,
p2_instqueue_reg_7__4_, p2_instqueue_reg_7__3_,
p2_instqueue_reg_7__2_, p2_instqueue_reg_7__1_,
p2_instqueue_reg_7__0_, p2_instqueue_reg_6__7_,
p2_instqueue_reg_6__6_, p2_instqueue_reg_6__5_,
p2_instqueue_reg_6__4_, p2_instqueue_reg_6__3_,
p2_instqueue_reg_6__2_, p2_instqueue_reg_6__1_,
p2_instqueue_reg_6__0_, p2_instqueue_reg_5__7_,
p2_instqueue_reg_5__6_, p2_instqueue_reg_5__5_,
p2_instqueue_reg_5__4_, p2_instqueue_reg_5__3_,
p2_instqueue_reg_5__2_, p2_instqueue_reg_5__1_,
p2_instqueue_reg_5__0_, p2_instqueue_reg_4__7_,
p2_instqueue_reg_4__6_, p2_instqueue_reg_4__5_,
p2_instqueue_reg_4__4_, p2_instqueue_reg_4__3_,
p2_instqueue_reg_4__2_, p2_instqueue_reg_4__1_,
p2_instqueue_reg_4__0_, p2_instqueue_reg_3__7_,
p2_instqueue_reg_3__6_, p2_instqueue_reg_3__5_,
p2_instqueue_reg_3__4_, p2_instqueue_reg_3__3_,
p2_instqueue_reg_3__2_, p2_instqueue_reg_3__1_,
p2_instqueue_reg_3__0_, p2_instqueue_reg_2__7_,
p2_instqueue_reg_2__6_, p2_instqueue_reg_2__5_,
p2_instqueue_reg_2__4_, p2_instqueue_reg_2__3_,
p2_instqueue_reg_2__2_, p2_instqueue_reg_2__1_,
p2_instqueue_reg_2__0_, p2_instqueue_reg_1__7_,
p2_instqueue_reg_1__6_, p2_instqueue_reg_1__5_,
p2_instqueue_reg_1__4_, p2_instqueue_reg_1__3_,
p2_instqueue_reg_1__2_, p2_instqueue_reg_1__1_,
p2_instqueue_reg_1__0_, p2_instqueue_reg_0__7_,
p2_instqueue_reg_0__6_, p2_instqueue_reg_0__5_,
p2_instqueue_reg_0__4_, p2_instqueue_reg_0__3_,
p2_instqueue_reg_0__2_, p2_instqueue_reg_0__1_,
p2_instqueue_reg_0__0_, p2_instqueuerd_addr_reg_4_,
p2_instqueuerd_addr_reg_3_, p2_instqueuerd_addr_reg_2_,
p2_instqueuerd_addr_reg_1_, p2_instqueuerd_addr_reg_0_,
p2_instqueuewr_addr_reg_4_, p2_instqueuewr_addr_reg_3_,
p2_instqueuewr_addr_reg_2_, p2_instqueuewr_addr_reg_1_,
p2_instqueuewr_addr_reg_0_, p2_instaddrpointer_reg_0_,
p2_instaddrpointer_reg_1_, p2_instaddrpointer_reg_2_,
p2_instaddrpointer_reg_3_, p2_instaddrpointer_reg_4_,
p2_instaddrpointer_reg_5_, p2_instaddrpointer_reg_6_,
p2_instaddrpointer_reg_7_, p2_instaddrpointer_reg_8_,
p2_instaddrpointer_reg_9_, p2_instaddrpointer_reg_10_,
p2_instaddrpointer_reg_11_, p2_instaddrpointer_reg_12_,
p2_instaddrpointer_reg_13_, p2_instaddrpointer_reg_14_,
p2_instaddrpointer_reg_15_, p2_instaddrpointer_reg_16_,
p2_instaddrpointer_reg_17_, p2_instaddrpointer_reg_18_,
p2_instaddrpointer_reg_19_, p2_instaddrpointer_reg_20_,
p2_instaddrpointer_reg_21_, p2_instaddrpointer_reg_22_,
p2_instaddrpointer_reg_23_, p2_instaddrpointer_reg_24_,
p2_instaddrpointer_reg_25_, p2_instaddrpointer_reg_26_,
p2_instaddrpointer_reg_27_, p2_instaddrpointer_reg_28_,
p2_instaddrpointer_reg_29_, p2_instaddrpointer_reg_30_,
p2_instaddrpointer_reg_31_, p2_phyaddrpointer_reg_0_,
p2_phyaddrpointer_reg_1_, p2_phyaddrpointer_reg_2_,
p2_phyaddrpointer_reg_3_, p2_phyaddrpointer_reg_4_,
p2_phyaddrpointer_reg_5_, p2_phyaddrpointer_reg_6_,
p2_phyaddrpointer_reg_7_, p2_phyaddrpointer_reg_8_,
p2_phyaddrpointer_reg_9_, p2_phyaddrpointer_reg_10_,
p2_phyaddrpointer_reg_11_, p2_phyaddrpointer_reg_12_,
p2_phyaddrpointer_reg_13_, p2_phyaddrpointer_reg_14_,
p2_phyaddrpointer_reg_15_, p2_phyaddrpointer_reg_16_,
p2_phyaddrpointer_reg_17_, p2_phyaddrpointer_reg_18_,
p2_phyaddrpointer_reg_19_, p2_phyaddrpointer_reg_20_,
p2_phyaddrpointer_reg_21_, p2_phyaddrpointer_reg_22_,
p2_phyaddrpointer_reg_23_, p2_phyaddrpointer_reg_24_,
p2_phyaddrpointer_reg_25_, p2_phyaddrpointer_reg_26_,
p2_phyaddrpointer_reg_27_, p2_phyaddrpointer_reg_28_,
p2_phyaddrpointer_reg_29_, p2_phyaddrpointer_reg_30_,
p2_phyaddrpointer_reg_31_, p2_lword_reg_15_, p2_lword_reg_14_,
p2_lword_reg_13_, p2_lword_reg_12_, p2_lword_reg_11_,
p2_lword_reg_10_, p2_lword_reg_9_, p2_lword_reg_8_, p2_lword_reg_7_,
p2_lword_reg_6_, p2_lword_reg_5_, p2_lword_reg_4_, p2_lword_reg_3_,
p2_lword_reg_2_, p2_lword_reg_1_, p2_lword_reg_0_, p2_uword_reg_14_,
p2_uword_reg_13_, p2_uword_reg_12_, p2_uword_reg_11_,
p2_uword_reg_10_, p2_uword_reg_9_, p2_uword_reg_8_, p2_uword_reg_7_,
p2_uword_reg_6_, p2_uword_reg_5_, p2_uword_reg_4_, p2_uword_reg_3_,
p2_uword_reg_2_, p2_uword_reg_1_, p2_uword_reg_0_, p2_datao_reg_0_,
p2_datao_reg_1_, p2_datao_reg_2_, p2_datao_reg_3_, p2_datao_reg_4_,
p2_datao_reg_5_, p2_datao_reg_6_, p2_datao_reg_7_, p2_datao_reg_8_,
p2_datao_reg_9_, p2_datao_reg_10_, p2_datao_reg_11_, p2_datao_reg_12_,
p2_datao_reg_13_, p2_datao_reg_14_, p2_datao_reg_15_,
p2_datao_reg_16_, p2_datao_reg_17_, p2_datao_reg_18_,
p2_datao_reg_19_, p2_datao_reg_20_, p2_datao_reg_21_,
p2_datao_reg_22_, p2_datao_reg_23_, p2_datao_reg_24_,
p2_datao_reg_25_, p2_datao_reg_26_, p2_datao_reg_27_,
p2_datao_reg_28_, p2_datao_reg_29_, p2_datao_reg_30_,
p2_datao_reg_31_, p2_eax_reg_0_, p2_eax_reg_1_, p2_eax_reg_2_,
p2_eax_reg_3_, p2_eax_reg_4_, p2_eax_reg_5_, p2_eax_reg_6_,
p2_eax_reg_7_, p2_eax_reg_8_, p2_eax_reg_9_, p2_eax_reg_10_,
p2_eax_reg_11_, p2_eax_reg_12_, p2_eax_reg_13_, p2_eax_reg_14_,
p2_eax_reg_15_, p2_eax_reg_16_, p2_eax_reg_17_, p2_eax_reg_18_,
p2_eax_reg_19_, p2_eax_reg_20_, p2_eax_reg_21_, p2_eax_reg_22_,
p2_eax_reg_23_, p2_eax_reg_24_, p2_eax_reg_25_, p2_eax_reg_26_,
p2_eax_reg_27_, p2_eax_reg_28_, p2_eax_reg_29_, p2_eax_reg_30_,
p2_eax_reg_31_, p2_ebx_reg_0_, p2_ebx_reg_1_, p2_ebx_reg_2_,
p2_ebx_reg_3_, p2_ebx_reg_4_, p2_ebx_reg_5_, p2_ebx_reg_6_,
p2_ebx_reg_7_, p2_ebx_reg_8_, p2_ebx_reg_9_, p2_ebx_reg_10_,
p2_ebx_reg_11_, p2_ebx_reg_12_, p2_ebx_reg_13_, p2_ebx_reg_14_,
p2_ebx_reg_15_, p2_ebx_reg_16_, p2_ebx_reg_17_, p2_ebx_reg_18_,
p2_ebx_reg_19_, p2_ebx_reg_20_, p2_ebx_reg_21_, p2_ebx_reg_22_,
p2_ebx_reg_23_, p2_ebx_reg_24_, p2_ebx_reg_25_, p2_ebx_reg_26_,
p2_ebx_reg_27_, p2_ebx_reg_28_, p2_ebx_reg_29_, p2_ebx_reg_30_,
p2_ebx_reg_31_, p2_reip_reg_0_, p2_reip_reg_1_, p2_reip_reg_2_,
p2_reip_reg_3_, p2_reip_reg_4_, p2_reip_reg_5_, p2_reip_reg_6_,
p2_reip_reg_7_, p2_reip_reg_8_, p2_reip_reg_9_, p2_reip_reg_10_,
p2_reip_reg_11_, p2_reip_reg_12_, p2_reip_reg_13_, p2_reip_reg_14_,
p2_reip_reg_15_, p2_reip_reg_16_, p2_reip_reg_17_, p2_reip_reg_18_,
p2_reip_reg_19_, p2_reip_reg_20_, p2_reip_reg_21_, p2_reip_reg_22_,
p2_reip_reg_23_, p2_reip_reg_24_, p2_reip_reg_25_, p2_reip_reg_26_,
p2_reip_reg_27_, p2_reip_reg_28_, p2_reip_reg_29_, p2_reip_reg_30_,
p2_reip_reg_31_, p2_byteenable_reg_3_, p2_byteenable_reg_2_,
p2_byteenable_reg_1_, p2_byteenable_reg_0_, p2_w_r_n_reg,
p2_flush_reg, p2_more_reg, p2_statebs16_reg, p2_requestpending_reg,
p2_d_c_n_reg, p2_m_io_n_reg, p2_codefetch_reg, p2_ads_n_reg,
p2_readrequest_reg, p2_memoryfetch_reg, p1_be_n_reg_3_,
p1_be_n_reg_2_, p1_be_n_reg_1_, p1_be_n_reg_0_, p1_state_reg_2_,
p1_state_reg_1_, p1_state_reg_0_, p1_datawidth_reg_0_,
p1_datawidth_reg_1_, p1_datawidth_reg_2_, p1_datawidth_reg_3_,
p1_datawidth_reg_4_, p1_datawidth_reg_5_, p1_datawidth_reg_6_,
p1_datawidth_reg_7_, p1_datawidth_reg_8_, p1_datawidth_reg_9_,
p1_datawidth_reg_10_, p1_datawidth_reg_11_, p1_datawidth_reg_12_,
p1_datawidth_reg_13_, p1_datawidth_reg_14_, p1_datawidth_reg_15_,
p1_datawidth_reg_16_, p1_datawidth_reg_17_, p1_datawidth_reg_18_,
p1_datawidth_reg_19_, p1_datawidth_reg_20_, p1_datawidth_reg_21_,
p1_datawidth_reg_22_, p1_datawidth_reg_23_, p1_datawidth_reg_24_,
p1_datawidth_reg_25_, p1_datawidth_reg_26_, p1_datawidth_reg_27_,
p1_datawidth_reg_28_, p1_datawidth_reg_29_, p1_datawidth_reg_30_,
p1_datawidth_reg_31_, p1_state2_reg_3_, p1_state2_reg_2_,
p1_state2_reg_1_, p1_state2_reg_0_, p1_instqueue_reg_15__7_,
p1_instqueue_reg_15__6_, p1_instqueue_reg_15__5_,
p1_instqueue_reg_15__4_, p1_instqueue_reg_15__3_,
p1_instqueue_reg_15__2_, p1_instqueue_reg_15__1_,
p1_instqueue_reg_15__0_, p1_instqueue_reg_14__7_,
p1_instqueue_reg_14__6_, p1_instqueue_reg_14__5_,
p1_instqueue_reg_14__4_, p1_instqueue_reg_14__3_,
p1_instqueue_reg_14__2_, p1_instqueue_reg_14__1_,
p1_instqueue_reg_14__0_, p1_instqueue_reg_13__7_,
p1_instqueue_reg_13__6_, p1_instqueue_reg_13__5_,
p1_instqueue_reg_13__4_, p1_instqueue_reg_13__3_,
p1_instqueue_reg_13__2_, p1_instqueue_reg_13__1_,
p1_instqueue_reg_13__0_, p1_instqueue_reg_12__7_,
p1_instqueue_reg_12__6_, p1_instqueue_reg_12__5_,
p1_instqueue_reg_12__4_, p1_instqueue_reg_12__3_,
p1_instqueue_reg_12__2_, p1_instqueue_reg_12__1_,
p1_instqueue_reg_12__0_, p1_instqueue_reg_11__7_,
p1_instqueue_reg_11__6_, p1_instqueue_reg_11__5_,
p1_instqueue_reg_11__4_, p1_instqueue_reg_11__3_,
p1_instqueue_reg_11__2_, p1_instqueue_reg_11__1_,
p1_instqueue_reg_11__0_, p1_instqueue_reg_10__7_,
p1_instqueue_reg_10__6_, p1_instqueue_reg_10__5_,
p1_instqueue_reg_10__4_, p1_instqueue_reg_10__3_,
p1_instqueue_reg_10__2_, p1_instqueue_reg_10__1_,
p1_instqueue_reg_10__0_, p1_instqueue_reg_9__7_,
p1_instqueue_reg_9__6_, p1_instqueue_reg_9__5_,
p1_instqueue_reg_9__4_, p1_instqueue_reg_9__3_,
p1_instqueue_reg_9__2_, p1_instqueue_reg_9__1_,
p1_instqueue_reg_9__0_, p1_instqueue_reg_8__7_,
p1_instqueue_reg_8__6_, p1_instqueue_reg_8__5_,
p1_instqueue_reg_8__4_, p1_instqueue_reg_8__3_,
p1_instqueue_reg_8__2_, p1_instqueue_reg_8__1_,
p1_instqueue_reg_8__0_, p1_instqueue_reg_7__7_,
p1_instqueue_reg_7__6_, p1_instqueue_reg_7__5_,
p1_instqueue_reg_7__4_, p1_instqueue_reg_7__3_,
p1_instqueue_reg_7__2_, p1_instqueue_reg_7__1_,
p1_instqueue_reg_7__0_, p1_instqueue_reg_6__7_,
p1_instqueue_reg_6__6_, p1_instqueue_reg_6__5_,
p1_instqueue_reg_6__4_, p1_instqueue_reg_6__3_,
p1_instqueue_reg_6__2_, p1_instqueue_reg_6__1_,
p1_instqueue_reg_6__0_, p1_instqueue_reg_5__7_,
p1_instqueue_reg_5__6_, p1_instqueue_reg_5__5_,
p1_instqueue_reg_5__4_, p1_instqueue_reg_5__3_,
p1_instqueue_reg_5__2_, p1_instqueue_reg_5__1_,
p1_instqueue_reg_5__0_, p1_instqueue_reg_4__7_,
p1_instqueue_reg_4__6_, p1_instqueue_reg_4__5_,
p1_instqueue_reg_4__4_, p1_instqueue_reg_4__3_,
p1_instqueue_reg_4__2_, p1_instqueue_reg_4__1_,
p1_instqueue_reg_4__0_, p1_instqueue_reg_3__7_,
p1_instqueue_reg_3__6_, p1_instqueue_reg_3__5_,
p1_instqueue_reg_3__4_, p1_instqueue_reg_3__3_,
p1_instqueue_reg_3__2_, p1_instqueue_reg_3__1_,
p1_instqueue_reg_3__0_, p1_instqueue_reg_2__7_,
p1_instqueue_reg_2__6_, p1_instqueue_reg_2__5_,
p1_instqueue_reg_2__4_, p1_instqueue_reg_2__3_,
p1_instqueue_reg_2__2_, p1_instqueue_reg_2__1_,
p1_instqueue_reg_2__0_, p1_instqueue_reg_1__7_,
p1_instqueue_reg_1__6_, p1_instqueue_reg_1__5_,
p1_instqueue_reg_1__4_, p1_instqueue_reg_1__3_,
p1_instqueue_reg_1__2_, p1_instqueue_reg_1__1_,
p1_instqueue_reg_1__0_, p1_instqueue_reg_0__7_,
p1_instqueue_reg_0__6_, p1_instqueue_reg_0__5_,
p1_instqueue_reg_0__4_, p1_instqueue_reg_0__3_,
p1_instqueue_reg_0__2_, p1_instqueue_reg_0__1_,
p1_instqueue_reg_0__0_, p1_instqueuerd_addr_reg_4_,
p1_instqueuerd_addr_reg_3_, p1_instqueuerd_addr_reg_2_,
p1_instqueuerd_addr_reg_1_, p1_instqueuerd_addr_reg_0_,
p1_instqueuewr_addr_reg_4_, p1_instqueuewr_addr_reg_3_,
p1_instqueuewr_addr_reg_2_, p1_instqueuewr_addr_reg_1_,
p1_instqueuewr_addr_reg_0_, p1_instaddrpointer_reg_0_,
p1_instaddrpointer_reg_1_, p1_instaddrpointer_reg_2_,
p1_instaddrpointer_reg_3_, p1_instaddrpointer_reg_4_,
p1_instaddrpointer_reg_5_, p1_instaddrpointer_reg_6_,
p1_instaddrpointer_reg_7_, p1_instaddrpointer_reg_8_,
p1_instaddrpointer_reg_9_, p1_instaddrpointer_reg_10_,
p1_instaddrpointer_reg_11_, p1_instaddrpointer_reg_12_,
p1_instaddrpointer_reg_13_, p1_instaddrpointer_reg_14_,
p1_instaddrpointer_reg_15_, p1_instaddrpointer_reg_16_,
p1_instaddrpointer_reg_17_, p1_instaddrpointer_reg_18_,
p1_instaddrpointer_reg_19_, p1_instaddrpointer_reg_20_,
p1_instaddrpointer_reg_21_, p1_instaddrpointer_reg_22_,
p1_instaddrpointer_reg_23_, p1_instaddrpointer_reg_24_,
p1_instaddrpointer_reg_25_, p1_instaddrpointer_reg_26_,
p1_instaddrpointer_reg_27_, p1_instaddrpointer_reg_28_,
p1_instaddrpointer_reg_29_, p1_instaddrpointer_reg_30_,
p1_instaddrpointer_reg_31_, p1_phyaddrpointer_reg_0_,
p1_phyaddrpointer_reg_1_, p1_phyaddrpointer_reg_2_,
p1_phyaddrpointer_reg_3_, p1_phyaddrpointer_reg_4_,
p1_phyaddrpointer_reg_5_, p1_phyaddrpointer_reg_6_,
p1_phyaddrpointer_reg_7_, p1_phyaddrpointer_reg_8_,
p1_phyaddrpointer_reg_9_, p1_phyaddrpointer_reg_10_,
p1_phyaddrpointer_reg_11_, p1_phyaddrpointer_reg_12_,
p1_phyaddrpointer_reg_13_, p1_phyaddrpointer_reg_14_,
p1_phyaddrpointer_reg_15_, p1_phyaddrpointer_reg_16_,
p1_phyaddrpointer_reg_17_, p1_phyaddrpointer_reg_18_,
p1_phyaddrpointer_reg_19_, p1_phyaddrpointer_reg_20_,
p1_phyaddrpointer_reg_21_, p1_phyaddrpointer_reg_22_,
p1_phyaddrpointer_reg_23_, p1_phyaddrpointer_reg_24_,
p1_phyaddrpointer_reg_25_, p1_phyaddrpointer_reg_26_,
p1_phyaddrpointer_reg_27_, p1_phyaddrpointer_reg_28_,
p1_phyaddrpointer_reg_29_, p1_phyaddrpointer_reg_30_,
p1_phyaddrpointer_reg_31_, p1_lword_reg_15_, p1_lword_reg_14_,
p1_lword_reg_13_, p1_lword_reg_12_, p1_lword_reg_11_,
p1_lword_reg_10_, p1_lword_reg_9_, p1_lword_reg_8_, p1_lword_reg_7_,
p1_lword_reg_6_, p1_lword_reg_5_, p1_lword_reg_4_, p1_lword_reg_3_,
p1_lword_reg_2_, p1_lword_reg_1_, p1_lword_reg_0_, p1_uword_reg_14_,
p1_uword_reg_13_, p1_uword_reg_12_, p1_uword_reg_11_,
p1_uword_reg_10_, p1_uword_reg_9_, p1_uword_reg_8_, p1_uword_reg_7_,
p1_uword_reg_6_, p1_uword_reg_5_, p1_uword_reg_4_, p1_uword_reg_3_,
p1_uword_reg_2_, p1_uword_reg_1_, p1_uword_reg_0_, p1_datao_reg_0_,
p1_datao_reg_1_, p1_datao_reg_2_, p1_datao_reg_3_, p1_datao_reg_4_,
p1_datao_reg_5_, p1_datao_reg_6_, p1_datao_reg_7_, p1_datao_reg_8_,
p1_datao_reg_9_, p1_datao_reg_10_, p1_datao_reg_11_, p1_datao_reg_12_,
p1_datao_reg_13_, p1_datao_reg_14_, p1_datao_reg_15_,
p1_datao_reg_16_, p1_datao_reg_17_, p1_datao_reg_18_,
p1_datao_reg_19_, p1_datao_reg_20_, p1_datao_reg_21_,
p1_datao_reg_22_, p1_datao_reg_23_, p1_datao_reg_24_,
p1_datao_reg_25_, p1_datao_reg_26_, p1_datao_reg_27_,
p1_datao_reg_28_, p1_datao_reg_29_, p1_datao_reg_30_,
p1_datao_reg_31_, p1_eax_reg_0_, p1_eax_reg_1_, p1_eax_reg_2_,
p1_eax_reg_3_, p1_eax_reg_4_, p1_eax_reg_5_, p1_eax_reg_6_,
p1_eax_reg_7_, p1_eax_reg_8_, p1_eax_reg_9_, p1_eax_reg_10_,
p1_eax_reg_11_, p1_eax_reg_12_, p1_eax_reg_13_, p1_eax_reg_14_,
p1_eax_reg_15_, p1_eax_reg_16_, p1_eax_reg_17_, p1_eax_reg_18_,
p1_eax_reg_19_, p1_eax_reg_20_, p1_eax_reg_21_, p1_eax_reg_22_,
p1_eax_reg_23_, p1_eax_reg_24_, p1_eax_reg_25_, p1_eax_reg_26_,
p1_eax_reg_27_, p1_eax_reg_28_, p1_eax_reg_29_, p1_eax_reg_30_,
p1_eax_reg_31_, p1_ebx_reg_0_, p1_ebx_reg_1_, p1_ebx_reg_2_,
p1_ebx_reg_3_, p1_ebx_reg_4_, p1_ebx_reg_5_, p1_ebx_reg_6_,
p1_ebx_reg_7_, p1_ebx_reg_8_, p1_ebx_reg_9_, p1_ebx_reg_10_,
p1_ebx_reg_11_, p1_ebx_reg_12_, p1_ebx_reg_13_, p1_ebx_reg_14_,
p1_ebx_reg_15_, p1_ebx_reg_16_, p1_ebx_reg_17_, p1_ebx_reg_18_,
p1_ebx_reg_19_, p1_ebx_reg_20_, p1_ebx_reg_21_, p1_ebx_reg_22_,
p1_ebx_reg_23_, p1_ebx_reg_24_, p1_ebx_reg_25_, p1_ebx_reg_26_,
p1_ebx_reg_27_, p1_ebx_reg_28_, p1_ebx_reg_29_, p1_ebx_reg_30_,
p1_ebx_reg_31_, p1_reip_reg_0_, p1_reip_reg_1_, p1_reip_reg_2_,
p1_reip_reg_3_, p1_reip_reg_4_, p1_reip_reg_5_, p1_reip_reg_6_,
p1_reip_reg_7_, p1_reip_reg_8_, p1_reip_reg_9_, p1_reip_reg_10_,
p1_reip_reg_11_, p1_reip_reg_12_, p1_reip_reg_13_, p1_reip_reg_14_,
p1_reip_reg_15_, p1_reip_reg_16_, p1_reip_reg_17_, p1_reip_reg_18_,
p1_reip_reg_19_, p1_reip_reg_20_, p1_reip_reg_21_, p1_reip_reg_22_,
p1_reip_reg_23_, p1_reip_reg_24_, p1_reip_reg_25_, p1_reip_reg_26_,
p1_reip_reg_27_, p1_reip_reg_28_, p1_reip_reg_29_, p1_reip_reg_30_,
p1_reip_reg_31_, p1_byteenable_reg_3_, p1_byteenable_reg_2_,
p1_byteenable_reg_1_, p1_byteenable_reg_0_, p1_w_r_n_reg,
p1_flush_reg, p1_more_reg, p1_statebs16_reg, p1_requestpending_reg,
p1_d_c_n_reg, p1_m_io_n_reg, p1_codefetch_reg, p1_ads_n_reg,
p1_readrequest_reg, p1_memoryfetch_reg, p1_address_reg_29_,
p1_address_reg_28_, p1_address_reg_27_, p1_address_reg_26_,
p1_address_reg_25_, p1_address_reg_24_, p1_address_reg_23_,
p1_address_reg_22_, p1_address_reg_21_, p1_address_reg_20_,
p1_address_reg_19_, p1_address_reg_18_, p1_address_reg_17_,
p1_address_reg_16_, p1_address_reg_15_, p1_address_reg_14_,
p1_address_reg_13_, p1_address_reg_12_, p1_address_reg_11_,
p1_address_reg_10_, p1_address_reg_9_, p1_address_reg_8_,
p1_address_reg_7_, p1_address_reg_6_, p1_address_reg_5_,
p1_address_reg_4_, p1_address_reg_3_, p1_address_reg_2_,
p1_address_reg_1_, p1_address_reg_0_;
output u355, u356, u357, u358, u359, u360, u361, u362, u363, u364, u366,
u367, u368, u369, u370, u371, u372, u373, u374, u375, u347, u348,
u349, u350, u351, u352, u353, u354, u365, u376, u247, u246, u245,
u244, u243, u242, u241, u240, u239, u238, u237, u236, u235, u234,
u233, u232, u231, u230, u229, u228, u227, u226, u225, u224, u223,
u222, u221, u220, u219, u218, u217, u216, u251, u252, u253, u254,
u255, u256, u257, u258, u259, u260, u261, u262, u263, u264, u265,
u266, u267, u268, u269, u270, u271, u272, u273, u274, u275, u276,
u277, u278, u279, u280, u281, u282, u212, u215, u213, u214, p3_u3274,
p3_u3275, p3_u3276, p3_u3277, p3_u3061, p3_u3060, p3_u3059, p3_u3058,
p3_u3057, p3_u3056, p3_u3055, p3_u3054, p3_u3053, p3_u3052, p3_u3051,
p3_u3050, p3_u3049, p3_u3048, p3_u3047, p3_u3046, p3_u3045, p3_u3044,
p3_u3043, p3_u3042, p3_u3041, p3_u3040, p3_u3039, p3_u3038, p3_u3037,
p3_u3036, p3_u3035, p3_u3034, p3_u3033, p3_u3032, p3_u3031, p3_u3030,
p3_u3029, p3_u3280, p3_u3281, p3_u3028, p3_u3027, p3_u3026, p3_u3025,
p3_u3024, p3_u3023, p3_u3022, p3_u3021, p3_u3020, p3_u3019, p3_u3018,
p3_u3017, p3_u3016, p3_u3015, p3_u3014, p3_u3013, p3_u3012, p3_u3011,
p3_u3010, p3_u3009, p3_u3008, p3_u3007, p3_u3006, p3_u3005, p3_u3004,
p3_u3003, p3_u3002, p3_u3001, p3_u3000, p3_u2999, p3_u3282, p3_u2998,
p3_u2997, p3_u2996, p3_u2995, p3_u2994, p3_u2993, p3_u2992, p3_u2991,
p3_u2990, p3_u2989, p3_u2988, p3_u2987, p3_u2986, p3_u2985, p3_u2984,
p3_u2983, p3_u2982, p3_u2981, p3_u2980, p3_u2979, p3_u2978, p3_u2977,
p3_u2976, p3_u2975, p3_u2974, p3_u2973, p3_u2972, p3_u2971, p3_u2970,
p3_u2969, p3_u2968, p3_u2967, p3_u2966, p3_u2965, p3_u2964, p3_u2963,
p3_u2962, p3_u2961, p3_u2960, p3_u2959, p3_u2958, p3_u2957, p3_u2956,
p3_u2955, p3_u2954, p3_u2953, p3_u2952, p3_u2951, p3_u2950, p3_u2949,
p3_u2948, p3_u2947, p3_u2946, p3_u2945, p3_u2944, p3_u2943, p3_u2942,
p3_u2941, p3_u2940, p3_u2939, p3_u2938, p3_u2937, p3_u2936, p3_u2935,
p3_u2934, p3_u2933, p3_u2932, p3_u2931, p3_u2930, p3_u2929, p3_u2928,
p3_u2927, p3_u2926, p3_u2925, p3_u2924, p3_u2923, p3_u2922, p3_u2921,
p3_u2920, p3_u2919, p3_u2918, p3_u2917, p3_u2916, p3_u2915, p3_u2914,
p3_u2913, p3_u2912, p3_u2911, p3_u2910, p3_u2909, p3_u2908, p3_u2907,
p3_u2906, p3_u2905, p3_u2904, p3_u2903, p3_u2902, p3_u2901, p3_u2900,
p3_u2899, p3_u2898, p3_u2897, p3_u2896, p3_u2895, p3_u2894, p3_u2893,
p3_u2892, p3_u2891, p3_u2890, p3_u2889, p3_u2888, p3_u2887, p3_u2886,
p3_u2885, p3_u2884, p3_u2883, p3_u2882, p3_u2881, p3_u2880, p3_u2879,
p3_u2878, p3_u2877, p3_u2876, p3_u2875, p3_u2874, p3_u2873, p3_u2872,
p3_u2871, p3_u2870, p3_u2869, p3_u2868, p3_u3284, p3_u3285, p3_u3288,
p3_u3289, p3_u3290, p3_u2867, p3_u2866, p3_u2865, p3_u2864, p3_u2863,
p3_u2862, p3_u2861, p3_u2860, p3_u2859, p3_u2858, p3_u2857, p3_u2856,
p3_u2855, p3_u2854, p3_u2853, p3_u2852, p3_u2851, p3_u2850, p3_u2849,
p3_u2848, p3_u2847, p3_u2846, p3_u2845, p3_u2844, p3_u2843, p3_u2842,
p3_u2841, p3_u2840, p3_u2839, p3_u2838, p3_u2837, p3_u2836, p3_u2835,
p3_u2834, p3_u2833, p3_u2832, p3_u2831, p3_u2830, p3_u2829, p3_u2828,
p3_u2827, p3_u2826, p3_u2825, p3_u2824, p3_u2823, p3_u2822, p3_u2821,
p3_u2820, p3_u2819, p3_u2818, p3_u2817, p3_u2816, p3_u2815, p3_u2814,
p3_u2813, p3_u2812, p3_u2811, p3_u2810, p3_u2809, p3_u2808, p3_u2807,
p3_u2806, p3_u2805, p3_u2804, p3_u2803, p3_u2802, p3_u2801, p3_u2800,
p3_u2799, p3_u2798, p3_u2797, p3_u2796, p3_u2795, p3_u2794, p3_u2793,
p3_u2792, p3_u2791, p3_u2790, p3_u2789, p3_u2788, p3_u2787, p3_u2786,
p3_u2785, p3_u2784, p3_u2783, p3_u2782, p3_u2781, p3_u2780, p3_u2779,
p3_u2778, p3_u2777, p3_u2776, p3_u2775, p3_u2774, p3_u2773, p3_u2772,
p3_u2771, p3_u2770, p3_u2769, p3_u2768, p3_u2767, p3_u2766, p3_u2765,
p3_u2764, p3_u2763, p3_u2762, p3_u2761, p3_u2760, p3_u2759, p3_u2758,
p3_u2757, p3_u2756, p3_u2755, p3_u2754, p3_u2753, p3_u2752, p3_u2751,
p3_u2750, p3_u2749, p3_u2748, p3_u2747, p3_u2746, p3_u2745, p3_u2744,
p3_u2743, p3_u2742, p3_u2741, p3_u2740, p3_u2739, p3_u2738, p3_u2737,
p3_u2736, p3_u2735, p3_u2734, p3_u2733, p3_u2732, p3_u2731, p3_u2730,
p3_u2729, p3_u2728, p3_u2727, p3_u2726, p3_u2725, p3_u2724, p3_u2723,
p3_u2722, p3_u2721, p3_u2720, p3_u2719, p3_u2718, p3_u2717, p3_u2716,
p3_u2715, p3_u2714, p3_u2713, p3_u2712, p3_u2711, p3_u2710, p3_u2709,
p3_u2708, p3_u2707, p3_u2706, p3_u2705, p3_u2704, p3_u2703, p3_u2702,
p3_u2701, p3_u2700, p3_u2699, p3_u2698, p3_u2697, p3_u2696, p3_u2695,
p3_u2694, p3_u2693, p3_u2692, p3_u2691, p3_u2690, p3_u2689, p3_u2688,
p3_u2687, p3_u2686, p3_u2685, p3_u2684, p3_u2683, p3_u2682, p3_u2681,
p3_u2680, p3_u2679, p3_u2678, p3_u2677, p3_u2676, p3_u2675, p3_u2674,
p3_u2673, p3_u2672, p3_u2671, p3_u2670, p3_u2669, p3_u2668, p3_u2667,
p3_u2666, p3_u2665, p3_u2664, p3_u2663, p3_u2662, p3_u2661, p3_u2660,
p3_u2659, p3_u2658, p3_u2657, p3_u2656, p3_u2655, p3_u2654, p3_u2653,
p3_u2652, p3_u2651, p3_u2650, p3_u2649, p3_u2648, p3_u2647, p3_u2646,
p3_u2645, p3_u2644, p3_u2643, p3_u2642, p3_u2641, p3_u2640, p3_u2639,
p3_u3292, p3_u2638, p3_u3293, p3_u3294, p3_u2637, p3_u3295, p3_u2636,
p3_u3296, p3_u2635, p3_u3297, p3_u2634, p3_u2633, p3_u3298, p3_u3299,
p2_u3585, p2_u3586, p2_u3587, p2_u3588, p2_u3241, p2_u3240, p2_u3239,
p2_u3238, p2_u3237, p2_u3236, p2_u3235, p2_u3234, p2_u3233, p2_u3232,
p2_u3231, p2_u3230, p2_u3229, p2_u3228, p2_u3227, p2_u3226, p2_u3225,
p2_u3224, p2_u3223, p2_u3222, p2_u3221, p2_u3220, p2_u3219, p2_u3218,
p2_u3217, p2_u3216, p2_u3215, p2_u3214, p2_u3213, p2_u3212, p2_u3211,
p2_u3210, p2_u3209, p2_u3591, p2_u3592, p2_u3208, p2_u3207, p2_u3206,
p2_u3205, p2_u3204, p2_u3203, p2_u3202, p2_u3201, p2_u3200, p2_u3199,
p2_u3198, p2_u3197, p2_u3196, p2_u3195, p2_u3194, p2_u3193, p2_u3192,
p2_u3191, p2_u3190, p2_u3189, p2_u3188, p2_u3187, p2_u3186, p2_u3185,
p2_u3184, p2_u3183, p2_u3182, p2_u3181, p2_u3180, p2_u3179, p2_u3593,
p2_u3178, p2_u3177, p2_u3176, p2_u3175, p2_u3174, p2_u3173, p2_u3172,
p2_u3171, p2_u3170, p2_u3169, p2_u3168, p2_u3167, p2_u3166, p2_u3165,
p2_u3164, p2_u3163, p2_u3162, p2_u3161, p2_u3160, p2_u3159, p2_u3158,
p2_u3157, p2_u3156, p2_u3155, p2_u3154, p2_u3153, p2_u3152, p2_u3151,
p2_u3150, p2_u3149, p2_u3148, p2_u3147, p2_u3146, p2_u3145, p2_u3144,
p2_u3143, p2_u3142, p2_u3141, p2_u3140, p2_u3139, p2_u3138, p2_u3137,
p2_u3136, p2_u3135, p2_u3134, p2_u3133, p2_u3132, p2_u3131, p2_u3130,
p2_u3129, p2_u3128, p2_u3127, p2_u3126, p2_u3125, p2_u3124, p2_u3123,
p2_u3122, p2_u3121, p2_u3120, p2_u3119, p2_u3118, p2_u3117, p2_u3116,
p2_u3115, p2_u3114, p2_u3113, p2_u3112, p2_u3111, p2_u3110, p2_u3109,
p2_u3108, p2_u3107, p2_u3106, p2_u3105, p2_u3104, p2_u3103, p2_u3102,
p2_u3101, p2_u3100, p2_u3099, p2_u3098, p2_u3097, p2_u3096, p2_u3095,
p2_u3094, p2_u3093, p2_u3092, p2_u3091, p2_u3090, p2_u3089, p2_u3088,
p2_u3087, p2_u3086, p2_u3085, p2_u3084, p2_u3083, p2_u3082, p2_u3081,
p2_u3080, p2_u3079, p2_u3078, p2_u3077, p2_u3076, p2_u3075, p2_u3074,
p2_u3073, p2_u3072, p2_u3071, p2_u3070, p2_u3069, p2_u3068, p2_u3067,
p2_u3066, p2_u3065, p2_u3064, p2_u3063, p2_u3062, p2_u3061, p2_u3060,
p2_u3059, p2_u3058, p2_u3057, p2_u3056, p2_u3055, p2_u3054, p2_u3053,
p2_u3052, p2_u3051, p2_u3050, p2_u3049, p2_u3048, p2_u3595, p2_u3596,
p2_u3599, p2_u3600, p2_u3601, p2_u3047, p2_u3602, p2_u3603, p2_u3604,
p2_u3605, p2_u3046, p2_u3045, p2_u3044, p2_u3043, p2_u3042, p2_u3041,
p2_u3040, p2_u3039, p2_u3038, p2_u3037, p2_u3036, p2_u3035, p2_u3034,
p2_u3033, p2_u3032, p2_u3031, p2_u3030, p2_u3029, p2_u3028, p2_u3027,
p2_u3026, p2_u3025, p2_u3024, p2_u3023, p2_u3022, p2_u3021, p2_u3020,
p2_u3019, p2_u3018, p2_u3017, p2_u3016, p2_u3015, p2_u3014, p2_u3013,
p2_u3012, p2_u3011, p2_u3010, p2_u3009, p2_u3008, p2_u3007, p2_u3006,
p2_u3005, p2_u3004, p2_u3003, p2_u3002, p2_u3001, p2_u3000, p2_u2999,
p2_u2998, p2_u2997, p2_u2996, p2_u2995, p2_u2994, p2_u2993, p2_u2992,
p2_u2991, p2_u2990, p2_u2989, p2_u2988, p2_u2987, p2_u2986, p2_u2985,
p2_u2984, p2_u2983, p2_u2982, p2_u2981, p2_u2980, p2_u2979, p2_u2978,
p2_u2977, p2_u2976, p2_u2975, p2_u2974, p2_u2973, p2_u2972, p2_u2971,
p2_u2970, p2_u2969, p2_u2968, p2_u2967, p2_u2966, p2_u2965, p2_u2964,
p2_u2963, p2_u2962, p2_u2961, p2_u2960, p2_u2959, p2_u2958, p2_u2957,
p2_u2956, p2_u2955, p2_u2954, p2_u2953, p2_u2952, p2_u2951, p2_u2950,
p2_u2949, p2_u2948, p2_u2947, p2_u2946, p2_u2945, p2_u2944, p2_u2943,
p2_u2942, p2_u2941, p2_u2940, p2_u2939, p2_u2938, p2_u2937, p2_u2936,
p2_u2935, p2_u2934, p2_u2933, p2_u2932, p2_u2931, p2_u2930, p2_u2929,
p2_u2928, p2_u2927, p2_u2926, p2_u2925, p2_u2924, p2_u2923, p2_u2922,
p2_u2921, p2_u2920, p2_u2919, p2_u2918, p2_u2917, p2_u2916, p2_u2915,
p2_u2914, p2_u2913, p2_u2912, p2_u2911, p2_u2910, p2_u2909, p2_u2908,
p2_u2907, p2_u2906, p2_u2905, p2_u2904, p2_u2903, p2_u2902, p2_u2901,
p2_u2900, p2_u2899, p2_u2898, p2_u2897, p2_u2896, p2_u2895, p2_u2894,
p2_u2893, p2_u2892, p2_u2891, p2_u2890, p2_u2889, p2_u2888, p2_u2887,
p2_u2886, p2_u2885, p2_u2884, p2_u2883, p2_u2882, p2_u2881, p2_u2880,
p2_u2879, p2_u2878, p2_u2877, p2_u2876, p2_u2875, p2_u2874, p2_u2873,
p2_u2872, p2_u2871, p2_u2870, p2_u2869, p2_u2868, p2_u2867, p2_u2866,
p2_u2865, p2_u2864, p2_u2863, p2_u2862, p2_u2861, p2_u2860, p2_u2859,
p2_u2858, p2_u2857, p2_u2856, p2_u2855, p2_u2854, p2_u2853, p2_u2852,
p2_u2851, p2_u2850, p2_u2849, p2_u2848, p2_u2847, p2_u2846, p2_u2845,
p2_u2844, p2_u2843, p2_u2842, p2_u2841, p2_u2840, p2_u2839, p2_u2838,
p2_u2837, p2_u2836, p2_u2835, p2_u2834, p2_u2833, p2_u2832, p2_u2831,
p2_u2830, p2_u2829, p2_u2828, p2_u2827, p2_u2826, p2_u2825, p2_u2824,
p2_u2823, p2_u2822, p2_u2821, p2_u2820, p2_u3608, p2_u2819, p2_u3609,
p2_u2818, p2_u3610, p2_u2817, p2_u3611, p2_u2816, p2_u2815, p2_u3612,
p2_u2814, p1_u3458, p1_u3459, p1_u3460, p1_u3461, p1_u3226, p1_u3225,
p1_u3224, p1_u3223, p1_u3222, p1_u3221, p1_u3220, p1_u3219, p1_u3218,
p1_u3217, p1_u3216, p1_u3215, p1_u3214, p1_u3213, p1_u3212, p1_u3211,
p1_u3210, p1_u3209, p1_u3208, p1_u3207, p1_u3206, p1_u3205, p1_u3204,
p1_u3203, p1_u3202, p1_u3201, p1_u3200, p1_u3199, p1_u3198, p1_u3197,
p1_u3196, p1_u3195, p1_u3194, p1_u3464, p1_u3465, p1_u3193, p1_u3192,
p1_u3191, p1_u3190, p1_u3189, p1_u3188, p1_u3187, p1_u3186, p1_u3185,
p1_u3184, p1_u3183, p1_u3182, p1_u3181, p1_u3180, p1_u3179, p1_u3178,
p1_u3177, p1_u3176, p1_u3175, p1_u3174, p1_u3173, p1_u3172, p1_u3171,
p1_u3170, p1_u3169, p1_u3168, p1_u3167, p1_u3166, p1_u3165, p1_u3164,
p1_u3466, p1_u3163, p1_u3162, p1_u3161, p1_u3160, p1_u3159, p1_u3158,
p1_u3157, p1_u3156, p1_u3155, p1_u3154, p1_u3153, p1_u3152, p1_u3151,
p1_u3150, p1_u3149, p1_u3148, p1_u3147, p1_u3146, p1_u3145, p1_u3144,
p1_u3143, p1_u3142, p1_u3141, p1_u3140, p1_u3139, p1_u3138, p1_u3137,
p1_u3136, p1_u3135, p1_u3134, p1_u3133, p1_u3132, p1_u3131, p1_u3130,
p1_u3129, p1_u3128, p1_u3127, p1_u3126, p1_u3125, p1_u3124, p1_u3123,
p1_u3122, p1_u3121, p1_u3120, p1_u3119, p1_u3118, p1_u3117, p1_u3116,
p1_u3115, p1_u3114, p1_u3113, p1_u3112, p1_u3111, p1_u3110, p1_u3109,
p1_u3108, p1_u3107, p1_u3106, p1_u3105, p1_u3104, p1_u3103, p1_u3102,
p1_u3101, p1_u3100, p1_u3099, p1_u3098, p1_u3097, p1_u3096, p1_u3095,
p1_u3094, p1_u3093, p1_u3092, p1_u3091, p1_u3090, p1_u3089, p1_u3088,
p1_u3087, p1_u3086, p1_u3085, p1_u3084, p1_u3083, p1_u3082, p1_u3081,
p1_u3080, p1_u3079, p1_u3078, p1_u3077, p1_u3076, p1_u3075, p1_u3074,
p1_u3073, p1_u3072, p1_u3071, p1_u3070, p1_u3069, p1_u3068, p1_u3067,
p1_u3066, p1_u3065, p1_u3064, p1_u3063, p1_u3062, p1_u3061, p1_u3060,
p1_u3059, p1_u3058, p1_u3057, p1_u3056, p1_u3055, p1_u3054, p1_u3053,
p1_u3052, p1_u3051, p1_u3050, p1_u3049, p1_u3048, p1_u3047, p1_u3046,
p1_u3045, p1_u3044, p1_u3043, p1_u3042, p1_u3041, p1_u3040, p1_u3039,
p1_u3038, p1_u3037, p1_u3036, p1_u3035, p1_u3034, p1_u3033, p1_u3468,
p1_u3469, p1_u3472, p1_u3473, p1_u3474, p1_u3032, p1_u3475, p1_u3476,
p1_u3477, p1_u3478, p1_u3031, p1_u3030, p1_u3029, p1_u3028, p1_u3027,
p1_u3026, p1_u3025, p1_u3024, p1_u3023, p1_u3022, p1_u3021, p1_u3020,
p1_u3019, p1_u3018, p1_u3017, p1_u3016, p1_u3015, p1_u3014, p1_u3013,
p1_u3012, p1_u3011, p1_u3010, p1_u3009, p1_u3008, p1_u3007, p1_u3006,
p1_u3005, p1_u3004, p1_u3003, p1_u3002, p1_u3001, p1_u3000, p1_u2999,
p1_u2998, p1_u2997, p1_u2996, p1_u2995, p1_u2994, p1_u2993, p1_u2992,
p1_u2991, p1_u2990, p1_u2989, p1_u2988, p1_u2987, p1_u2986, p1_u2985,
p1_u2984, p1_u2983, p1_u2982, p1_u2981, p1_u2980, p1_u2979, p1_u2978,
p1_u2977, p1_u2976, p1_u2975, p1_u2974, p1_u2973, p1_u2972, p1_u2971,
p1_u2970, p1_u2969, p1_u2968, p1_u2967, p1_u2966, p1_u2965, p1_u2964,
p1_u2963, p1_u2962, p1_u2961, p1_u2960, p1_u2959, p1_u2958, p1_u2957,
p1_u2956, p1_u2955, p1_u2954, p1_u2953, p1_u2952, p1_u2951, p1_u2950,
p1_u2949, p1_u2948, p1_u2947, p1_u2946, p1_u2945, p1_u2944, p1_u2943,
p1_u2942, p1_u2941, p1_u2940, p1_u2939, p1_u2938, p1_u2937, p1_u2936,
p1_u2935, p1_u2934, p1_u2933, p1_u2932, p1_u2931, p1_u2930, p1_u2929,
p1_u2928, p1_u2927, p1_u2926, p1_u2925, p1_u2924, p1_u2923, p1_u2922,
p1_u2921, p1_u2920, p1_u2919, p1_u2918, p1_u2917, p1_u2916, p1_u2915,
p1_u2914, p1_u2913, p1_u2912, p1_u2911, p1_u2910, p1_u2909, p1_u2908,
p1_u2907, p1_u2906, p1_u2905, p1_u2904, p1_u2903, p1_u2902, p1_u2901,
p1_u2900, p1_u2899, p1_u2898, p1_u2897, p1_u2896, p1_u2895, p1_u2894,
p1_u2893, p1_u2892, p1_u2891, p1_u2890, p1_u2889, p1_u2888, p1_u2887,
p1_u2886, p1_u2885, p1_u2884, p1_u2883, p1_u2882, p1_u2881, p1_u2880,
p1_u2879, p1_u2878, p1_u2877, p1_u2876, p1_u2875, p1_u2874, p1_u2873,
p1_u2872, p1_u2871, p1_u2870, p1_u2869, p1_u2868, p1_u2867, p1_u2866,
p1_u2865, p1_u2864, p1_u2863, p1_u2862, p1_u2861, p1_u2860, p1_u2859,
p1_u2858, p1_u2857, p1_u2856, p1_u2855, p1_u2854, p1_u2853, p1_u2852,
p1_u2851, p1_u2850, p1_u2849, p1_u2848, p1_u2847, p1_u2846, p1_u2845,
p1_u2844, p1_u2843, p1_u2842, p1_u2841, p1_u2840, p1_u2839, p1_u2838,
p1_u2837, p1_u2836, p1_u2835, p1_u2834, p1_u2833, p1_u2832, p1_u2831,
p1_u2830, p1_u2829, p1_u2828, p1_u2827, p1_u2826, p1_u2825, p1_u2824,
p1_u2823, p1_u2822, p1_u2821, p1_u2820, p1_u2819, p1_u2818, p1_u2817,
p1_u2816, p1_u2815, p1_u2814, p1_u2813, p1_u2812, p1_u2811, p1_u2810,
p1_u2809, p1_u2808, p1_u3481, p1_u2807, p1_u3482, p1_u3483, p1_u2806,
p1_u3484, p1_u2805, p1_u3485, p1_u2804, p1_u3486, p1_u2803, p1_u2802,
p1_u3487, p1_u2801;
wire   n53114, n53115, n53116, n53117, n53118, n53119, n53120, n53121,
n53122, n53123, n53124, n53125, n53126, n53127, n53128, n53129,
n53130, n53131, n53132, n53133, n53134, n53135, n53136, n53137,
n53138, n53139, n53140, n53141, n53142, n53143, n53144, n53145,
n53146, n53147, n53148, n53149, n53150, n53151, n53152, n53153,
n53154, n53155, n53156, n53157, n53158, n53159, n53160, n53161,
n53162, n53163, n53164, n53165, n53166, n53167, n53168, n53169,
n53170, n25181, n25182, n25183, n25184, n25186, n25188, n25190,
n25192, n25194, n25196, n25198, n25200, n25202, n25204, n25206,
n25208, n25210, n25212, n25214, n25216, n25218, n25220, n25222,
n25224, n25226, n25228, n25230, n25232, n25234, n25236, n25238,
n25240, n25242, n25244, n25246, n25248, n25250, n25252, n25254,
n25256, n25258, n25260, n25262, n25264, n25266, n25268, n25270,
n25272, n25274, n25276, n25278, n25280, n25282, n25284, n25286,
n25288, n25290, n25292, n25294, n25296, n25298, n25300, n25302,
n25304, n25306, n25308, n25310, n25312, n25314, n25316, n25318,
n25320, n25322, n25324, n25326, n25328, n25330, n25332, n25334,
n25336, n25338, n25340, n25342, n25344, n25346, n25348, n25350,
n25352, n25354, n25356, n25358, n25360, n25362, n25364, n25366,
n25368, n25370, n25372, n25374, n25376, n25378, n25380, n25382,
n25384, n25386, n25388, n25390, n25392, n25394, n25396, n25398,
n25400, n25402, n25404, n25406, n25408, n25410, n25412, n25414,
n25416, n25418, n25420, n25422, n25424, n25426, n25428, n25430,
n25432, n25434, n25436, n25438, n25440, n25442, n25444, n25446,
n25448, n25450, n25452, n25454, n25456, n25458, n25460, n25462,
n25464, n25466, n25468, n25470, n25472, n25474, n25476, n25478,
n25480, n25482, n25484, n25486, n25488, n25490, n25492, n25494,
n25496, n25498, n25500, n25502, n25504, n25506, n25508, n25510,
n25512, n25514, n25516, n25518, n25520, n25522, n25524, n25526,
n25528, n25530, n25532, n25534, n25536, n25538, n25540, n25542,
n25544, n25546, n25548, n25550, n25552, n25554, n25556, n25558,
n25560, n25562, n25564, n25566, n25568, n25570, n25572, n25574,
n25576, n25578, n25580, n25582, n25584, n25586, n25588, n25590,
n25592, n25594, n25596, n25598, n25600, n25602, n25604, n25606,
n25608, n25610, n25612, n25614, n25616, n25618, n25620, n25622,
n25624, n25626, n25628, n25630, n25632, n25634, n25636, n25638,
n25640, n25642, n25644, n25646, n25648, n25650, n25652, n25654,
n25656, n25658, n25660, n25662, n25664, n25666, n25668, n25670,
n25672, n25674, n25676, n25678, n25680, n25682, n25684, n25686,
n25688, n25690, n25692, n25694, n25696, n25698, n25700, n25702,
n25704, n25706, n25708, n25710, n25712, n25714, n25716, n25718,
n25720, n25722, n25724, n25726, n25728, n25730, n25732, n25734,
n25736, n25738, n25740, n25742, n25744, n25746, n25748, n25750,
n25752, n25754, n25756, n25758, n25760, n25762, n25764, n25766,
n25768, n25770, n25772, n25774, n25776, n25778, n25780, n25782,
n25784, n25786, n25788, n25790, n25792, n25794, n25796, n25798,
n25800, n25802, n25804, n25806, n25808, n25810, n25812, n25814,
n25816, n25818, n25820, n25822, n25824, n25826, n25828, n25830,
n25832, n25834, n25836, n25838, n25840, n25842, n25844, n25846,
n25848, n25850, n25852, n25854, n25856, n25858, n25860, n25862,
n25864, n25866, n25868, n25870, n25872, n25874, n25876, n25878,
n25880, n25882, n25884, n25886, n25888, n25890, n25892, n25894,
n25896, n25898, n25900, n25902, n25904, n25906, n25908, n25910,
n25912, n25914, n25916, n25918, n25920, n25922, n25924, n25926,
n25928, n25930, n25932, n25934, n25936, n25938, n25940, n25942,
n25944, n25946, n25948, n25950, n25952, n25954, n25956, n25958,
n25960, n25962, n25964, n25966, n25968, n25970, n25972, n25974,
n25976, n25978, n25980, n25982, n25984, n25986, n25988, n25990,
n25992, n25994, n25996, n25998, n26000, n26002, n26004, n26006,
n26008, n26010, n26012, n26014, n26016, n26018, n26020, n26022,
n26024, n26026, n26028, n26030, n26032, n26034, n26036, n26038,
n26040, n26042, n26044, n26046, n26048, n26050, n26052, n26054,
n26056, n26058, n26060, n26062, n26064, n26066, n26068, n26070,
n26072, n26074, n26076, n26078, n26080, n26082, n26084, n26086,
n26088, n26090, n26092, n26094, n26096, n26098, n26100, n26102,
n26104, n26106, n26108, n26110, n26112, n26114, n26116, n26118,
n26120, n26122, n26124, n26126, n26128, n26130, n26132, n26134,
n26136, n26138, n26140, n26142, n26144, n26146, n26148, n26150,
n26152, n26154, n26156, n26158, n26160, n26162, n26164, n26166,
n26168, n26170, n26172, n26174, n26176, n26178, n26180, n26182,
n26184, n26186, n26188, n26190, n26192, n26194, n26196, n26198,
n26200, n26202, n26204, n26206, n26208, n26210, n26212, n26214,
n26216, n26218, n26220, n26222, n26224, n26226, n26228, n26230,
n26232, n26234, n26236, n26238, n26240, n26242, n26244, n26246,
n26248, n26250, n26252, n26254, n26256, n26258, n26260, n26262,
n26264, n26266, n26268, n26270, n26272, n26274, n26276, n26278,
n26280, n26282, n26284, n26286, n26288, n26290, n26292, n26294,
n26296, n26298, n26300, n26302, n26304, n26306, n26308, n26310,
n26312, n26314, n26316, n26318, n26320, n26322, n26324, n26326,
n26328, n26330, n26332, n26334, n26336, n26338, n26340, n26342,
n26344, n26346, n26348, n26350, n26352, n26354, n26356, n26358,
n26360, n26362, n26364, n26366, n26368, n26370, n26372, n26374,
n26376, n26378, n26380, n26382, n26384, n26386, n26388, n26390,
n26392, n26394, n26396, n26398, n26400, n26402, n26404, n26406,
n26408, n26410, n26412, n26414, n26416, n26418, n26420, n26422,
n26424, n26426, n26428, n26430, n26432, n26434, n26436, n26438,
n26440, n26442, n26444, n26446, n26448, n26450, n26452, n26454,
n26456, n26458, n26460, n26462, n26464, n26466, n26468, n26470,
n26472, n26474, n26476, n26478, n26480, n26482, n26484, n26486,
n26488, n26490, n26492, n26494, n26496, n26498, n26500, n26502,
n26504, n26506, n26508, n26510, n26512, n26514, n26516, n26518,
n26520, n26522, n26524, n26526, n26528, n26530, n26532, n26534,
n26536, n26538, n26540, n26542, n26544, n26546, n26548, n26550,
n26552, n26554, n26556, n26558, n26560, n26562, n26564, n26566,
n26568, n26570, n26572, n26574, n26576, n26578, n26580, n26582,
n26584, n26586, n26588, n26590, n26592, n26594, n26596, n26598,
n26600, n26602, n26604, n26606, n26608, n26610, n26612, n26614,
n26616, n26618, n26620, n26622, n26624, n26626, n26628, n26630,
n26632, n26634, n26636, n26638, n26640, n26642, n26644, n26646,
n26648, n26650, n26652, n26654, n26656, n26658, n26660, n26662,
n26664, n26666, n26668, n26670, n26672, n26674, n26676, n26678,
n26680, n26682, n26684, n26686, n26688, n26690, n26692, n26694,
n26696, n26698, n26700, n26702, n26704, n26706, n26708, n26710,
n26712, n26714, n26716, n26718, n26720, n26722, n26724, n26726,
n26728, n26730, n26732, n26734, n26736, n26738, n26740, n26742,
n26744, n26746, n26748, n26750, n26752, n26754, n26756, n26758,
n26760, n26762, n26764, n26766, n26768, n26770, n26772, n26774,
n26776, n26778, n26780, n26782, n26784, n26786, n26788, n26790,
n26792, n26794, n26796, n26798, n26800, n26802, n26804, n26806,
n26808, n26810, n26812, n26814, n26816, n26818, n26820, n26822,
n26824, n26826, n26828, n26830, n26832, n26834, n26836, n26838,
n26840, n26842, n26844, n26846, n26848, n26850, n26852, n26854,
n26856, n26858, n26860, n26862, n26864, n26866, n26868, n26870,
n26872, n26874, n26876, n26878, n26880, n26882, n26884, n26886,
n26888, n26890, n26892, n26894, n26896, n26898, n26900, n26902,
n26904, n26906, n26908, n26910, n26912, n26914, n26916, n26918,
n26920, n26922, n26924, n26926, n26928, n26930, n26932, n26934,
n26936, n26938, n26940, n26942, n26944, n26946, n26948, n26950,
n26952, n26954, n26956, n26958, n26960, n26962, n26964, n26966,
n26968, n26970, n26972, n26974, n26976, n26978, n26980, n26982,
n26984, n26986, n26988, n26990, n26992, n26994, n26996, n26998,
n27000, n27002, n27004, n27006, n27008, n27010, n27012, n27014,
n27016, n27018, n27020, n27022, n27024, n27026, n27028, n27030,
n27032, n27034, n27036, n27038, n27040, n27042, n27044, n27046,
n27048, n27050, n27052, n27054, n27056, n27058, n27060, n27062,
n27064, n27066, n27068, n27070, n27072, n27074, n27076, n27078,
n27080, n27082, n27084, n27086, n27088, n27090, n27092, n27094,
n27096, n27098, n27100, n27102, n27104, n27106, n27108, n27110,
n27112, n27114, n27116, n27118, n27120, n27122, n27124, n27126,
n27128, n27130, n27132, n27134, n27136, n27138, n27140, n27142,
n27144, n27146, n27148, n27150, n27152, n27154, n27156, n27158,
n27160, n27162, n27164, n27166, n27168, n27170, n27172, n27174,
n27176, n27178, n27180, n27182, n27184, n27186, n27188, n27190,
n27192, n27194, n27196, n27198, n27200, n27202, n27204, n27206,
n27208, n27210, n27212, n27214, n27216, n27218, n27220, n27222,
n27224, n27226, n27228, n27230, n27232, n27234, n27236, n27238,
n27240, n27242, n27244, n27246, n27248, n27250, n27252, n27254,
n27256, n27258, n27260, n27262, n27264, n27266, n27268, n27270,
n27272, n27274, n27276, n27278, n27280, n27282, n27284, n27286,
n27288, n27290, n27292, n27294, n27296, n27298, n27300, n27302,
n27304, n27306, n27308, n27310, n27312, n27314, n27316, n27318,
n27320, n27322, n27324, n27326, n27328, n27330, n27332, n27334,
n27336, n27338, n27340, n27342, n27344, n27346, n27348, n27350,
n27352, n27354, n27356, n27358, n27360, n27362, n27364, n27366,
n27368, n27370, n27372, n27374, n27376, n27378, n27380, n27382,
n27384, n27386, n27388, n27390, n27392, n27394, n27396, n27398,
n27400, n27402, n27404, n27406, n27408, n27410, n27412, n27414,
n27416, n27418, n27420, n27422, n27424, n27426, n27428, n27430,
n27432, n27434, n27436, n27438, n27440, n27442, n27444, n27446,
n27448, n27450, n27452, n27454, n27456, n27458, n27460, n27462,
n27464, n27466, n27468, n27470, n27472, n27474, n27476, n27478,
n27480, n27482, n27484, n27486, n27488, n27490, n27492, n27494,
n27496, n27498, n27500, n27502, n27504, n27506, n27508, n27510,
n27512, n27514, n27516, n27518, n27520, n27522, n27524, n27526,
n27528, n27530, n27532, n27534, n27536, n27538, n27540, n27542,
n27544, n27546, n27548, n27550, n27552, n27554, n27556, n27558,
n27560, n27562, n27564, n27566, n27568, n27570, n27572, n27574,
n27576, n27578, n27580, n27582, n27584, n27586, n27588, n27590,
n27592, n27594, n27596, n27598, n27600, n27602, n27604, n27606,
n27608, n27610, n27612, n27614, n27616, n27618, n27620, n27622,
n27624, n27626, n27628, n27630, n27632, n27634, n27636, n27638,
n27640, n27642, n27644, n27646, n27648, n27650, n27652, n27654,
n27656, n27658, n27660, n27662, n27664, n27666, n27668, n27670,
n27672, n27674, n27676, n27678, n27680, n27682, n27684, n27686,
n27688, n27690, n27692, n27694, n27696, n27698, n27700, n27702,
n27704, n27706, n27708, n27710, n27712, n27714, n27716, n27718,
n27720, n27722, n27724, n27726, n27728, n27730, n27732, n27734,
n27736, n27738, n27740, n27742, n27744, n27746, n27748, n27750,
n27752, n27754, n27756, n27758, n27760, n27762, n27764, n27766,
n27768, n27770, n27772, n27774, n27776, n27778, n27780, n27782,
n27784, n27786, n27788, n27790, n27792, n27794, n27796, n27798,
n27800, n27802, n27804, n27806, n27808, n27810, n27812, n27814,
n27816, n27818, n27820, n27822, n27824, n27826, n27828, n27830,
n27832, n27834, n27836, n27838, n27840, n27842, n27844, n27846,
n27848, n27850, n27852, n27854, n27856, n27858, n27860, n27862,
n27864, n27866, n27868, n27870, n27872, n27874, n27876, n27878,
n27880, n27881, n27882, n27883, n27884, n27885, n27886, n27887,
n27888, n27889, n27890, n27891, n27892, n27893, n27894, n27895,
n27896, n27897, n27898, n27899, n27901, n27903, n27905, n27907,
n27909, n27911, n27913, n27915, n27917, n27919, n27921, n27923,
n27925, n27927, n27929, n27931, n27933, n27935, n27937, n27939,
n27941, n27943, n27945, n27947, n27949, n27951, n27953, n27955,
n27957, n27959, n27961, n27963, n27965, n27967, n27969, n27971,
n27973, n27975, n27977, n27979, n27981, n27983, n27985, n27987,
n27989, n27991, n27993, n27995, n27997, n27999, n28001, n28003,
n28005, n28007, n28009, n28011, n28013, n28015, n28017, n28019,
n28021, n28023, n28025, n28027, n28029, n28031, n28033, n28035,
n28037, n28039, n28041, n28043, n28045, n28047, n28049, n28051,
n28053, n28055, n28057, n28059, n28061, n28063, n28065, n28067,
n28069, n28071, n28073, n28075, n28077, n28079, n28081, n28083,
n28085, n28087, n28089, n28090, n28091, n28092, n28093, n28094,
n28095, n28096, n28097, n28098, n28099, n28100, n28101, n28102,
n28103, n28104, n28105, n28106, n28107, n28108, n28109, n28110,
n28111, n28112, n28113, n28114, n28115, n28116, n28117, n28118,
n28119, n28120, n28121, n28122, n28123, n28124, n28125, n28126,
n28127, n28128, n28129, n28130, n28132, n28133, n28134, n28135,
n28136, n28137, n28138, n28139, n28140, n28141, n28142, n28143,
n28144, n28145, n28146, n28147, n28148, n28149, n28150, n28151,
n28152, n28153, n28154, n28155, n28156, n28157, n28158, n28159,
n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167,
n28168, n28169, n28170, n28171, n28172, n28173, n28174, n28175,
n28176, n28177, n28178, n28179, n28180, n28181, n28182, n28183,
n28184, n28185, n28186, n28188, n28189, n28190, n28191, n28192,
n28193, n28194, n28195, n28196, n28197, n28198, n28199, n28200,
n28201, n28202, n28203, n28204, n28205, n28206, n28207, n28208,
n28209, n28210, n28211, n28212, n28213, n28214, n28215, n28216,
n28217, n28218, n28219, n28220, n28221, n28222, n28223, n28224,
n28225, n28226, n28227, n28228, n28229, n28230, n28231, n28232,
n28233, n28234, n28235, n28236, n28237, n28238, n28239, n28240,
n28241, n28242, n28243, n28244, n28245, n28246, n28247, n28248,
n28249, n28250, n28251, n28252, n28253, n28254, n28255, n28256,
n28257, n28258, n28259, n28260, n28261, n28262, n28263, n28264,
n28265, n28266, n28267, n28268, n28269, n28270, n28271, n28272,
n28273, n28274, n28275, n28276, n28277, n28278, n28279, n28280,
n28281, n28282, n28283, n28284, n28285, n28286, n28287, n28288,
n28289, n28290, n28291, n28292, n28293, n28294, n28295, n28296,
n28297, n28298, n28299, n28300, n28301, n28302, n28303, n28304,
n28305, n28306, n28307, n28308, n28309, n28310, n28311, n28312,
n28313, n28314, n28315, n28316, n28317, n28318, n28319, n28320,
n28321, n28322, n28323, n28324, n28325, n28326, n28327, n28328,
n28329, n28330, n28331, n28332, n28333, n28334, n28335, n28336,
n28337, n28338, n28339, n28340, n28341, n28342, n28343, n28344,
n28345, n28346, n28347, n28348, n28349, n28350, n28351, n28352,
n28353, n28354, n28355, n28356, n28357, n28358, n28359, n28360,
n28361, n28362, n28363, n28364, n28365, n28366, n28367, n28368,
n28369, n28370, n28371, n28372, n28373, n28374, n28375, n28376,
n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384,
n28385, n28386, n28387, n28388, n28389, n28390, n28391, n28392,
n28393, n28394, n28395, n28396, n28397, n28398, n28399, n28400,
n28401, n28402, n28403, n28404, n28405, n28406, n28407, n28408,
n28409, n28410, n28411, n28412, n28413, n28414, n28415, n28416,
n28417, n28418, n28419, n28420, n28421, n28422, n28423, n28424,
n28425, n28426, n28427, n28428, n28429, n28430, n28431, n28432,
n28433, n28434, n28435, n28436, n28437, n28438, n28439, n28440,
n28441, n28442, n28443, n28444, n28445, n28446, n28447, n28448,
n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456,
n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464,
n28465, n28466, n28467, n28468, n28469, n28470, n28471, n28472,
n28473, n28474, n28475, n28476, n28477, n28478, n28479, n28480,
n28481, n28482, n28483, n28484, n28485, n28486, n28487, n28488,
n28489, n28490, n28491, n28492, n28493, n28494, n28495, n28496,
n28497, n28498, n28499, n28500, n28501, n28502, n28503, n28504,
n28505, n28506, n28507, n28508, n28509, n28510, n28511, n28512,
n28513, n28514, n28515, n28516, n28517, n28518, n28519, n28520,
n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528,
n28529, n28530, n28531, n28532, n28533, n28534, n28535, n28536,
n28537, n28538, n28539, n28540, n28541, n28542, n28543, n28544,
n28545, n28546, n28547, n28548, n28549, n28550, n28551, n28552,
n28553, n28554, n28555, n28556, n28557, n28558, n28559, n28560,
n28561, n28562, n28563, n28564, n28565, n28566, n28567, n28568,
n28569, n28570, n28571, n28572, n28573, n28574, n28575, n28576,
n28577, n28578, n28579, n28580, n28581, n28582, n28583, n28584,
n28585, n28586, n28587, n28588, n28589, n28590, n28591, n28592,
n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600,
n28601, n28602, n28603, n28604, n28605, n28606, n28607, n28608,
n28609, n28610, n28611, n28612, n28613, n28614, n28615, n28616,
n28617, n28618, n28619, n28620, n28621, n28622, n28623, n28624,
n28625, n28626, n28627, n28628, n28629, n28630, n28631, n28632,
n28633, n28634, n28635, n28636, n28637, n28638, n28639, n28640,
n28641, n28642, n28643, n28644, n28645, n28646, n28647, n28648,
n28649, n28650, n28651, n28652, n28653, n28654, n28655, n28656,
n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664,
n28665, n28666, n28667, n28668, n28669, n28670, n28671, n28672,
n28673, n28674, n28675, n28676, n28677, n28678, n28679, n28680,
n28681, n28682, n28683, n28684, n28685, n28686, n28687, n28688,
n28689, n28690, n28691, n28692, n28693, n28694, n28695, n28696,
n28697, n28698, n28699, n28700, n28701, n28702, n28703, n28704,
n28705, n28706, n28707, n28708, n28709, n28710, n28711, n28712,
n28713, n28714, n28715, n28716, n28717, n28718, n28719, n28720,
n28721, n28722, n28723, n28724, n28725, n28726, n28727, n28728,
n28729, n28730, n28731, n28732, n28733, n28734, n28735, n28736,
n28737, n28738, n28739, n28740, n28741, n28742, n28743, n28744,
n28745, n28746, n28747, n28748, n28749, n28750, n28751, n28752,
n28753, n28754, n28755, n28756, n28757, n28758, n28759, n28760,
n28761, n28762, n28763, n28764, n28765, n28766, n28767, n28768,
n28769, n28770, n28771, n28772, n28773, n28774, n28775, n28776,
n28777, n28778, n28779, n28780, n28781, n28782, n28783, n28784,
n28785, n28786, n28787, n28788, n28789, n28790, n28791, n28792,
n28793, n28794, n28795, n28796, n28797, n28798, n28799, n28800,
n28801, n28802, n28803, n28804, n28805, n28806, n28807, n28808,
n28809, n28810, n28811, n28812, n28813, n28814, n28815, n28816,
n28817, n28818, n28819, n28820, n28821, n28822, n28823, n28824,
n28825, n28826, n28827, n28828, n28829, n28830, n28831, n28832,
n28833, n28834, n28835, n28836, n28837, n28838, n28839, n28840,
n28841, n28842, n28843, n28844, n28845, n28846, n28847, n28848,
n28849, n28850, n28851, n28852, n28853, n28854, n28855, n28856,
n28857, n28858, n28859, n28860, n28861, n28862, n28863, n28864,
n28865, n28866, n28867, n28868, n28869, n28870, n28871, n28872,
n28873, n28874, n28875, n28876, n28877, n28878, n28879, n28880,
n28881, n28882, n28883, n28884, n28885, n28886, n28887, n28888,
n28889, n28890, n28891, n28892, n28893, n28894, n28895, n28896,
n28897, n28898, n28899, n28900, n28901, n28902, n28903, n28904,
n28905, n28906, n28907, n28908, n28909, n28910, n28911, n28912,
n28913, n28914, n28915, n28916, n28917, n28918, n28919, n28920,
n28921, n28922, n28923, n28924, n28925, n28926, n28927, n28928,
n28929, n28930, n28931, n28932, n28933, n28934, n28935, n28936,
n28937, n28938, n28939, n28940, n28941, n28942, n28943, n28944,
n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952,
n28953, n28954, n28955, n28956, n28957, n28958, n28959, n28960,
n28961, n28962, n28963, n28964, n28965, n28966, n28967, n28968,
n28969, n28970, n28971, n28972, n28973, n28974, n28975, n28976,
n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984,
n28985, n28986, n28987, n28988, n28989, n28990, n28991, n28992,
n28993, n28994, n28995, n28996, n28997, n28998, n28999, n29000,
n29001, n29002, n29003, n29004, n29005, n29006, n29007, n29008,
n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016,
n29017, n29018, n29019, n29020, n29021, n29022, n29023, n29024,
n29025, n29026, n29027, n29028, n29029, n29030, n29031, n29032,
n29033, n29034, n29035, n29036, n29037, n29038, n29039, n29040,
n29041, n29042, n29043, n29044, n29045, n29046, n29047, n29048,
n29049, n29050, n29051, n29052, n29053, n29054, n29055, n29056,
n29057, n29058, n29059, n29060, n29061, n29062, n29063, n29064,
n29065, n29066, n29067, n29068, n29069, n29070, n29071, n29072,
n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080,
n29081, n29082, n29083, n29084, n29085, n29086, n29087, n29088,
n29089, n29090, n29091, n29092, n29093, n29094, n29095, n29096,
n29097, n29098, n29099, n29100, n29101, n29102, n29103, n29104,
n29105, n29106, n29107, n29108, n29109, n29110, n29111, n29112,
n29113, n29114, n29115, n29116, n29117, n29118, n29119, n29120,
n29121, n29122, n29123, n29124, n29125, n29126, n29127, n29128,
n29129, n29130, n29131, n29132, n29133, n29134, n29135, n29136,
n29137, n29138, n29139, n29140, n29141, n29142, n29143, n29144,
n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152,
n29153, n29154, n29155, n29156, n29157, n29158, n29159, n29160,
n29161, n29162, n29163, n29164, n29165, n29166, n29167, n29168,
n29169, n29170, n29171, n29172, n29173, n29174, n29175, n29176,
n29177, n29178, n29179, n29180, n29181, n29182, n29183, n29184,
n29185, n29186, n29187, n29188, n29189, n29190, n29191, n29192,
n29193, n29194, n29195, n29196, n29197, n29198, n29199, n29200,
n29201, n29202, n29203, n29204, n29205, n29206, n29207, n29208,
n29209, n29210, n29211, n29212, n29213, n29214, n29215, n29216,
n29217, n29218, n29219, n29220, n29221, n29222, n29223, n29224,
n29225, n29226, n29227, n29228, n29229, n29230, n29231, n29232,
n29233, n29234, n29235, n29236, n29237, n29238, n29239, n29240,
n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248,
n29249, n29250, n29251, n29252, n29253, n29254, n29255, n29256,
n29257, n29258, n29259, n29260, n29261, n29262, n29263, n29264,
n29265, n29266, n29267, n29268, n29269, n29270, n29271, n29272,
n29273, n29274, n29275, n29276, n29277, n29278, n29279, n29280,
n29281, n29282, n29283, n29284, n29285, n29286, n29287, n29288,
n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296,
n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304,
n29305, n29306, n29307, n29308, n29309, n29310, n29311, n29312,
n29313, n29314, n29315, n29316, n29317, n29318, n29319, n29320,
n29321, n29322, n29323, n29324, n29325, n29326, n29327, n29328,
n29329, n29330, n29331, n29332, n29333, n29334, n29335, n29336,
n29337, n29338, n29339, n29340, n29341, n29342, n29343, n29344,
n29345, n29346, n29347, n29348, n29349, n29350, n29351, n29352,
n29353, n29354, n29355, n29356, n29357, n29358, n29359, n29360,
n29361, n29362, n29363, n29364, n29365, n29366, n29367, n29368,
n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376,
n29377, n29378, n29379, n29380, n29381, n29382, n29383, n29384,
n29385, n29386, n29387, n29388, n29389, n29390, n29391, n29392,
n29393, n29394, n29395, n29396, n29397, n29398, n29399, n29400,
n29401, n29402, n29403, n29404, n29405, n29406, n29407, n29408,
n29409, n29410, n29411, n29412, n29413, n29414, n29415, n29416,
n29417, n29418, n29419, n29420, n29421, n29422, n29423, n29424,
n29425, n29426, n29427, n29428, n29429, n29430, n29431, n29432,
n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440,
n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448,
n29449, n29450, n29451, n29452, n29453, n29454, n29455, n29456,
n29457, n29458, n29459, n29460, n29461, n29462, n29463, n29464,
n29465, n29466, n29467, n29468, n29469, n29470, n29471, n29472,
n29473, n29474, n29475, n29476, n29477, n29478, n29479, n29480,
n29481, n29482, n29483, n29484, n29485, n29486, n29487, n29488,
n29489, n29490, n29491, n29492, n29493, n29494, n29495, n29496,
n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504,
n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512,
n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520,
n29521, n29522, n29523, n29524, n29525, n29526, n29527, n29528,
n29529, n29530, n29531, n29532, n29533, n29534, n29535, n29536,
n29537, n29538, n29539, n29540, n29541, n29542, n29543, n29544,
n29545, n29546, n29547, n29548, n29549, n29550, n29551, n29552,
n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560,
n29561, n29562, n29563, n29564, n29565, n29566, n29567, n29568,
n29569, n29570, n29571, n29572, n29573, n29574, n29575, n29576,
n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584,
n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592,
n29593, n29594, n29595, n29596, n29597, n29598, n29599, n29600,
n29601, n29602, n29603, n29604, n29605, n29606, n29607, n29608,
n29609, n29610, n29611, n29612, n29613, n29614, n29615, n29616,
n29617, n29618, n29619, n29620, n29621, n29622, n29623, n29624,
n29625, n29626, n29627, n29628, n29629, n29630, n29631, n29632,
n29633, n29634, n29635, n29636, n29637, n29638, n29639, n29640,
n29641, n29642, n29643, n29644, n29645, n29646, n29647, n29648,
n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656,
n29657, n29658, n29659, n29660, n29661, n29662, n29663, n29664,
n29665, n29666, n29667, n29668, n29669, n29670, n29671, n29672,
n29673, n29674, n29675, n29676, n29677, n29678, n29679, n29680,
n29681, n29682, n29683, n29684, n29685, n29686, n29687, n29688,
n29689, n29690, n29691, n29692, n29693, n29694, n29695, n29696,
n29697, n29698, n29699, n29700, n29701, n29702, n29703, n29704,
n29705, n29706, n29707, n29708, n29709, n29710, n29711, n29712,
n29713, n29714, n29715, n29716, n29717, n29718, n29719, n29720,
n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728,
n29729, n29730, n29731, n29732, n29733, n29734, n29735, n29736,
n29737, n29738, n29739, n29740, n29741, n29742, n29743, n29744,
n29745, n29746, n29747, n29748, n29749, n29750, n29751, n29752,
n29753, n29754, n29755, n29756, n29757, n29758, n29759, n29760,
n29761, n29762, n29763, n29764, n29765, n29766, n29767, n29768,
n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776,
n29777, n29778, n29779, n29780, n29781, n29782, n29783, n29784,
n29785, n29786, n29787, n29788, n29789, n29790, n29791, n29792,
n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800,
n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808,
n29809, n29810, n29811, n29812, n29813, n29814, n29815, n29816,
n29817, n29818, n29819, n29820, n29821, n29822, n29823, n29824,
n29825, n29826, n29827, n29828, n29829, n29830, n29831, n29832,
n29833, n29834, n29835, n29836, n29837, n29838, n29839, n29840,
n29841, n29842, n29843, n29844, n29845, n29846, n29847, n29848,
n29849, n29850, n29851, n29852, n29853, n29854, n29855, n29856,
n29857, n29858, n29859, n29860, n29861, n29862, n29863, n29864,
n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872,
n29873, n29874, n29875, n29876, n29877, n29878, n29879, n29880,
n29881, n29882, n29883, n29884, n29885, n29886, n29887, n29888,
n29889, n29890, n29891, n29892, n29893, n29894, n29895, n29896,
n29897, n29898, n29899, n29900, n29901, n29902, n29903, n29904,
n29905, n29906, n29907, n29908, n29909, n29910, n29911, n29912,
n29913, n29914, n29915, n29916, n29917, n29918, n29919, n29920,
n29921, n29922, n29923, n29924, n29925, n29926, n29927, n29928,
n29929, n29930, n29931, n29932, n29933, n29934, n29935, n29936,
n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944,
n29945, n29946, n29947, n29948, n29949, n29950, n29951, n29952,
n29953, n29954, n29955, n29956, n29957, n29958, n29959, n29960,
n29961, n29962, n29963, n29964, n29965, n29966, n29967, n29968,
n29969, n29970, n29971, n29972, n29973, n29974, n29975, n29976,
n29977, n29978, n29979, n29980, n29981, n29982, n29983, n29984,
n29985, n29986, n29987, n29988, n29989, n29990, n29991, n29992,
n29993, n29994, n29995, n29996, n29997, n29998, n29999, n30000,
n30001, n30002, n30003, n30004, n30005, n30006, n30007, n30008,
n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016,
n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024,
n30025, n30026, n30027, n30028, n30029, n30030, n30031, n30032,
n30033, n30034, n30035, n30036, n30037, n30038, n30039, n30040,
n30041, n30042, n30043, n30044, n30045, n30046, n30047, n30048,
n30049, n30050, n30051, n30052, n30053, n30054, n30055, n30056,
n30057, n30058, n30059, n30060, n30061, n30062, n30063, n30064,
n30065, n30066, n30067, n30068, n30069, n30070, n30071, n30072,
n30073, n30074, n30075, n30076, n30077, n30078, n30079, n30080,
n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088,
n30089, n30090, n30091, n30092, n30093, n30094, n30095, n30096,
n30097, n30098, n30099, n30100, n30101, n30102, n30103, n30104,
n30105, n30106, n30107, n30108, n30109, n30110, n30111, n30112,
n30113, n30114, n30115, n30116, n30117, n30118, n30119, n30120,
n30121, n30122, n30123, n30124, n30125, n30126, n30127, n30128,
n30129, n30130, n30131, n30132, n30133, n30134, n30135, n30136,
n30137, n30138, n30139, n30140, n30141, n30142, n30143, n30144,
n30145, n30146, n30147, n30148, n30149, n30150, n30151, n30152,
n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160,
n30161, n30162, n30163, n30164, n30165, n30166, n30167, n30168,
n30169, n30170, n30171, n30172, n30173, n30174, n30175, n30176,
n30177, n30178, n30179, n30180, n30181, n30182, n30183, n30184,
n30185, n30186, n30187, n30188, n30189, n30190, n30191, n30192,
n30193, n30194, n30195, n30196, n30197, n30198, n30199, n30200,
n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208,
n30209, n30210, n30211, n30212, n30213, n30214, n30215, n30216,
n30217, n30218, n30219, n30220, n30221, n30222, n30223, n30224,
n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232,
n30233, n30234, n30235, n30236, n30237, n30238, n30239, n30240,
n30241, n30242, n30243, n30244, n30245, n30246, n30247, n30248,
n30249, n30250, n30251, n30252, n30253, n30254, n30255, n30256,
n30257, n30258, n30259, n30260, n30261, n30262, n30263, n30264,
n30265, n30266, n30267, n30268, n30269, n30270, n30271, n30272,
n30273, n30274, n30275, n30276, n30277, n30278, n30279, n30280,
n30281, n30282, n30283, n30284, n30285, n30286, n30287, n30288,
n30289, n30290, n30291, n30292, n30293, n30294, n30295, n30296,
n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304,
n30305, n30306, n30307, n30308, n30309, n30310, n30311, n30312,
n30313, n30314, n30315, n30316, n30317, n30318, n30319, n30320,
n30321, n30322, n30323, n30324, n30325, n30326, n30327, n30328,
n30329, n30330, n30331, n30332, n30333, n30334, n30335, n30336,
n30337, n30338, n30339, n30340, n30341, n30342, n30343, n30344,
n30345, n30346, n30347, n30348, n30349, n30350, n30351, n30352,
n30353, n30354, n30355, n30356, n30357, n30358, n30359, n30360,
n30361, n30362, n30363, n30364, n30365, n30366, n30367, n30368,
n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376,
n30377, n30378, n30379, n30380, n30381, n30382, n30383, n30384,
n30385, n30386, n30387, n30388, n30389, n30390, n30391, n30392,
n30393, n30394, n30395, n30396, n30397, n30398, n30399, n30400,
n30401, n30402, n30403, n30404, n30405, n30406, n30407, n30408,
n30409, n30410, n30411, n30412, n30413, n30414, n30415, n30416,
n30417, n30418, n30419, n30420, n30421, n30422, n30423, n30424,
n30425, n30426, n30427, n30428, n30429, n30430, n30431, n30432,
n30433, n30434, n30435, n30436, n30437, n30438, n30439, n30440,
n30441, n30442, n30443, n30444, n30445, n30446, n30447, n30448,
n30449, n30450, n30451, n30452, n30453, n30454, n30455, n30456,
n30457, n30458, n30459, n30460, n30461, n30462, n30463, n30464,
n30465, n30466, n30467, n30468, n30469, n30470, n30471, n30472,
n30473, n30474, n30475, n30476, n30477, n30478, n30479, n30480,
n30481, n30482, n30483, n30484, n30485, n30486, n30487, n30488,
n30489, n30490, n30491, n30492, n30493, n30494, n30495, n30496,
n30497, n30498, n30499, n30500, n30501, n30502, n30503, n30504,
n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512,
n30513, n30514, n30515, n30516, n30517, n30518, n30519, n30520,
n30521, n30522, n30523, n30524, n30525, n30526, n30527, n30528,
n30529, n30530, n30531, n30532, n30533, n30534, n30535, n30536,
n30537, n30538, n30539, n30540, n30541, n30542, n30543, n30544,
n30545, n30546, n30547, n30548, n30549, n30550, n30551, n30552,
n30553, n30554, n30555, n30556, n30557, n30558, n30559, n30560,
n30561, n30562, n30563, n30564, n30565, n30566, n30567, n30568,
n30569, n30570, n30571, n30572, n30573, n30574, n30575, n30576,
n30577, n30578, n30579, n30580, n30581, n30582, n30583, n30584,
n30585, n30586, n30587, n30588, n30589, n30590, n30591, n30592,
n30593, n30594, n30595, n30596, n30597, n30598, n30599, n30600,
n30601, n30602, n30603, n30604, n30605, n30606, n30607, n30608,
n30609, n30610, n30611, n30612, n30613, n30614, n30615, n30616,
n30617, n30618, n30619, n30620, n30621, n30622, n30623, n30624,
n30625, n30626, n30627, n30628, n30629, n30630, n30631, n30632,
n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640,
n30641, n30642, n30643, n30644, n30645, n30646, n30647, n30648,
n30649, n30650, n30651, n30652, n30653, n30654, n30655, n30656,
n30657, n30658, n30659, n30660, n30661, n30662, n30663, n30664,
n30665, n30666, n30667, n30668, n30669, n30670, n30671, n30672,
n30673, n30674, n30675, n30676, n30677, n30678, n30679, n30680,
n30681, n30682, n30683, n30684, n30685, n30686, n30687, n30688,
n30689, n30690, n30691, n30692, n30693, n30694, n30695, n30696,
n30697, n30698, n30699, n30700, n30701, n30702, n30703, n30704,
n30705, n30706, n30707, n30708, n30709, n30710, n30711, n30712,
n30713, n30714, n30715, n30716, n30717, n30718, n30719, n30720,
n30721, n30722, n30723, n30724, n30725, n30726, n30727, n30728,
n30729, n30730, n30731, n30732, n30733, n30734, n30735, n30736,
n30737, n30738, n30739, n30740, n30741, n30742, n30743, n30744,
n30745, n30746, n30747, n30748, n30749, n30750, n30751, n30752,
n30753, n30754, n30755, n30756, n30757, n30758, n30759, n30760,
n30761, n30762, n30763, n30764, n30765, n30766, n30767, n30768,
n30769, n30770, n30771, n30772, n30773, n30774, n30775, n30776,
n30777, n30778, n30779, n30780, n30781, n30782, n30783, n30784,
n30785, n30786, n30787, n30788, n30789, n30790, n30791, n30792,
n30793, n30794, n30795, n30796, n30797, n30798, n30799, n30800,
n30801, n30802, n30803, n30804, n30805, n30806, n30807, n30808,
n30809, n30810, n30811, n30812, n30813, n30814, n30815, n30816,
n30817, n30818, n30819, n30820, n30821, n30822, n30823, n30824,
n30825, n30826, n30827, n30828, n30829, n30830, n30831, n30832,
n30833, n30834, n30835, n30836, n30837, n30838, n30839, n30840,
n30841, n30842, n30843, n30844, n30845, n30846, n30847, n30848,
n30849, n30850, n30851, n30852, n30853, n30854, n30855, n30856,
n30857, n30858, n30859, n30860, n30861, n30862, n30863, n30864,
n30865, n30866, n30867, n30868, n30869, n30870, n30871, n30872,
n30873, n30874, n30875, n30876, n30877, n30878, n30879, n30880,
n30881, n30882, n30883, n30884, n30885, n30886, n30887, n30888,
n30889, n30890, n30891, n30892, n30893, n30894, n30895, n30896,
n30897, n30898, n30899, n30900, n30901, n30902, n30903, n30904,
n30905, n30906, n30907, n30908, n30909, n30910, n30911, n30912,
n30913, n30914, n30915, n30916, n30917, n30918, n30919, n30920,
n30921, n30922, n30923, n30924, n30925, n30926, n30927, n30928,
n30929, n30930, n30931, n30932, n30933, n30934, n30935, n30936,
n30937, n30938, n30939, n30940, n30941, n30942, n30943, n30944,
n30945, n30946, n30947, n30948, n30949, n30950, n30951, n30952,
n30953, n30954, n30955, n30956, n30957, n30958, n30959, n30960,
n30961, n30962, n30963, n30964, n30965, n30966, n30967, n30968,
n30969, n30970, n30971, n30972, n30973, n30974, n30975, n30976,
n30977, n30978, n30979, n30980, n30981, n30982, n30983, n30984,
n30985, n30986, n30987, n30988, n30989, n30990, n30991, n30992,
n30993, n30994, n30995, n30996, n30997, n30998, n30999, n31000,
n31001, n31002, n31003, n31004, n31005, n31006, n31007, n31008,
n31009, n31010, n31011, n31012, n31013, n31014, n31015, n31016,
n31017, n31018, n31019, n31020, n31021, n31022, n31023, n31024,
n31025, n31026, n31027, n31028, n31029, n31030, n31031, n31032,
n31033, n31034, n31035, n31036, n31037, n31038, n31039, n31040,
n31041, n31042, n31043, n31044, n31045, n31046, n31047, n31048,
n31049, n31050, n31051, n31052, n31053, n31054, n31055, n31056,
n31057, n31058, n31059, n31060, n31061, n31062, n31063, n31064,
n31065, n31066, n31067, n31068, n31069, n31070, n31071, n31072,
n31073, n31074, n31075, n31076, n31077, n31078, n31079, n31080,
n31081, n31082, n31083, n31084, n31085, n31086, n31087, n31088,
n31089, n31090, n31091, n31092, n31093, n31094, n31095, n31096,
n31097, n31098, n31099, n31100, n31101, n31102, n31103, n31104,
n31105, n31106, n31107, n31108, n31109, n31110, n31111, n31112,
n31113, n31114, n31115, n31116, n31117, n31118, n31119, n31120,
n31121, n31122, n31123, n31124, n31125, n31126, n31127, n31128,
n31129, n31130, n31131, n31132, n31133, n31134, n31135, n31136,
n31137, n31138, n31139, n31140, n31141, n31142, n31143, n31144,
n31145, n31146, n31147, n31148, n31149, n31150, n31151, n31152,
n31153, n31154, n31155, n31156, n31157, n31158, n31159, n31160,
n31161, n31162, n31163, n31164, n31165, n31166, n31167, n31168,
n31169, n31170, n31171, n31172, n31173, n31174, n31175, n31176,
n31177, n31178, n31179, n31180, n31181, n31182, n31183, n31184,
n31185, n31186, n31187, n31188, n31189, n31190, n31191, n31192,
n31193, n31194, n31195, n31196, n31197, n31198, n31199, n31200,
n31201, n31202, n31203, n31204, n31205, n31206, n31207, n31208,
n31209, n31210, n31211, n31212, n31213, n31214, n31215, n31216,
n31217, n31218, n31219, n31220, n31221, n31222, n31223, n31224,
n31225, n31226, n31227, n31228, n31229, n31230, n31231, n31232,
n31233, n31234, n31235, n31236, n31237, n31238, n31239, n31240,
n31241, n31242, n31243, n31244, n31245, n31246, n31247, n31248,
n31249, n31250, n31251, n31252, n31253, n31254, n31255, n31256,
n31257, n31258, n31259, n31260, n31261, n31262, n31263, n31264,
n31265, n31266, n31267, n31268, n31269, n31270, n31271, n31272,
n31273, n31274, n31275, n31276, n31277, n31278, n31279, n31280,
n31281, n31282, n31283, n31284, n31285, n31286, n31287, n31288,
n31289, n31290, n31291, n31292, n31293, n31294, n31295, n31296,
n31297, n31298, n31299, n31300, n31301, n31302, n31303, n31304,
n31305, n31306, n31307, n31308, n31309, n31310, n31311, n31312,
n31313, n31314, n31315, n31316, n31317, n31318, n31319, n31320,
n31321, n31322, n31323, n31324, n31325, n31326, n31327, n31328,
n31329, n31330, n31331, n31332, n31333, n31334, n31335, n31336,
n31337, n31338, n31339, n31340, n31341, n31342, n31343, n31344,
n31345, n31346, n31347, n31348, n31349, n31350, n31351, n31352,
n31353, n31354, n31355, n31356, n31357, n31358, n31359, n31360,
n31361, n31362, n31363, n31364, n31365, n31366, n31367, n31368,
n31369, n31370, n31371, n31372, n31373, n31374, n31375, n31376,
n31377, n31378, n31379, n31380, n31381, n31382, n31383, n31384,
n31385, n31386, n31387, n31388, n31389, n31390, n31391, n31392,
n31393, n31394, n31395, n31396, n31397, n31398, n31399, n31400,
n31401, n31402, n31403, n31404, n31405, n31406, n31407, n31408,
n31409, n31410, n31411, n31412, n31413, n31414, n31415, n31416,
n31417, n31418, n31419, n31420, n31421, n31422, n31423, n31424,
n31425, n31426, n31427, n31428, n31429, n31430, n31431, n31432,
n31433, n31434, n31435, n31436, n31437, n31438, n31439, n31440,
n31441, n31442, n31443, n31444, n31445, n31446, n31447, n31448,
n31449, n31450, n31451, n31452, n31453, n31454, n31455, n31456,
n31457, n31458, n31459, n31460, n31461, n31462, n31463, n31464,
n31465, n31466, n31467, n31468, n31469, n31470, n31471, n31472,
n31473, n31474, n31475, n31476, n31477, n31478, n31479, n31480,
n31481, n31482, n31483, n31484, n31485, n31486, n31487, n31488,
n31489, n31490, n31491, n31492, n31493, n31494, n31495, n31496,
n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504,
n31505, n31506, n31507, n31508, n31509, n31510, n31511, n31512,
n31513, n31514, n31515, n31516, n31517, n31518, n31519, n31520,
n31521, n31522, n31523, n31524, n31525, n31526, n31527, n31528,
n31529, n31530, n31531, n31532, n31533, n31534, n31535, n31536,
n31537, n31538, n31539, n31540, n31541, n31542, n31543, n31544,
n31545, n31546, n31547, n31548, n31549, n31550, n31551, n31552,
n31553, n31554, n31555, n31556, n31557, n31558, n31559, n31560,
n31561, n31562, n31563, n31564, n31565, n31566, n31567, n31568,
n31569, n31570, n31571, n31572, n31573, n31574, n31575, n31576,
n31577, n31578, n31579, n31580, n31581, n31582, n31583, n31584,
n31585, n31586, n31587, n31588, n31589, n31590, n31591, n31592,
n31593, n31594, n31595, n31596, n31597, n31598, n31599, n31600,
n31601, n31602, n31603, n31604, n31605, n31606, n31607, n31608,
n31609, n31610, n31611, n31612, n31613, n31614, n31615, n31616,
n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624,
n31625, n31626, n31627, n31628, n31629, n31630, n31631, n31632,
n31633, n31634, n31635, n31636, n31637, n31638, n31639, n31640,
n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31648,
n31649, n31650, n31651, n31652, n31653, n31654, n31655, n31656,
n31657, n31658, n31659, n31660, n31661, n31662, n31663, n31664,
n31665, n31666, n31667, n31668, n31669, n31670, n31671, n31672,
n31673, n31674, n31675, n31676, n31677, n31678, n31679, n31680,
n31681, n31682, n31683, n31684, n31685, n31686, n31687, n31688,
n31689, n31690, n31691, n31692, n31693, n31694, n31695, n31696,
n31697, n31698, n31699, n31700, n31701, n31702, n31703, n31704,
n31705, n31706, n31707, n31708, n31709, n31710, n31711, n31712,
n31713, n31714, n31715, n31716, n31717, n31718, n31719, n31720,
n31721, n31722, n31723, n31724, n31725, n31726, n31727, n31728,
n31729, n31730, n31731, n31732, n31733, n31734, n31735, n31736,
n31737, n31738, n31739, n31740, n31741, n31742, n31743, n31744,
n31745, n31746, n31747, n31748, n31749, n31750, n31751, n31752,
n31753, n31754, n31755, n31756, n31757, n31758, n31759, n31760,
n31761, n31762, n31763, n31764, n31765, n31766, n31767, n31768,
n31769, n31770, n31771, n31772, n31773, n31774, n31775, n31776,
n31777, n31778, n31779, n31780, n31781, n31782, n31783, n31784,
n31785, n31786, n31787, n31788, n31789, n31790, n31791, n31792,
n31793, n31794, n31795, n31796, n31797, n31798, n31799, n31800,
n31801, n31802, n31803, n31804, n31805, n31806, n31807, n31808,
n31809, n31810, n31811, n31812, n31813, n31814, n31815, n31816,
n31817, n31818, n31819, n31820, n31821, n31822, n31823, n31824,
n31825, n31826, n31827, n31828, n31829, n31830, n31831, n31832,
n31833, n31834, n31835, n31836, n31837, n31838, n31839, n31840,
n31841, n31842, n31843, n31844, n31845, n31846, n31847, n31848,
n31849, n31850, n31851, n31852, n31853, n31854, n31855, n31856,
n31857, n31858, n31859, n31860, n31861, n31862, n31863, n31864,
n31865, n31866, n31867, n31868, n31869, n31870, n31871, n31872,
n31873, n31874, n31875, n31876, n31877, n31878, n31879, n31880,
n31881, n31882, n31883, n31884, n31885, n31886, n31887, n31888,
n31889, n31890, n31891, n31892, n31893, n31894, n31895, n31896,
n31897, n31898, n31899, n31900, n31901, n31902, n31903, n31904,
n31905, n31906, n31907, n31908, n31909, n31910, n31911, n31912,
n31913, n31914, n31915, n31916, n31917, n31918, n31919, n31920,
n31921, n31922, n31923, n31924, n31925, n31926, n31927, n31928,
n31929, n31930, n31931, n31932, n31933, n31934, n31935, n31936,
n31937, n31938, n31939, n31940, n31941, n31942, n31943, n31944,
n31945, n31946, n31947, n31948, n31949, n31950, n31951, n31952,
n31953, n31954, n31955, n31956, n31957, n31958, n31959, n31960,
n31961, n31962, n31963, n31964, n31965, n31966, n31967, n31968,
n31969, n31970, n31971, n31972, n31973, n31974, n31975, n31976,
n31977, n31978, n31979, n31980, n31981, n31982, n31983, n31984,
n31985, n31986, n31987, n31988, n31989, n31990, n31991, n31992,
n31993, n31994, n31995, n31996, n31997, n31998, n31999, n32000,
n32001, n32002, n32003, n32004, n32005, n32006, n32007, n32008,
n32009, n32010, n32011, n32012, n32013, n32014, n32015, n32016,
n32017, n32018, n32019, n32020, n32021, n32022, n32023, n32024,
n32025, n32026, n32027, n32028, n32029, n32030, n32031, n32032,
n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32040,
n32041, n32042, n32043, n32044, n32045, n32046, n32047, n32048,
n32049, n32050, n32051, n32052, n32053, n32054, n32055, n32056,
n32057, n32058, n32059, n32060, n32061, n32062, n32063, n32064,
n32065, n32066, n32067, n32068, n32069, n32070, n32071, n32072,
n32073, n32074, n32075, n32076, n32077, n32078, n32079, n32080,
n32081, n32082, n32083, n32084, n32085, n32086, n32087, n32088,
n32089, n32090, n32091, n32092, n32093, n32094, n32095, n32096,
n32097, n32098, n32099, n32100, n32101, n32102, n32103, n32104,
n32105, n32106, n32107, n32108, n32109, n32110, n32111, n32112,
n32113, n32114, n32115, n32116, n32117, n32118, n32119, n32120,
n32121, n32122, n32123, n32124, n32125, n32126, n32127, n32128,
n32129, n32130, n32131, n32132, n32133, n32134, n32135, n32136,
n32137, n32138, n32139, n32140, n32141, n32142, n32143, n32144,
n32145, n32146, n32147, n32148, n32149, n32150, n32151, n32152,
n32153, n32154, n32155, n32156, n32157, n32158, n32159, n32160,
n32161, n32162, n32163, n32164, n32165, n32166, n32167, n32168,
n32169, n32170, n32171, n32172, n32173, n32174, n32175, n32176,
n32177, n32178, n32179, n32180, n32181, n32182, n32183, n32184,
n32185, n32186, n32187, n32188, n32189, n32190, n32191, n32192,
n32193, n32194, n32195, n32196, n32197, n32198, n32199, n32200,
n32201, n32202, n32203, n32204, n32205, n32206, n32207, n32208,
n32209, n32210, n32211, n32212, n32213, n32214, n32215, n32216,
n32217, n32218, n32219, n32220, n32221, n32222, n32223, n32224,
n32225, n32226, n32227, n32228, n32229, n32230, n32231, n32232,
n32233, n32234, n32235, n32236, n32237, n32238, n32239, n32240,
n32241, n32242, n32243, n32244, n32245, n32246, n32247, n32248,
n32249, n32250, n32251, n32252, n32253, n32254, n32255, n32256,
n32257, n32258, n32259, n32260, n32261, n32262, n32263, n32264,
n32265, n32266, n32267, n32268, n32269, n32270, n32271, n32272,
n32273, n32274, n32275, n32276, n32277, n32278, n32279, n32280,
n32281, n32282, n32283, n32284, n32285, n32286, n32287, n32288,
n32289, n32290, n32291, n32292, n32293, n32294, n32295, n32296,
n32297, n32298, n32299, n32300, n32301, n32302, n32303, n32304,
n32305, n32306, n32307, n32308, n32309, n32310, n32311, n32312,
n32313, n32314, n32315, n32316, n32317, n32318, n32319, n32320,
n32321, n32322, n32323, n32324, n32325, n32326, n32327, n32328,
n32329, n32330, n32331, n32332, n32333, n32334, n32335, n32336,
n32337, n32338, n32339, n32340, n32341, n32342, n32343, n32344,
n32345, n32346, n32347, n32348, n32349, n32350, n32351, n32352,
n32353, n32354, n32355, n32356, n32357, n32358, n32359, n32360,
n32361, n32362, n32363, n32364, n32365, n32366, n32367, n32368,
n32369, n32370, n32371, n32372, n32373, n32374, n32375, n32376,
n32377, n32378, n32379, n32380, n32381, n32382, n32383, n32384,
n32385, n32386, n32387, n32388, n32389, n32390, n32391, n32392,
n32393, n32394, n32395, n32396, n32397, n32398, n32399, n32400,
n32401, n32402, n32403, n32404, n32405, n32406, n32407, n32408,
n32409, n32410, n32411, n32412, n32413, n32414, n32415, n32416,
n32417, n32418, n32419, n32420, n32421, n32422, n32423, n32424,
n32425, n32426, n32427, n32428, n32429, n32430, n32431, n32432,
n32433, n32434, n32435, n32436, n32437, n32438, n32439, n32440,
n32441, n32442, n32443, n32444, n32445, n32446, n32447, n32448,
n32449, n32450, n32451, n32452, n32453, n32454, n32455, n32456,
n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464,
n32465, n32466, n32467, n32468, n32469, n32470, n32471, n32472,
n32473, n32474, n32475, n32476, n32477, n32478, n32479, n32480,
n32481, n32482, n32483, n32484, n32485, n32486, n32487, n32488,
n32489, n32490, n32491, n32492, n32493, n32494, n32495, n32496,
n32497, n32498, n32499, n32500, n32501, n32502, n32503, n32504,
n32505, n32506, n32507, n32508, n32509, n32510, n32511, n32512,
n32513, n32514, n32515, n32516, n32517, n32518, n32519, n32520,
n32521, n32522, n32523, n32524, n32525, n32526, n32527, n32528,
n32529, n32530, n32531, n32532, n32533, n32534, n32535, n32536,
n32537, n32538, n32539, n32540, n32541, n32542, n32543, n32544,
n32545, n32546, n32547, n32548, n32549, n32550, n32551, n32552,
n32553, n32554, n32555, n32556, n32557, n32558, n32559, n32560,
n32561, n32562, n32563, n32564, n32565, n32566, n32567, n32568,
n32569, n32570, n32571, n32572, n32573, n32574, n32575, n32576,
n32577, n32578, n32579, n32580, n32581, n32582, n32583, n32584,
n32585, n32586, n32587, n32588, n32589, n32590, n32591, n32592,
n32593, n32594, n32595, n32596, n32597, n32598, n32599, n32600,
n32601, n32602, n32603, n32604, n32605, n32606, n32607, n32608,
n32609, n32610, n32611, n32612, n32613, n32614, n32615, n32616,
n32617, n32618, n32619, n32620, n32621, n32622, n32623, n32624,
n32625, n32626, n32627, n32628, n32629, n32630, n32631, n32632,
n32633, n32634, n32635, n32636, n32637, n32638, n32639, n32640,
n32641, n32642, n32643, n32644, n32645, n32646, n32647, n32648,
n32649, n32650, n32651, n32652, n32653, n32654, n32655, n32656,
n32657, n32658, n32659, n32660, n32661, n32662, n32663, n32664,
n32665, n32666, n32667, n32668, n32669, n32670, n32671, n32672,
n32673, n32674, n32675, n32676, n32677, n32678, n32679, n32680,
n32681, n32682, n32683, n32684, n32685, n32686, n32687, n32688,
n32689, n32690, n32691, n32692, n32693, n32694, n32695, n32696,
n32697, n32698, n32699, n32700, n32701, n32702, n32703, n32704,
n32705, n32706, n32707, n32708, n32709, n32710, n32711, n32712,
n32713, n32714, n32715, n32716, n32717, n32718, n32719, n32720,
n32721, n32722, n32723, n32724, n32725, n32726, n32727, n32728,
n32729, n32730, n32731, n32732, n32733, n32734, n32735, n32736,
n32737, n32738, n32739, n32740, n32741, n32742, n32743, n32744,
n32745, n32746, n32747, n32748, n32749, n32750, n32751, n32752,
n32753, n32754, n32755, n32756, n32757, n32758, n32759, n32760,
n32761, n32762, n32763, n32764, n32765, n32766, n32767, n32768,
n32769, n32770, n32771, n32772, n32773, n32774, n32775, n32776,
n32777, n32778, n32779, n32780, n32781, n32782, n32783, n32784,
n32785, n32786, n32787, n32788, n32789, n32790, n32791, n32792,
n32793, n32794, n32795, n32796, n32797, n32798, n32799, n32800,
n32801, n32802, n32803, n32804, n32805, n32806, n32807, n32808,
n32809, n32810, n32811, n32812, n32813, n32814, n32815, n32816,
n32817, n32818, n32819, n32820, n32821, n32822, n32823, n32824,
n32825, n32826, n32827, n32828, n32829, n32830, n32831, n32832,
n32833, n32834, n32835, n32836, n32837, n32838, n32839, n32840,
n32841, n32842, n32843, n32844, n32845, n32846, n32847, n32848,
n32849, n32850, n32851, n32852, n32853, n32854, n32855, n32856,
n32857, n32858, n32859, n32860, n32861, n32862, n32863, n32864,
n32865, n32866, n32867, n32868, n32869, n32870, n32871, n32872,
n32873, n32874, n32875, n32876, n32877, n32878, n32879, n32880,
n32881, n32882, n32883, n32884, n32885, n32886, n32887, n32888,
n32889, n32890, n32891, n32892, n32893, n32894, n32895, n32896,
n32897, n32898, n32899, n32900, n32901, n32902, n32903, n32904,
n32905, n32906, n32907, n32908, n32909, n32910, n32911, n32912,
n32913, n32914, n32915, n32916, n32917, n32918, n32919, n32920,
n32921, n32922, n32923, n32924, n32925, n32926, n32927, n32928,
n32929, n32930, n32931, n32932, n32933, n32934, n32935, n32936,
n32937, n32938, n32939, n32940, n32941, n32942, n32943, n32944,
n32945, n32946, n32947, n32948, n32949, n32950, n32951, n32952,
n32953, n32954, n32955, n32956, n32957, n32958, n32959, n32960,
n32961, n32962, n32963, n32964, n32965, n32966, n32967, n32968,
n32969, n32970, n32971, n32972, n32973, n32974, n32975, n32976,
n32977, n32978, n32979, n32980, n32981, n32982, n32983, n32984,
n32985, n32986, n32987, n32988, n32989, n32990, n32991, n32992,
n32993, n32994, n32995, n32996, n32997, n32998, n32999, n33000,
n33001, n33002, n33003, n33004, n33005, n33006, n33007, n33008,
n33009, n33010, n33011, n33012, n33013, n33014, n33015, n33016,
n33017, n33018, n33019, n33020, n33021, n33022, n33023, n33024,
n33025, n33026, n33027, n33028, n33029, n33030, n33031, n33032,
n33033, n33034, n33035, n33036, n33037, n33038, n33039, n33040,
n33041, n33042, n33043, n33044, n33045, n33046, n33047, n33048,
n33049, n33050, n33051, n33052, n33053, n33054, n33055, n33056,
n33057, n33058, n33059, n33060, n33061, n33062, n33063, n33064,
n33065, n33066, n33067, n33068, n33069, n33070, n33071, n33072,
n33073, n33074, n33075, n33076, n33077, n33078, n33079, n33080,
n33081, n33082, n33083, n33084, n33085, n33086, n33087, n33088,
n33089, n33090, n33091, n33092, n33093, n33094, n33095, n33096,
n33097, n33098, n33099, n33100, n33101, n33102, n33103, n33104,
n33105, n33106, n33107, n33108, n33109, n33110, n33111, n33112,
n33113, n33114, n33115, n33116, n33117, n33118, n33119, n33120,
n33121, n33122, n33123, n33124, n33125, n33126, n33127, n33128,
n33129, n33130, n33131, n33132, n33133, n33134, n33135, n33136,
n33137, n33138, n33139, n33140, n33141, n33142, n33143, n33144,
n33145, n33146, n33147, n33148, n33149, n33150, n33151, n33152,
n33153, n33154, n33155, n33156, n33157, n33158, n33159, n33160,
n33161, n33162, n33163, n33164, n33165, n33166, n33167, n33168,
n33169, n33170, n33171, n33172, n33173, n33174, n33175, n33176,
n33177, n33178, n33179, n33180, n33181, n33182, n33183, n33184,
n33185, n33186, n33187, n33188, n33189, n33190, n33191, n33192,
n33193, n33194, n33195, n33196, n33197, n33198, n33199, n33200,
n33201, n33202, n33203, n33204, n33205, n33206, n33207, n33208,
n33209, n33210, n33211, n33212, n33213, n33214, n33215, n33216,
n33217, n33218, n33219, n33220, n33221, n33222, n33223, n33224,
n33225, n33226, n33227, n33228, n33229, n33230, n33231, n33232,
n33233, n33234, n33235, n33236, n33237, n33238, n33239, n33240,
n33241, n33242, n33243, n33244, n33245, n33246, n33247, n33248,
n33249, n33250, n33251, n33252, n33253, n33254, n33255, n33256,
n33257, n33258, n33259, n33260, n33261, n33262, n33263, n33264,
n33265, n33266, n33267, n33268, n33269, n33270, n33271, n33272,
n33273, n33274, n33275, n33276, n33277, n33278, n33279, n33280,
n33281, n33282, n33283, n33284, n33285, n33286, n33287, n33288,
n33289, n33290, n33291, n33292, n33293, n33294, n33295, n33296,
n33297, n33298, n33299, n33300, n33301, n33302, n33303, n33304,
n33305, n33306, n33307, n33308, n33309, n33310, n33311, n33312,
n33313, n33314, n33315, n33316, n33317, n33318, n33319, n33320,
n33321, n33322, n33323, n33324, n33325, n33326, n33327, n33328,
n33329, n33330, n33331, n33332, n33333, n33334, n33335, n33336,
n33337, n33338, n33339, n33340, n33341, n33342, n33343, n33344,
n33345, n33346, n33347, n33348, n33349, n33350, n33351, n33352,
n33353, n33354, n33355, n33356, n33357, n33358, n33359, n33360,
n33361, n33362, n33363, n33364, n33365, n33366, n33367, n33368,
n33369, n33370, n33371, n33372, n33373, n33374, n33375, n33376,
n33377, n33378, n33379, n33380, n33381, n33382, n33383, n33384,
n33385, n33386, n33387, n33388, n33389, n33390, n33391, n33392,
n33393, n33394, n33395, n33396, n33397, n33398, n33399, n33400,
n33401, n33402, n33403, n33404, n33405, n33406, n33407, n33408,
n33409, n33410, n33411, n33412, n33413, n33414, n33415, n33416,
n33417, n33418, n33419, n33420, n33421, n33422, n33423, n33424,
n33425, n33426, n33427, n33428, n33429, n33430, n33431, n33432,
n33433, n33434, n33435, n33436, n33437, n33438, n33439, n33440,
n33441, n33442, n33443, n33444, n33445, n33446, n33447, n33448,
n33449, n33450, n33451, n33452, n33453, n33454, n33455, n33456,
n33457, n33458, n33459, n33460, n33461, n33462, n33463, n33464,
n33465, n33466, n33467, n33468, n33469, n33470, n33471, n33472,
n33473, n33474, n33475, n33476, n33477, n33478, n33479, n33480,
n33481, n33482, n33483, n33484, n33485, n33486, n33487, n33488,
n33489, n33490, n33491, n33492, n33493, n33494, n33495, n33496,
n33497, n33498, n33499, n33500, n33501, n33502, n33503, n33504,
n33505, n33506, n33507, n33508, n33509, n33510, n33511, n33512,
n33513, n33514, n33515, n33516, n33517, n33518, n33519, n33520,
n33521, n33522, n33523, n33524, n33525, n33526, n33527, n33528,
n33529, n33530, n33531, n33532, n33533, n33534, n33535, n33536,
n33537, n33538, n33539, n33540, n33541, n33542, n33543, n33544,
n33545, n33546, n33547, n33548, n33549, n33550, n33551, n33552,
n33553, n33554, n33555, n33556, n33557, n33558, n33559, n33560,
n33561, n33562, n33563, n33564, n33565, n33566, n33567, n33568,
n33569, n33570, n33571, n33572, n33573, n33574, n33575, n33576,
n33577, n33578, n33579, n33580, n33581, n33582, n33583, n33584,
n33585, n33586, n33587, n33588, n33589, n33590, n33591, n33592,
n33593, n33594, n33595, n33596, n33597, n33598, n33599, n33600,
n33601, n33602, n33603, n33604, n33605, n33606, n33607, n33608,
n33609, n33610, n33611, n33612, n33613, n33614, n33615, n33616,
n33617, n33618, n33619, n33620, n33621, n33622, n33623, n33624,
n33625, n33626, n33627, n33628, n33629, n33630, n33631, n33632,
n33633, n33634, n33635, n33636, n33637, n33638, n33639, n33640,
n33641, n33642, n33643, n33644, n33645, n33646, n33647, n33648,
n33649, n33650, n33651, n33652, n33653, n33654, n33655, n33656,
n33657, n33658, n33659, n33660, n33661, n33662, n33663, n33664,
n33665, n33666, n33667, n33668, n33669, n33670, n33671, n33672,
n33673, n33674, n33675, n33676, n33677, n33678, n33679, n33680,
n33681, n33682, n33683, n33684, n33685, n33686, n33687, n33688,
n33689, n33690, n33691, n33692, n33693, n33694, n33695, n33696,
n33697, n33698, n33699, n33700, n33701, n33702, n33703, n33704,
n33705, n33706, n33707, n33708, n33709, n33710, n33711, n33712,
n33713, n33714, n33715, n33716, n33717, n33718, n33719, n33720,
n33721, n33722, n33723, n33724, n33725, n33726, n33727, n33728,
n33729, n33730, n33731, n33732, n33733, n33734, n33735, n33736,
n33737, n33738, n33739, n33740, n33741, n33742, n33743, n33744,
n33745, n33746, n33747, n33748, n33749, n33750, n33751, n33752,
n33753, n33754, n33755, n33756, n33757, n33758, n33759, n33760,
n33761, n33762, n33763, n33764, n33765, n33766, n33767, n33768,
n33769, n33770, n33771, n33772, n33773, n33774, n33775, n33776,
n33777, n33778, n33779, n33780, n33781, n33782, n33783, n33784,
n33785, n33786, n33787, n33788, n33789, n33790, n33791, n33792,
n33793, n33794, n33795, n33796, n33797, n33798, n33799, n33800,
n33801, n33802, n33803, n33804, n33805, n33806, n33807, n33808,
n33809, n33810, n33811, n33812, n33813, n33814, n33815, n33816,
n33817, n33818, n33819, n33820, n33821, n33822, n33823, n33824,
n33825, n33826, n33827, n33828, n33829, n33830, n33831, n33832,
n33833, n33834, n33835, n33836, n33837, n33838, n33839, n33840,
n33841, n33842, n33843, n33844, n33845, n33846, n33847, n33848,
n33849, n33850, n33851, n33852, n33853, n33854, n33855, n33856,
n33857, n33858, n33859, n33860, n33861, n33862, n33863, n33864,
n33865, n33866, n33867, n33868, n33869, n33870, n33871, n33872,
n33873, n33874, n33875, n33876, n33877, n33878, n33879, n33880,
n33881, n33882, n33883, n33884, n33885, n33886, n33887, n33888,
n33889, n33890, n33891, n33892, n33893, n33894, n33895, n33896,
n33897, n33898, n33899, n33900, n33901, n33902, n33903, n33904,
n33905, n33906, n33907, n33908, n33909, n33910, n33911, n33912,
n33913, n33914, n33915, n33916, n33917, n33918, n33919, n33920,
n33921, n33922, n33923, n33924, n33925, n33926, n33927, n33928,
n33929, n33930, n33931, n33932, n33933, n33934, n33935, n33936,
n33937, n33938, n33939, n33940, n33941, n33942, n33943, n33944,
n33945, n33946, n33947, n33948, n33949, n33950, n33951, n33952,
n33953, n33954, n33955, n33956, n33957, n33958, n33959, n33960,
n33961, n33962, n33963, n33964, n33965, n33966, n33967, n33968,
n33969, n33970, n33971, n33972, n33973, n33974, n33975, n33976,
n33977, n33978, n33979, n33980, n33981, n33982, n33983, n33984,
n33985, n33986, n33987, n33988, n33989, n33990, n33991, n33992,
n33993, n33994, n33995, n33996, n33997, n33998, n33999, n34000,
n34001, n34002, n34003, n34004, n34005, n34006, n34007, n34008,
n34009, n34010, n34011, n34012, n34013, n34014, n34015, n34016,
n34017, n34018, n34019, n34020, n34021, n34022, n34023, n34024,
n34025, n34026, n34027, n34028, n34029, n34030, n34031, n34032,
n34033, n34034, n34035, n34036, n34037, n34038, n34039, n34040,
n34041, n34042, n34043, n34044, n34045, n34046, n34047, n34048,
n34049, n34050, n34051, n34052, n34053, n34054, n34055, n34056,
n34057, n34058, n34059, n34060, n34061, n34062, n34063, n34064,
n34065, n34066, n34067, n34068, n34069, n34070, n34071, n34072,
n34073, n34074, n34075, n34076, n34077, n34078, n34079, n34080,
n34081, n34082, n34083, n34084, n34085, n34086, n34087, n34088,
n34089, n34090, n34091, n34092, n34093, n34094, n34095, n34096,
n34097, n34098, n34099, n34100, n34101, n34102, n34103, n34104,
n34105, n34106, n34107, n34108, n34109, n34110, n34111, n34112,
n34113, n34114, n34115, n34116, n34117, n34118, n34119, n34120,
n34121, n34122, n34123, n34124, n34125, n34126, n34127, n34128,
n34129, n34130, n34131, n34132, n34133, n34134, n34135, n34136,
n34137, n34138, n34139, n34140, n34141, n34142, n34143, n34144,
n34145, n34146, n34147, n34148, n34149, n34150, n34151, n34152,
n34153, n34154, n34155, n34156, n34157, n34158, n34159, n34160,
n34161, n34162, n34163, n34164, n34165, n34166, n34167, n34168,
n34169, n34170, n34171, n34172, n34173, n34174, n34175, n34176,
n34177, n34178, n34179, n34180, n34181, n34182, n34183, n34184,
n34185, n34186, n34187, n34188, n34189, n34190, n34191, n34192,
n34193, n34194, n34195, n34196, n34197, n34198, n34199, n34200,
n34201, n34202, n34203, n34204, n34205, n34206, n34207, n34208,
n34209, n34210, n34211, n34212, n34213, n34214, n34215, n34216,
n34217, n34218, n34219, n34220, n34221, n34222, n34223, n34224,
n34225, n34226, n34227, n34228, n34229, n34230, n34231, n34232,
n34233, n34234, n34235, n34236, n34237, n34238, n34239, n34240,
n34241, n34242, n34243, n34244, n34245, n34246, n34247, n34248,
n34249, n34250, n34251, n34252, n34253, n34254, n34255, n34256,
n34257, n34258, n34259, n34260, n34261, n34262, n34263, n34264,
n34265, n34266, n34267, n34268, n34269, n34270, n34271, n34272,
n34273, n34274, n34275, n34276, n34277, n34278, n34279, n34280,
n34281, n34282, n34283, n34284, n34285, n34286, n34287, n34288,
n34289, n34290, n34291, n34292, n34293, n34294, n34295, n34296,
n34297, n34298, n34299, n34300, n34301, n34302, n34303, n34304,
n34305, n34306, n34307, n34308, n34309, n34310, n34311, n34312,
n34313, n34314, n34315, n34316, n34317, n34318, n34319, n34320,
n34321, n34322, n34323, n34324, n34325, n34326, n34327, n34328,
n34329, n34330, n34331, n34332, n34333, n34334, n34335, n34336,
n34337, n34338, n34339, n34340, n34341, n34342, n34343, n34344,
n34345, n34346, n34347, n34348, n34349, n34350, n34351, n34352,
n34353, n34354, n34355, n34356, n34357, n34358, n34359, n34360,
n34361, n34362, n34363, n34364, n34365, n34366, n34367, n34368,
n34369, n34370, n34371, n34372, n34373, n34374, n34375, n34376,
n34377, n34378, n34379, n34380, n34381, n34382, n34383, n34384,
n34385, n34386, n34387, n34388, n34389, n34390, n34391, n34392,
n34393, n34394, n34395, n34396, n34397, n34398, n34399, n34400,
n34401, n34402, n34403, n34404, n34405, n34406, n34407, n34408,
n34409, n34410, n34411, n34412, n34413, n34414, n34415, n34416,
n34417, n34418, n34419, n34420, n34421, n34422, n34423, n34424,
n34425, n34426, n34427, n34428, n34429, n34430, n34431, n34432,
n34433, n34434, n34435, n34436, n34437, n34438, n34439, n34440,
n34441, n34442, n34443, n34444, n34445, n34446, n34447, n34448,
n34449, n34450, n34451, n34452, n34453, n34454, n34455, n34456,
n34457, n34458, n34459, n34460, n34461, n34462, n34463, n34464,
n34465, n34466, n34467, n34468, n34469, n34470, n34471, n34472,
n34473, n34474, n34475, n34476, n34477, n34478, n34479, n34480,
n34481, n34482, n34483, n34484, n34485, n34486, n34487, n34488,
n34489, n34490, n34491, n34492, n34493, n34494, n34495, n34496,
n34497, n34498, n34499, n34500, n34501, n34502, n34503, n34504,
n34505, n34506, n34507, n34508, n34509, n34510, n34511, n34512,
n34513, n34514, n34515, n34516, n34517, n34518, n34519, n34520,
n34521, n34522, n34523, n34524, n34525, n34526, n34527, n34528,
n34529, n34530, n34531, n34532, n34533, n34534, n34535, n34536,
n34537, n34538, n34539, n34540, n34541, n34542, n34543, n34544,
n34545, n34546, n34547, n34548, n34549, n34550, n34551, n34552,
n34553, n34554, n34555, n34556, n34557, n34558, n34559, n34560,
n34561, n34562, n34563, n34564, n34565, n34566, n34567, n34568,
n34569, n34570, n34571, n34572, n34573, n34574, n34575, n34576,
n34577, n34578, n34579, n34580, n34581, n34582, n34583, n34584,
n34585, n34586, n34587, n34588, n34589, n34590, n34591, n34592,
n34593, n34594, n34595, n34596, n34597, n34598, n34599, n34600,
n34601, n34602, n34603, n34604, n34605, n34606, n34607, n34608,
n34609, n34610, n34611, n34612, n34613, n34614, n34615, n34616,
n34617, n34618, n34619, n34620, n34621, n34622, n34623, n34624,
n34625, n34626, n34627, n34628, n34629, n34630, n34631, n34632,
n34633, n34634, n34635, n34636, n34637, n34638, n34639, n34640,
n34641, n34642, n34643, n34644, n34645, n34646, n34647, n34648,
n34649, n34650, n34651, n34652, n34653, n34654, n34655, n34656,
n34657, n34658, n34659, n34660, n34661, n34662, n34663, n34664,
n34665, n34666, n34667, n34668, n34669, n34670, n34671, n34672,
n34673, n34674, n34675, n34676, n34677, n34678, n34679, n34680,
n34681, n34682, n34683, n34684, n34685, n34686, n34687, n34688,
n34689, n34690, n34691, n34692, n34693, n34694, n34695, n34696,
n34697, n34698, n34699, n34700, n34701, n34702, n34703, n34704,
n34705, n34706, n34707, n34708, n34709, n34710, n34711, n34712,
n34713, n34714, n34715, n34716, n34717, n34718, n34719, n34720,
n34721, n34722, n34723, n34724, n34725, n34726, n34727, n34728,
n34729, n34730, n34731, n34732, n34733, n34734, n34735, n34736,
n34737, n34738, n34739, n34740, n34741, n34742, n34743, n34744,
n34745, n34746, n34747, n34748, n34749, n34750, n34751, n34752,
n34753, n34754, n34755, n34756, n34757, n34758, n34759, n34760,
n34761, n34762, n34763, n34764, n34765, n34766, n34767, n34768,
n34769, n34770, n34771, n34772, n34773, n34774, n34775, n34776,
n34777, n34778, n34779, n34780, n34781, n34782, n34783, n34784,
n34785, n34786, n34787, n34788, n34789, n34790, n34791, n34792,
n34793, n34794, n34795, n34796, n34797, n34798, n34799, n34800,
n34801, n34802, n34803, n34804, n34805, n34806, n34807, n34808,
n34809, n34810, n34811, n34812, n34813, n34814, n34815, n34816,
n34817, n34818, n34819, n34820, n34821, n34822, n34823, n34824,
n34825, n34826, n34827, n34828, n34829, n34830, n34831, n34832,
n34833, n34834, n34835, n34836, n34837, n34838, n34839, n34840,
n34841, n34842, n34843, n34844, n34845, n34846, n34847, n34848,
n34849, n34850, n34851, n34852, n34853, n34854, n34855, n34856,
n34857, n34858, n34859, n34860, n34861, n34862, n34863, n34864,
n34865, n34866, n34867, n34868, n34869, n34870, n34871, n34872,
n34873, n34874, n34875, n34876, n34877, n34878, n34879, n34880,
n34881, n34882, n34883, n34884, n34885, n34886, n34887, n34888,
n34889, n34890, n34891, n34892, n34893, n34894, n34895, n34896,
n34897, n34898, n34899, n34900, n34901, n34902, n34903, n34904,
n34905, n34906, n34907, n34908, n34909, n34910, n34911, n34912,
n34913, n34914, n34915, n34916, n34917, n34918, n34919, n34920,
n34921, n34922, n34923, n34924, n34925, n34926, n34927, n34928,
n34929, n34930, n34931, n34932, n34933, n34934, n34935, n34936,
n34937, n34938, n34939, n34940, n34941, n34942, n34943, n34944,
n34945, n34946, n34947, n34948, n34949, n34950, n34951, n34952,
n34953, n34954, n34955, n34956, n34957, n34958, n34959, n34960,
n34961, n34962, n34963, n34964, n34965, n34966, n34967, n34968,
n34969, n34970, n34971, n34972, n34973, n34974, n34975, n34976,
n34977, n34978, n34979, n34980, n34981, n34982, n34983, n34984,
n34985, n34986, n34987, n34988, n34989, n34990, n34991, n34992,
n34993, n34994, n34995, n34996, n34997, n34998, n34999, n35000,
n35001, n35002, n35003, n35004, n35005, n35006, n35007, n35008,
n35009, n35010, n35011, n35012, n35013, n35014, n35015, n35016,
n35017, n35018, n35019, n35020, n35021, n35022, n35023, n35024,
n35025, n35026, n35027, n35028, n35029, n35030, n35031, n35032,
n35033, n35034, n35035, n35036, n35037, n35038, n35039, n35040,
n35041, n35042, n35043, n35044, n35045, n35046, n35047, n35048,
n35049, n35050, n35051, n35052, n35053, n35054, n35055, n35056,
n35057, n35058, n35059, n35060, n35061, n35062, n35063, n35064,
n35065, n35066, n35067, n35068, n35069, n35070, n35071, n35072,
n35073, n35074, n35075, n35076, n35077, n35078, n35079, n35080,
n35081, n35082, n35083, n35084, n35085, n35086, n35087, n35088,
n35089, n35090, n35091, n35092, n35093, n35094, n35095, n35096,
n35097, n35098, n35099, n35100, n35101, n35102, n35103, n35104,
n35105, n35106, n35107, n35108, n35109, n35110, n35111, n35112,
n35113, n35114, n35115, n35116, n35117, n35118, n35119, n35120,
n35121, n35122, n35123, n35124, n35125, n35126, n35127, n35128,
n35129, n35130, n35131, n35132, n35133, n35134, n35135, n35136,
n35137, n35138, n35139, n35140, n35141, n35142, n35143, n35144,
n35145, n35146, n35147, n35148, n35149, n35150, n35151, n35152,
n35153, n35154, n35155, n35156, n35157, n35158, n35159, n35160,
n35161, n35162, n35163, n35164, n35165, n35166, n35167, n35168,
n35169, n35170, n35171, n35172, n35173, n35174, n35175, n35176,
n35177, n35178, n35179, n35180, n35181, n35182, n35183, n35184,
n35185, n35186, n35187, n35188, n35189, n35190, n35191, n35192,
n35193, n35194, n35195, n35196, n35197, n35198, n35199, n35200,
n35201, n35202, n35203, n35204, n35205, n35206, n35207, n35208,
n35209, n35210, n35211, n35212, n35213, n35214, n35215, n35216,
n35217, n35218, n35219, n35220, n35221, n35222, n35223, n35224,
n35225, n35226, n35227, n35228, n35229, n35230, n35231, n35232,
n35233, n35234, n35235, n35236, n35237, n35238, n35239, n35240,
n35241, n35242, n35243, n35244, n35245, n35246, n35247, n35248,
n35249, n35250, n35251, n35252, n35253, n35254, n35255, n35256,
n35257, n35258, n35259, n35260, n35261, n35262, n35263, n35264,
n35265, n35266, n35267, n35268, n35269, n35270, n35271, n35272,
n35273, n35274, n35275, n35276, n35277, n35278, n35279, n35280,
n35281, n35282, n35283, n35284, n35285, n35286, n35287, n35288,
n35289, n35290, n35291, n35292, n35293, n35294, n35295, n35296,
n35297, n35298, n35299, n35300, n35301, n35302, n35303, n35304,
n35305, n35306, n35307, n35308, n35309, n35310, n35311, n35312,
n35313, n35314, n35315, n35316, n35317, n35318, n35319, n35320,
n35321, n35322, n35323, n35324, n35325, n35326, n35327, n35328,
n35329, n35330, n35331, n35332, n35333, n35334, n35335, n35336,
n35337, n35338, n35339, n35340, n35341, n35342, n35343, n35344,
n35345, n35346, n35347, n35348, n35349, n35350, n35351, n35352,
n35353, n35354, n35355, n35356, n35357, n35358, n35359, n35360,
n35361, n35362, n35363, n35364, n35365, n35366, n35367, n35368,
n35369, n35370, n35371, n35372, n35373, n35374, n35375, n35376,
n35377, n35378, n35379, n35380, n35381, n35382, n35383, n35384,
n35385, n35386, n35387, n35388, n35389, n35390, n35391, n35392,
n35393, n35394, n35395, n35396, n35397, n35398, n35399, n35400,
n35401, n35402, n35403, n35404, n35405, n35406, n35407, n35408,
n35409, n35410, n35411, n35412, n35413, n35414, n35415, n35416,
n35417, n35418, n35419, n35420, n35421, n35422, n35423, n35424,
n35425, n35426, n35427, n35428, n35429, n35430, n35431, n35432,
n35433, n35434, n35435, n35436, n35437, n35438, n35439, n35440,
n35441, n35442, n35443, n35444, n35445, n35446, n35447, n35448,
n35449, n35450, n35451, n35452, n35453, n35454, n35455, n35456,
n35457, n35458, n35459, n35460, n35461, n35462, n35463, n35464,
n35465, n35466, n35467, n35468, n35469, n35470, n35471, n35472,
n35473, n35474, n35475, n35476, n35477, n35478, n35479, n35480,
n35481, n35482, n35483, n35484, n35485, n35486, n35487, n35488,
n35489, n35490, n35491, n35492, n35493, n35494, n35495, n35496,
n35497, n35498, n35499, n35500, n35501, n35502, n35503, n35504,
n35505, n35506, n35507, n35508, n35509, n35510, n35511, n35512,
n35513, n35514, n35515, n35516, n35517, n35518, n35519, n35520,
n35521, n35522, n35523, n35524, n35525, n35526, n35527, n35528,
n35529, n35530, n35531, n35532, n35533, n35534, n35535, n35536,
n35537, n35538, n35539, n35540, n35541, n35542, n35543, n35544,
n35545, n35546, n35547, n35548, n35549, n35550, n35551, n35552,
n35553, n35554, n35555, n35556, n35557, n35558, n35559, n35560,
n35561, n35562, n35563, n35564, n35565, n35566, n35567, n35568,
n35569, n35570, n35571, n35572, n35573, n35574, n35575, n35576,
n35577, n35578, n35579, n35580, n35581, n35582, n35583, n35584,
n35585, n35586, n35587, n35588, n35589, n35590, n35591, n35592,
n35593, n35594, n35595, n35596, n35597, n35598, n35599, n35600,
n35601, n35602, n35603, n35604, n35605, n35606, n35607, n35608,
n35609, n35610, n35611, n35612, n35613, n35614, n35615, n35616,
n35617, n35618, n35619, n35620, n35621, n35622, n35623, n35624,
n35625, n35626, n35627, n35628, n35629, n35630, n35631, n35632,
n35633, n35634, n35635, n35636, n35637, n35638, n35639, n35640,
n35641, n35642, n35643, n35644, n35645, n35646, n35647, n35648,
n35649, n35650, n35651, n35652, n35653, n35654, n35655, n35656,
n35657, n35658, n35659, n35660, n35661, n35662, n35663, n35664,
n35665, n35666, n35667, n35668, n35669, n35670, n35671, n35672,
n35673, n35674, n35675, n35676, n35677, n35678, n35679, n35680,
n35681, n35682, n35683, n35684, n35685, n35686, n35687, n35688,
n35689, n35690, n35691, n35692, n35693, n35694, n35695, n35696,
n35697, n35698, n35699, n35700, n35701, n35702, n35703, n35704,
n35705, n35706, n35707, n35708, n35709, n35710, n35711, n35712,
n35713, n35714, n35715, n35716, n35717, n35718, n35719, n35720,
n35721, n35722, n35723, n35724, n35725, n35726, n35727, n35728,
n35729, n35730, n35731, n35732, n35733, n35734, n35735, n35736,
n35737, n35738, n35739, n35740, n35741, n35742, n35743, n35744,
n35745, n35746, n35747, n35748, n35749, n35750, n35751, n35752,
n35753, n35754, n35755, n35756, n35757, n35758, n35759, n35760,
n35761, n35762, n35763, n35764, n35765, n35766, n35767, n35768,
n35769, n35770, n35771, n35772, n35773, n35774, n35775, n35776,
n35777, n35778, n35779, n35780, n35781, n35782, n35783, n35784,
n35785, n35786, n35787, n35788, n35789, n35790, n35791, n35792,
n35793, n35794, n35795, n35796, n35797, n35798, n35799, n35800,
n35801, n35802, n35803, n35804, n35805, n35806, n35807, n35808,
n35809, n35810, n35811, n35812, n35813, n35814, n35815, n35816,
n35817, n35818, n35819, n35820, n35821, n35822, n35823, n35824,
n35825, n35826, n35827, n35828, n35829, n35830, n35831, n35832,
n35833, n35834, n35835, n35836, n35837, n35838, n35839, n35840,
n35841, n35842, n35843, n35844, n35845, n35846, n35847, n35848,
n35849, n35850, n35851, n35852, n35853, n35854, n35855, n35856,
n35857, n35858, n35859, n35860, n35861, n35862, n35863, n35864,
n35865, n35866, n35867, n35868, n35869, n35870, n35871, n35872,
n35873, n35874, n35875, n35876, n35877, n35878, n35879, n35880,
n35881, n35882, n35883, n35884, n35885, n35886, n35887, n35888,
n35889, n35890, n35891, n35892, n35893, n35894, n35895, n35896,
n35897, n35898, n35899, n35900, n35901, n35902, n35903, n35904,
n35905, n35906, n35907, n35908, n35909, n35910, n35911, n35912,
n35913, n35914, n35915, n35916, n35917, n35918, n35919, n35920,
n35921, n35922, n35923, n35924, n35925, n35926, n35927, n35928,
n35929, n35930, n35931, n35932, n35933, n35934, n35935, n35936,
n35937, n35938, n35939, n35940, n35941, n35942, n35943, n35944,
n35945, n35946, n35947, n35948, n35949, n35950, n35951, n35952,
n35953, n35954, n35955, n35956, n35957, n35958, n35959, n35960,
n35961, n35962, n35963, n35964, n35965, n35966, n35967, n35968,
n35969, n35970, n35971, n35972, n35973, n35974, n35975, n35976,
n35977, n35978, n35979, n35980, n35981, n35982, n35983, n35984,
n35985, n35986, n35987, n35988, n35989, n35990, n35991, n35992,
n35993, n35994, n35995, n35996, n35997, n35998, n35999, n36000,
n36001, n36002, n36003, n36004, n36005, n36006, n36007, n36008,
n36009, n36010, n36011, n36012, n36013, n36014, n36015, n36016,
n36017, n36018, n36019, n36020, n36021, n36022, n36023, n36024,
n36025, n36026, n36027, n36028, n36029, n36030, n36031, n36032,
n36033, n36034, n36035, n36036, n36037, n36038, n36039, n36040,
n36041, n36042, n36043, n36044, n36045, n36046, n36047, n36048,
n36049, n36050, n36051, n36052, n36053, n36054, n36055, n36056,
n36057, n36058, n36059, n36060, n36061, n36062, n36063, n36064,
n36065, n36066, n36067, n36068, n36069, n36070, n36071, n36072,
n36073, n36074, n36075, n36076, n36077, n36078, n36079, n36080,
n36081, n36082, n36083, n36084, n36085, n36086, n36087, n36088,
n36089, n36090, n36091, n36092, n36093, n36094, n36095, n36096,
n36097, n36098, n36099, n36100, n36101, n36102, n36103, n36104,
n36105, n36106, n36107, n36108, n36109, n36110, n36111, n36112,
n36113, n36114, n36115, n36116, n36117, n36118, n36119, n36120,
n36121, n36122, n36123, n36124, n36125, n36126, n36127, n36128,
n36129, n36130, n36131, n36132, n36133, n36134, n36135, n36136,
n36137, n36138, n36139, n36140, n36141, n36142, n36143, n36144,
n36145, n36146, n36147, n36148, n36149, n36150, n36151, n36152,
n36153, n36154, n36155, n36156, n36157, n36158, n36159, n36160,
n36161, n36162, n36163, n36164, n36165, n36166, n36167, n36168,
n36169, n36170, n36171, n36172, n36173, n36174, n36175, n36176,
n36177, n36178, n36179, n36180, n36181, n36182, n36183, n36184,
n36185, n36186, n36187, n36188, n36189, n36190, n36191, n36192,
n36193, n36194, n36195, n36196, n36197, n36198, n36199, n36200,
n36201, n36202, n36203, n36204, n36205, n36206, n36207, n36208,
n36209, n36210, n36211, n36212, n36213, n36214, n36215, n36216,
n36217, n36218, n36219, n36220, n36221, n36222, n36223, n36224,
n36225, n36226, n36227, n36228, n36229, n36230, n36231, n36232,
n36233, n36234, n36235, n36236, n36237, n36238, n36239, n36240,
n36241, n36242, n36243, n36244, n36245, n36246, n36247, n36248,
n36249, n36250, n36251, n36252, n36253, n36254, n36255, n36256,
n36257, n36258, n36259, n36260, n36261, n36262, n36263, n36264,
n36265, n36266, n36267, n36268, n36269, n36270, n36271, n36272,
n36273, n36274, n36275, n36276, n36277, n36278, n36279, n36280,
n36281, n36282, n36283, n36284, n36285, n36286, n36287, n36288,
n36289, n36290, n36291, n36292, n36293, n36294, n36295, n36296,
n36297, n36298, n36299, n36300, n36301, n36302, n36303, n36304,
n36305, n36306, n36307, n36308, n36309, n36310, n36311, n36312,
n36313, n36314, n36315, n36316, n36317, n36318, n36319, n36320,
n36321, n36322, n36323, n36324, n36325, n36326, n36327, n36328,
n36329, n36330, n36331, n36332, n36333, n36334, n36335, n36336,
n36337, n36338, n36339, n36340, n36341, n36342, n36343, n36344,
n36345, n36346, n36347, n36348, n36349, n36350, n36351, n36352,
n36353, n36354, n36355, n36356, n36357, n36358, n36359, n36360,
n36361, n36362, n36363, n36364, n36365, n36366, n36367, n36368,
n36369, n36370, n36371, n36372, n36373, n36374, n36375, n36376,
n36377, n36378, n36379, n36380, n36381, n36382, n36383, n36384,
n36385, n36386, n36387, n36388, n36389, n36390, n36391, n36392,
n36393, n36394, n36395, n36396, n36397, n36398, n36399, n36400,
n36401, n36402, n36403, n36404, n36405, n36406, n36407, n36408,
n36409, n36410, n36411, n36412, n36413, n36414, n36415, n36416,
n36417, n36418, n36419, n36420, n36421, n36422, n36423, n36424,
n36425, n36426, n36427, n36428, n36429, n36430, n36431, n36432,
n36433, n36434, n36435, n36436, n36437, n36438, n36439, n36440,
n36441, n36442, n36443, n36444, n36445, n36446, n36447, n36448,
n36449, n36450, n36451, n36452, n36453, n36454, n36455, n36456,
n36457, n36458, n36459, n36460, n36461, n36462, n36463, n36464,
n36465, n36466, n36467, n36468, n36469, n36470, n36471, n36472,
n36473, n36474, n36475, n36476, n36477, n36478, n36479, n36480,
n36481, n36482, n36483, n36484, n36485, n36486, n36487, n36488,
n36489, n36490, n36491, n36492, n36493, n36494, n36495, n36496,
n36497, n36498, n36499, n36500, n36501, n36502, n36503, n36504,
n36505, n36506, n36507, n36508, n36509, n36510, n36511, n36512,
n36513, n36514, n36515, n36516, n36517, n36518, n36519, n36520,
n36521, n36522, n36523, n36524, n36525, n36526, n36527, n36528,
n36529, n36530, n36531, n36532, n36533, n36534, n36535, n36536,
n36537, n36538, n36539, n36540, n36541, n36542, n36543, n36544,
n36545, n36546, n36547, n36548, n36549, n36550, n36551, n36552,
n36553, n36554, n36555, n36556, n36557, n36558, n36559, n36560,
n36561, n36562, n36563, n36564, n36565, n36566, n36567, n36568,
n36569, n36570, n36571, n36572, n36573, n36574, n36575, n36576,
n36577, n36578, n36579, n36580, n36581, n36582, n36583, n36584,
n36585, n36586, n36587, n36588, n36589, n36590, n36591, n36592,
n36593, n36594, n36595, n36596, n36597, n36598, n36599, n36600,
n36601, n36602, n36603, n36604, n36605, n36606, n36607, n36608,
n36609, n36610, n36611, n36612, n36613, n36614, n36615, n36616,
n36617, n36618, n36619, n36620, n36621, n36622, n36623, n36624,
n36625, n36626, n36627, n36628, n36629, n36630, n36631, n36632,
n36633, n36634, n36635, n36636, n36637, n36638, n36639, n36640,
n36641, n36642, n36643, n36644, n36645, n36646, n36647, n36648,
n36649, n36650, n36651, n36652, n36653, n36654, n36655, n36656,
n36657, n36658, n36659, n36660, n36661, n36662, n36663, n36664,
n36665, n36666, n36667, n36668, n36669, n36670, n36671, n36672,
n36673, n36674, n36675, n36676, n36677, n36678, n36679, n36680,
n36681, n36682, n36683, n36684, n36685, n36686, n36687, n36688,
n36689, n36690, n36691, n36692, n36693, n36694, n36695, n36696,
n36697, n36698, n36699, n36700, n36701, n36702, n36703, n36704,
n36705, n36706, n36707, n36708, n36709, n36710, n36711, n36712,
n36713, n36714, n36715, n36716, n36717, n36718, n36719, n36720,
n36721, n36722, n36723, n36724, n36725, n36726, n36727, n36728,
n36729, n36730, n36731, n36732, n36733, n36734, n36735, n36736,
n36737, n36738, n36739, n36740, n36741, n36742, n36743, n36744,
n36745, n36746, n36747, n36748, n36749, n36750, n36751, n36752,
n36753, n36754, n36755, n36756, n36757, n36758, n36759, n36760,
n36761, n36762, n36763, n36764, n36765, n36766, n36767, n36768,
n36769, n36770, n36771, n36772, n36773, n36774, n36775, n36776,
n36777, n36778, n36779, n36780, n36781, n36782, n36783, n36784,
n36785, n36786, n36787, n36788, n36789, n36790, n36791, n36792,
n36793, n36794, n36795, n36796, n36797, n36798, n36799, n36800,
n36801, n36802, n36803, n36804, n36805, n36806, n36807, n36808,
n36809, n36810, n36811, n36812, n36813, n36814, n36815, n36816,
n36817, n36818, n36819, n36820, n36821, n36822, n36823, n36824,
n36825, n36826, n36827, n36828, n36829, n36830, n36831, n36832,
n36833, n36834, n36835, n36836, n36837, n36838, n36839, n36840,
n36841, n36842, n36843, n36844, n36845, n36846, n36847, n36848,
n36849, n36850, n36851, n36852, n36853, n36854, n36855, n36856,
n36857, n36858, n36859, n36860, n36861, n36862, n36863, n36864,
n36865, n36866, n36867, n36868, n36869, n36870, n36871, n36872,
n36873, n36874, n36875, n36876, n36877, n36878, n36879, n36880,
n36881, n36882, n36883, n36884, n36885, n36886, n36887, n36888,
n36889, n36890, n36891, n36892, n36893, n36894, n36895, n36896,
n36897, n36898, n36899, n36900, n36901, n36902, n36903, n36904,
n36905, n36906, n36907, n36908, n36909, n36910, n36911, n36912,
n36913, n36914, n36915, n36916, n36917, n36918, n36919, n36920,
n36921, n36922, n36923, n36924, n36925, n36926, n36927, n36928,
n36929, n36930, n36931, n36932, n36933, n36934, n36935, n36936,
n36937, n36938, n36939, n36940, n36941, n36942, n36943, n36944,
n36945, n36946, n36947, n36948, n36949, n36950, n36951, n36952,
n36953, n36954, n36955, n36956, n36957, n36958, n36959, n36960,
n36961, n36962, n36963, n36964, n36965, n36966, n36967, n36968,
n36969, n36970, n36971, n36972, n36973, n36974, n36975, n36976,
n36977, n36978, n36979, n36980, n36981, n36982, n36983, n36984,
n36985, n36986, n36987, n36988, n36989, n36990, n36991, n36992,
n36993, n36994, n36995, n36996, n36997, n36998, n36999, n37000,
n37001, n37002, n37003, n37004, n37005, n37006, n37007, n37008,
n37009, n37010, n37011, n37012, n37013, n37014, n37015, n37016,
n37017, n37018, n37019, n37020, n37021, n37022, n37023, n37024,
n37025, n37026, n37027, n37028, n37029, n37030, n37031, n37032,
n37033, n37034, n37035, n37036, n37037, n37038, n37039, n37040,
n37041, n37042, n37043, n37044, n37045, n37046, n37047, n37048,
n37049, n37050, n37051, n37052, n37053, n37054, n37055, n37056,
n37057, n37058, n37059, n37060, n37061, n37062, n37063, n37064,
n37065, n37066, n37067, n37068, n37069, n37070, n37071, n37072,
n37073, n37074, n37075, n37076, n37077, n37078, n37079, n37080,
n37081, n37082, n37083, n37084, n37085, n37086, n37087, n37088,
n37089, n37090, n37091, n37092, n37093, n37094, n37095, n37096,
n37097, n37098, n37099, n37100, n37101, n37102, n37103, n37104,
n37105, n37106, n37107, n37108, n37109, n37110, n37111, n37112,
n37113, n37114, n37115, n37116, n37117, n37118, n37119, n37120,
n37121, n37122, n37123, n37124, n37125, n37126, n37127, n37128,
n37129, n37130, n37131, n37132, n37133, n37134, n37135, n37136,
n37137, n37138, n37139, n37140, n37141, n37142, n37143, n37144,
n37145, n37146, n37147, n37148, n37149, n37150, n37151, n37152,
n37153, n37154, n37155, n37156, n37157, n37158, n37159, n37160,
n37161, n37162, n37163, n37164, n37165, n37166, n37167, n37168,
n37169, n37170, n37171, n37172, n37173, n37174, n37175, n37176,
n37177, n37178, n37179, n37180, n37181, n37182, n37183, n37184,
n37185, n37186, n37187, n37188, n37189, n37190, n37191, n37192,
n37193, n37194, n37195, n37196, n37197, n37198, n37199, n37200,
n37201, n37202, n37203, n37204, n37205, n37206, n37207, n37208,
n37209, n37210, n37211, n37212, n37213, n37214, n37215, n37216,
n37217, n37218, n37219, n37220, n37221, n37222, n37223, n37224,
n37225, n37226, n37227, n37228, n37229, n37230, n37231, n37232,
n37233, n37234, n37235, n37236, n37237, n37238, n37239, n37240,
n37241, n37242, n37243, n37244, n37245, n37246, n37247, n37248,
n37249, n37250, n37251, n37252, n37253, n37254, n37255, n37256,
n37257, n37258, n37259, n37260, n37261, n37262, n37263, n37264,
n37265, n37266, n37267, n37268, n37269, n37270, n37271, n37272,
n37273, n37274, n37275, n37276, n37277, n37278, n37279, n37280,
n37281, n37282, n37283, n37284, n37285, n37286, n37287, n37288,
n37289, n37290, n37291, n37292, n37293, n37294, n37295, n37296,
n37297, n37298, n37299, n37300, n37301, n37302, n37303, n37304,
n37305, n37306, n37307, n37308, n37309, n37310, n37311, n37312,
n37313, n37314, n37315, n37316, n37317, n37318, n37319, n37320,
n37321, n37322, n37323, n37324, n37325, n37326, n37327, n37328,
n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336,
n37337, n37338, n37339, n37340, n37341, n37342, n37343, n37344,
n37345, n37346, n37347, n37348, n37349, n37350, n37351, n37352,
n37353, n37354, n37355, n37356, n37357, n37358, n37359, n37360,
n37361, n37362, n37363, n37364, n37365, n37366, n37367, n37368,
n37369, n37370, n37371, n37372, n37373, n37374, n37375, n37376,
n37377, n37378, n37379, n37380, n37381, n37382, n37383, n37384,
n37385, n37386, n37387, n37388, n37389, n37390, n37391, n37392,
n37393, n37394, n37395, n37396, n37397, n37398, n37399, n37400,
n37401, n37402, n37403, n37404, n37405, n37406, n37407, n37408,
n37409, n37410, n37411, n37412, n37413, n37414, n37415, n37416,
n37417, n37418, n37419, n37420, n37421, n37422, n37423, n37424,
n37425, n37426, n37427, n37428, n37429, n37430, n37431, n37432,
n37433, n37434, n37435, n37436, n37437, n37438, n37439, n37440,
n37441, n37442, n37443, n37444, n37445, n37446, n37447, n37448,
n37449, n37450, n37451, n37452, n37453, n37454, n37455, n37456,
n37457, n37458, n37459, n37460, n37461, n37462, n37463, n37464,
n37465, n37466, n37467, n37468, n37469, n37470, n37471, n37472,
n37473, n37474, n37475, n37476, n37477, n37478, n37479, n37480,
n37481, n37482, n37483, n37484, n37485, n37486, n37487, n37488,
n37489, n37490, n37491, n37492, n37493, n37494, n37495, n37496,
n37497, n37498, n37499, n37500, n37501, n37502, n37503, n37504,
n37505, n37506, n37507, n37508, n37509, n37510, n37511, n37512,
n37513, n37514, n37515, n37516, n37517, n37518, n37519, n37520,
n37521, n37522, n37523, n37524, n37525, n37526, n37527, n37528,
n37529, n37530, n37531, n37532, n37533, n37534, n37535, n37536,
n37537, n37538, n37539, n37540, n37541, n37542, n37543, n37544,
n37545, n37546, n37547, n37548, n37549, n37550, n37551, n37552,
n37553, n37554, n37555, n37556, n37557, n37558, n37559, n37560,
n37561, n37562, n37563, n37564, n37565, n37566, n37567, n37568,
n37569, n37570, n37571, n37572, n37573, n37574, n37575, n37576,
n37577, n37578, n37579, n37580, n37581, n37582, n37583, n37584,
n37585, n37586, n37587, n37588, n37589, n37590, n37591, n37592,
n37593, n37594, n37595, n37596, n37597, n37598, n37599, n37600,
n37601, n37602, n37603, n37604, n37605, n37606, n37607, n37608,
n37609, n37610, n37611, n37612, n37613, n37614, n37615, n37616,
n37617, n37618, n37619, n37620, n37621, n37622, n37623, n37624,
n37625, n37626, n37627, n37628, n37629, n37630, n37631, n37632,
n37633, n37634, n37635, n37636, n37637, n37638, n37639, n37640,
n37641, n37642, n37643, n37644, n37645, n37646, n37647, n37648,
n37649, n37650, n37651, n37652, n37653, n37654, n37655, n37656,
n37657, n37658, n37659, n37660, n37661, n37662, n37663, n37664,
n37665, n37666, n37667, n37668, n37669, n37670, n37671, n37672,
n37673, n37674, n37675, n37676, n37677, n37678, n37679, n37680,
n37681, n37682, n37683, n37684, n37685, n37686, n37687, n37688,
n37689, n37690, n37691, n37692, n37693, n37694, n37695, n37696,
n37697, n37698, n37699, n37700, n37701, n37702, n37703, n37704,
n37705, n37706, n37707, n37708, n37709, n37710, n37711, n37712,
n37713, n37714, n37715, n37716, n37717, n37718, n37719, n37720,
n37721, n37722, n37723, n37724, n37725, n37726, n37727, n37728,
n37729, n37730, n37731, n37732, n37733, n37734, n37735, n37736,
n37737, n37738, n37739, n37740, n37741, n37742, n37743, n37744,
n37745, n37746, n37747, n37748, n37749, n37750, n37751, n37752,
n37753, n37754, n37755, n37756, n37757, n37758, n37759, n37760,
n37761, n37762, n37763, n37764, n37765, n37766, n37767, n37768,
n37769, n37770, n37771, n37772, n37773, n37774, n37775, n37776,
n37777, n37778, n37779, n37780, n37781, n37782, n37783, n37784,
n37785, n37786, n37787, n37788, n37789, n37790, n37791, n37792,
n37793, n37794, n37795, n37796, n37797, n37798, n37799, n37800,
n37801, n37802, n37803, n37804, n37805, n37806, n37807, n37808,
n37809, n37810, n37811, n37812, n37813, n37814, n37815, n37816,
n37817, n37818, n37819, n37820, n37821, n37822, n37823, n37824,
n37825, n37826, n37827, n37828, n37829, n37830, n37831, n37832,
n37833, n37834, n37835, n37836, n37837, n37838, n37839, n37840,
n37841, n37842, n37843, n37844, n37845, n37846, n37847, n37848,
n37849, n37850, n37851, n37852, n37853, n37854, n37855, n37856,
n37857, n37858, n37859, n37860, n37861, n37862, n37863, n37864,
n37865, n37866, n37867, n37868, n37869, n37870, n37871, n37872,
n37873, n37874, n37875, n37876, n37877, n37878, n37879, n37880,
n37881, n37882, n37883, n37884, n37885, n37886, n37887, n37888,
n37889, n37890, n37891, n37892, n37893, n37894, n37895, n37896,
n37897, n37898, n37899, n37900, n37901, n37902, n37903, n37904,
n37905, n37906, n37907, n37908, n37909, n37910, n37911, n37912,
n37913, n37914, n37915, n37916, n37917, n37918, n37919, n37920,
n37921, n37922, n37923, n37924, n37925, n37926, n37927, n37928,
n37929, n37930, n37931, n37932, n37933, n37934, n37935, n37936,
n37937, n37938, n37939, n37940, n37941, n37942, n37943, n37944,
n37945, n37946, n37947, n37948, n37949, n37950, n37951, n37952,
n37953, n37954, n37955, n37956, n37957, n37958, n37959, n37960,
n37961, n37962, n37963, n37964, n37965, n37966, n37967, n37968,
n37969, n37970, n37971, n37972, n37973, n37974, n37975, n37976,
n37977, n37978, n37979, n37980, n37981, n37982, n37983, n37984,
n37985, n37986, n37987, n37988, n37989, n37990, n37991, n37992,
n37993, n37994, n37995, n37996, n37997, n37998, n37999, n38000,
n38001, n38002, n38003, n38004, n38005, n38006, n38007, n38008,
n38009, n38010, n38011, n38012, n38013, n38014, n38015, n38016,
n38017, n38018, n38019, n38020, n38021, n38022, n38023, n38024,
n38025, n38026, n38027, n38028, n38029, n38030, n38031, n38032,
n38033, n38034, n38035, n38036, n38037, n38038, n38039, n38040,
n38041, n38042, n38043, n38044, n38045, n38046, n38047, n38048,
n38049, n38050, n38051, n38052, n38053, n38054, n38055, n38056,
n38057, n38058, n38059, n38060, n38061, n38062, n38063, n38064,
n38065, n38066, n38067, n38068, n38069, n38070, n38071, n38072,
n38073, n38074, n38075, n38076, n38077, n38078, n38079, n38080,
n38081, n38082, n38083, n38084, n38085, n38086, n38087, n38088,
n38089, n38090, n38091, n38092, n38093, n38094, n38095, n38096,
n38097, n38098, n38099, n38100, n38101, n38102, n38103, n38104,
n38105, n38106, n38107, n38108, n38109, n38110, n38111, n38112,
n38113, n38114, n38115, n38116, n38117, n38118, n38119, n38120,
n38121, n38122, n38123, n38124, n38125, n38126, n38127, n38128,
n38129, n38130, n38131, n38132, n38133, n38134, n38135, n38136,
n38137, n38138, n38139, n38140, n38141, n38142, n38143, n38144,
n38145, n38146, n38147, n38148, n38149, n38150, n38151, n38152,
n38153, n38154, n38155, n38156, n38157, n38158, n38159, n38160,
n38161, n38162, n38163, n38164, n38165, n38166, n38167, n38168,
n38169, n38170, n38171, n38172, n38173, n38174, n38175, n38176,
n38177, n38178, n38179, n38180, n38181, n38182, n38183, n38184,
n38185, n38186, n38187, n38188, n38189, n38190, n38191, n38192,
n38193, n38194, n38195, n38196, n38197, n38198, n38199, n38200,
n38201, n38202, n38203, n38204, n38205, n38206, n38207, n38208,
n38209, n38210, n38211, n38212, n38213, n38214, n38215, n38216,
n38217, n38218, n38219, n38220, n38221, n38222, n38223, n38224,
n38225, n38226, n38227, n38228, n38229, n38230, n38231, n38232,
n38233, n38234, n38235, n38236, n38237, n38238, n38239, n38240,
n38241, n38242, n38243, n38244, n38245, n38246, n38247, n38248,
n38249, n38250, n38251, n38252, n38253, n38254, n38255, n38256,
n38257, n38258, n38259, n38260, n38261, n38262, n38263, n38264,
n38265, n38266, n38267, n38268, n38269, n38270, n38271, n38272,
n38273, n38274, n38275, n38276, n38277, n38278, n38279, n38280,
n38281, n38282, n38283, n38284, n38285, n38286, n38287, n38288,
n38289, n38290, n38291, n38292, n38293, n38294, n38295, n38296,
n38297, n38298, n38299, n38300, n38301, n38302, n38303, n38304,
n38305, n38306, n38307, n38308, n38309, n38310, n38311, n38312,
n38313, n38314, n38315, n38316, n38317, n38318, n38319, n38320,
n38321, n38322, n38323, n38324, n38325, n38326, n38327, n38328,
n38329, n38330, n38331, n38332, n38333, n38334, n38335, n38336,
n38337, n38338, n38339, n38340, n38341, n38342, n38343, n38344,
n38345, n38346, n38347, n38348, n38349, n38350, n38351, n38352,
n38353, n38354, n38355, n38356, n38357, n38358, n38359, n38360,
n38361, n38362, n38363, n38364, n38365, n38366, n38367, n38368,
n38369, n38370, n38371, n38372, n38373, n38374, n38375, n38376,
n38377, n38378, n38379, n38380, n38381, n38382, n38383, n38384,
n38385, n38386, n38387, n38388, n38389, n38390, n38391, n38392,
n38393, n38394, n38395, n38396, n38397, n38398, n38399, n38400,
n38401, n38402, n38403, n38404, n38405, n38406, n38407, n38408,
n38409, n38410, n38411, n38412, n38413, n38414, n38415, n38416,
n38417, n38418, n38419, n38420, n38421, n38422, n38423, n38424,
n38425, n38426, n38427, n38428, n38429, n38430, n38431, n38432,
n38433, n38434, n38435, n38436, n38437, n38438, n38439, n38440,
n38441, n38442, n38443, n38444, n38445, n38446, n38447, n38448,
n38449, n38450, n38451, n38452, n38453, n38454, n38455, n38456,
n38457, n38458, n38459, n38460, n38461, n38462, n38463, n38464,
n38465, n38466, n38467, n38468, n38469, n38470, n38471, n38472,
n38473, n38474, n38475, n38476, n38477, n38478, n38479, n38480,
n38481, n38482, n38483, n38484, n38485, n38486, n38487, n38488,
n38489, n38490, n38491, n38492, n38493, n38494, n38495, n38496,
n38497, n38498, n38499, n38500, n38501, n38502, n38503, n38504,
n38505, n38506, n38507, n38508, n38509, n38510, n38511, n38512,
n38513, n38514, n38515, n38516, n38517, n38518, n38519, n38520,
n38521, n38522, n38523, n38524, n38525, n38526, n38527, n38528,
n38529, n38530, n38531, n38532, n38533, n38534, n38535, n38536,
n38537, n38538, n38539, n38540, n38541, n38542, n38543, n38544,
n38545, n38546, n38547, n38548, n38549, n38550, n38551, n38552,
n38553, n38554, n38555, n38556, n38557, n38558, n38559, n38560,
n38561, n38562, n38563, n38564, n38565, n38566, n38567, n38568,
n38569, n38570, n38571, n38572, n38573, n38574, n38575, n38576,
n38577, n38578, n38579, n38580, n38581, n38582, n38583, n38584,
n38585, n38586, n38587, n38588, n38589, n38590, n38591, n38592,
n38593, n38594, n38595, n38596, n38597, n38598, n38599, n38600,
n38601, n38602, n38603, n38604, n38605, n38606, n38607, n38608,
n38609, n38610, n38611, n38612, n38613, n38614, n38615, n38616,
n38617, n38618, n38619, n38620, n38621, n38622, n38623, n38624,
n38625, n38626, n38627, n38628, n38629, n38630, n38631, n38632,
n38633, n38634, n38635, n38636, n38637, n38638, n38639, n38640,
n38641, n38642, n38643, n38644, n38645, n38646, n38647, n38648,
n38649, n38650, n38651, n38652, n38653, n38654, n38655, n38656,
n38657, n38658, n38659, n38660, n38661, n38662, n38663, n38664,
n38665, n38666, n38667, n38668, n38669, n38670, n38671, n38672,
n38673, n38674, n38675, n38676, n38677, n38678, n38679, n38680,
n38681, n38682, n38683, n38684, n38685, n38686, n38687, n38688,
n38689, n38690, n38691, n38692, n38693, n38694, n38695, n38696,
n38697, n38698, n38699, n38700, n38701, n38702, n38703, n38704,
n38705, n38706, n38707, n38708, n38709, n38710, n38711, n38712,
n38713, n38714, n38715, n38716, n38717, n38718, n38719, n38720,
n38721, n38722, n38723, n38724, n38725, n38726, n38727, n38728,
n38729, n38730, n38731, n38732, n38733, n38734, n38735, n38736,
n38737, n38738, n38739, n38740, n38741, n38742, n38743, n38744,
n38745, n38746, n38747, n38748, n38749, n38750, n38751, n38752,
n38753, n38754, n38755, n38756, n38757, n38758, n38759, n38760,
n38761, n38762, n38763, n38764, n38765, n38766, n38767, n38768,
n38769, n38770, n38771, n38772, n38773, n38774, n38775, n38776,
n38777, n38778, n38779, n38780, n38781, n38782, n38783, n38784,
n38785, n38786, n38787, n38788, n38789, n38790, n38791, n38792,
n38793, n38794, n38795, n38796, n38797, n38798, n38799, n38800,
n38801, n38802, n38803, n38804, n38805, n38806, n38807, n38808,
n38809, n38810, n38811, n38812, n38813, n38814, n38815, n38816,
n38817, n38818, n38819, n38820, n38821, n38822, n38823, n38824,
n38825, n38826, n38827, n38828, n38829, n38830, n38831, n38832,
n38833, n38834, n38835, n38836, n38837, n38838, n38839, n38840,
n38841, n38842, n38843, n38844, n38845, n38846, n38847, n38848,
n38849, n38850, n38851, n38852, n38853, n38854, n38855, n38856,
n38857, n38858, n38859, n38860, n38861, n38862, n38863, n38864,
n38865, n38866, n38867, n38868, n38869, n38870, n38871, n38872,
n38873, n38874, n38875, n38876, n38877, n38878, n38879, n38880,
n38881, n38882, n38883, n38884, n38885, n38886, n38887, n38888,
n38889, n38890, n38891, n38892, n38893, n38894, n38895, n38896,
n38897, n38898, n38899, n38900, n38901, n38902, n38903, n38904,
n38905, n38906, n38907, n38908, n38909, n38910, n38911, n38912,
n38913, n38914, n38915, n38916, n38917, n38918, n38919, n38920,
n38921, n38922, n38923, n38924, n38925, n38926, n38927, n38928,
n38929, n38930, n38931, n38932, n38933, n38934, n38935, n38936,
n38937, n38938, n38939, n38940, n38941, n38942, n38943, n38944,
n38945, n38946, n38947, n38948, n38949, n38950, n38951, n38952,
n38953, n38954, n38955, n38956, n38957, n38958, n38959, n38960,
n38961, n38962, n38963, n38964, n38965, n38966, n38967, n38968,
n38969, n38970, n38971, n38972, n38973, n38974, n38975, n38976,
n38977, n38978, n38979, n38980, n38981, n38982, n38983, n38984,
n38985, n38986, n38987, n38988, n38989, n38990, n38991, n38992,
n38993, n38994, n38995, n38996, n38997, n38998, n38999, n39000,
n39001, n39002, n39003, n39004, n39005, n39006, n39007, n39008,
n39009, n39010, n39011, n39012, n39013, n39014, n39015, n39016,
n39017, n39018, n39019, n39020, n39021, n39022, n39023, n39024,
n39025, n39026, n39027, n39028, n39029, n39030, n39031, n39032,
n39033, n39034, n39035, n39036, n39037, n39038, n39039, n39040,
n39041, n39042, n39043, n39044, n39045, n39046, n39047, n39048,
n39049, n39050, n39051, n39052, n39053, n39054, n39055, n39056,
n39057, n39058, n39059, n39060, n39061, n39062, n39063, n39064,
n39065, n39066, n39067, n39068, n39069, n39070, n39071, n39072,
n39073, n39074, n39075, n39076, n39077, n39078, n39079, n39080,
n39081, n39082, n39083, n39084, n39085, n39086, n39087, n39088,
n39089, n39090, n39091, n39092, n39093, n39094, n39095, n39096,
n39097, n39098, n39099, n39100, n39101, n39102, n39103, n39104,
n39105, n39106, n39107, n39108, n39109, n39110, n39111, n39112,
n39113, n39114, n39115, n39116, n39117, n39118, n39119, n39120,
n39121, n39122, n39123, n39124, n39125, n39126, n39127, n39128,
n39129, n39130, n39131, n39132, n39133, n39134, n39135, n39136,
n39137, n39138, n39139, n39140, n39141, n39142, n39143, n39144,
n39145, n39146, n39147, n39148, n39149, n39150, n39151, n39152,
n39153, n39154, n39155, n39156, n39157, n39158, n39159, n39160,
n39161, n39162, n39163, n39164, n39165, n39166, n39167, n39168,
n39169, n39170, n39171, n39172, n39173, n39174, n39175, n39176,
n39177, n39178, n39179, n39180, n39181, n39182, n39183, n39184,
n39185, n39186, n39187, n39188, n39189, n39190, n39191, n39192,
n39193, n39194, n39195, n39196, n39197, n39198, n39199, n39200,
n39201, n39202, n39203, n39204, n39205, n39206, n39207, n39208,
n39209, n39210, n39211, n39212, n39213, n39214, n39215, n39216,
n39217, n39218, n39219, n39220, n39221, n39222, n39223, n39224,
n39225, n39226, n39227, n39228, n39229, n39230, n39231, n39232,
n39233, n39234, n39235, n39236, n39237, n39238, n39239, n39240,
n39241, n39242, n39243, n39244, n39245, n39246, n39247, n39248,
n39249, n39250, n39251, n39252, n39253, n39254, n39255, n39256,
n39257, n39258, n39259, n39260, n39261, n39262, n39263, n39264,
n39265, n39266, n39267, n39268, n39269, n39270, n39271, n39272,
n39273, n39274, n39275, n39276, n39277, n39278, n39279, n39280,
n39281, n39282, n39283, n39284, n39285, n39286, n39287, n39288,
n39289, n39290, n39291, n39292, n39293, n39294, n39295, n39296,
n39297, n39298, n39299, n39300, n39301, n39302, n39303, n39304,
n39305, n39306, n39307, n39308, n39309, n39310, n39311, n39312,
n39313, n39314, n39315, n39316, n39317, n39318, n39319, n39320,
n39321, n39322, n39323, n39324, n39325, n39326, n39327, n39328,
n39329, n39330, n39331, n39332, n39333, n39334, n39335, n39336,
n39337, n39338, n39339, n39340, n39341, n39342, n39343, n39344,
n39345, n39346, n39347, n39348, n39349, n39350, n39351, n39352,
n39353, n39354, n39355, n39356, n39357, n39358, n39359, n39360,
n39361, n39362, n39363, n39364, n39365, n39366, n39367, n39368,
n39369, n39370, n39371, n39372, n39373, n39374, n39375, n39376,
n39377, n39378, n39379, n39380, n39381, n39382, n39383, n39384,
n39385, n39386, n39387, n39388, n39389, n39390, n39391, n39392,
n39393, n39394, n39395, n39396, n39397, n39398, n39399, n39400,
n39401, n39402, n39403, n39404, n39405, n39406, n39407, n39408,
n39409, n39410, n39411, n39412, n39413, n39414, n39415, n39416,
n39417, n39418, n39419, n39420, n39421, n39422, n39423, n39424,
n39425, n39426, n39427, n39428, n39429, n39430, n39431, n39432,
n39433, n39434, n39435, n39436, n39437, n39438, n39439, n39440,
n39441, n39442, n39443, n39444, n39445, n39446, n39447, n39448,
n39449, n39450, n39451, n39452, n39453, n39454, n39455, n39456,
n39457, n39458, n39459, n39460, n39461, n39462, n39463, n39464,
n39465, n39466, n39467, n39468, n39469, n39470, n39471, n39472,
n39473, n39474, n39475, n39476, n39477, n39478, n39479, n39480,
n39481, n39482, n39483, n39484, n39485, n39486, n39487, n39488,
n39489, n39490, n39491, n39492, n39493, n39494, n39495, n39496,
n39497, n39498, n39499, n39500, n39501, n39502, n39503, n39504,
n39505, n39506, n39507, n39508, n39509, n39510, n39511, n39512,
n39513, n39514, n39515, n39516, n39517, n39518, n39519, n39520,
n39521, n39522, n39523, n39524, n39525, n39526, n39527, n39528,
n39529, n39530, n39531, n39532, n39533, n39534, n39535, n39536,
n39537, n39538, n39539, n39540, n39541, n39542, n39543, n39544,
n39545, n39546, n39547, n39548, n39549, n39550, n39551, n39552,
n39553, n39554, n39555, n39556, n39557, n39558, n39559, n39560,
n39561, n39562, n39563, n39564, n39565, n39566, n39567, n39568,
n39569, n39570, n39571, n39572, n39573, n39574, n39575, n39576,
n39577, n39578, n39579, n39580, n39581, n39582, n39583, n39584,
n39585, n39586, n39587, n39588, n39589, n39590, n39591, n39592,
n39593, n39594, n39595, n39596, n39597, n39598, n39599, n39600,
n39601, n39602, n39603, n39604, n39605, n39606, n39607, n39608,
n39609, n39610, n39611, n39612, n39613, n39614, n39615, n39616,
n39617, n39618, n39619, n39620, n39621, n39622, n39623, n39624,
n39625, n39626, n39627, n39628, n39629, n39630, n39631, n39632,
n39633, n39634, n39635, n39636, n39637, n39638, n39639, n39640,
n39641, n39642, n39643, n39644, n39645, n39646, n39647, n39648,
n39649, n39650, n39651, n39652, n39653, n39654, n39655, n39656,
n39657, n39658, n39659, n39660, n39661, n39662, n39663, n39664,
n39665, n39666, n39667, n39668, n39669, n39670, n39671, n39672,
n39673, n39674, n39675, n39676, n39677, n39678, n39679, n39680,
n39681, n39682, n39683, n39684, n39685, n39686, n39687, n39688,
n39689, n39690, n39691, n39692, n39693, n39694, n39695, n39696,
n39697, n39698, n39699, n39700, n39701, n39702, n39703, n39704,
n39705, n39706, n39707, n39708, n39709, n39710, n39711, n39712,
n39713, n39714, n39715, n39716, n39717, n39718, n39719, n39720,
n39721, n39722, n39723, n39724, n39725, n39726, n39727, n39728,
n39729, n39730, n39731, n39732, n39733, n39734, n39735, n39736,
n39737, n39738, n39739, n39740, n39741, n39742, n39743, n39744,
n39745, n39746, n39747, n39748, n39749, n39750, n39751, n39752,
n39753, n39754, n39755, n39756, n39757, n39758, n39759, n39760,
n39761, n39762, n39763, n39764, n39765, n39766, n39767, n39768,
n39769, n39770, n39771, n39772, n39773, n39774, n39775, n39776,
n39777, n39778, n39779, n39780, n39781, n39782, n39783, n39784,
n39785, n39786, n39787, n39788, n39789, n39790, n39791, n39792,
n39793, n39794, n39795, n39796, n39797, n39798, n39799, n39800,
n39801, n39802, n39803, n39804, n39805, n39806, n39807, n39808,
n39809, n39810, n39811, n39812, n39813, n39814, n39815, n39816,
n39817, n39818, n39819, n39820, n39821, n39822, n39823, n39824,
n39825, n39826, n39827, n39828, n39829, n39830, n39831, n39832,
n39833, n39834, n39835, n39836, n39837, n39838, n39839, n39840,
n39841, n39842, n39843, n39844, n39845, n39846, n39847, n39848,
n39849, n39850, n39851, n39852, n39853, n39854, n39855, n39856,
n39857, n39858, n39859, n39860, n39861, n39862, n39863, n39864,
n39865, n39866, n39867, n39868, n39869, n39870, n39871, n39872,
n39873, n39874, n39875, n39876, n39877, n39878, n39879, n39880,
n39881, n39882, n39883, n39884, n39885, n39886, n39887, n39888,
n39889, n39890, n39891, n39892, n39893, n39894, n39895, n39896,
n39897, n39898, n39899, n39900, n39901, n39902, n39903, n39904,
n39905, n39906, n39907, n39908, n39909, n39910, n39911, n39912,
n39913, n39914, n39915, n39916, n39917, n39918, n39919, n39920,
n39921, n39922, n39923, n39924, n39925, n39926, n39927, n39928,
n39929, n39930, n39931, n39932, n39933, n39934, n39935, n39936,
n39937, n39938, n39939, n39940, n39941, n39942, n39943, n39944,
n39945, n39946, n39947, n39948, n39949, n39950, n39951, n39952,
n39953, n39954, n39955, n39956, n39957, n39958, n39959, n39960,
n39961, n39962, n39963, n39964, n39965, n39966, n39967, n39968,
n39969, n39970, n39971, n39972, n39973, n39974, n39975, n39976,
n39977, n39978, n39979, n39980, n39981, n39982, n39983, n39984,
n39985, n39986, n39987, n39988, n39989, n39990, n39991, n39992,
n39993, n39994, n39995, n39996, n39997, n39998, n39999, n40000,
n40001, n40002, n40003, n40004, n40005, n40006, n40007, n40008,
n40009, n40010, n40011, n40012, n40013, n40014, n40015, n40016,
n40017, n40018, n40019, n40020, n40021, n40022, n40023, n40024,
n40025, n40026, n40027, n40028, n40029, n40030, n40031, n40032,
n40033, n40034, n40035, n40036, n40037, n40038, n40039, n40040,
n40041, n40042, n40043, n40044, n40045, n40046, n40047, n40048,
n40049, n40050, n40051, n40052, n40053, n40054, n40055, n40056,
n40057, n40058, n40059, n40060, n40061, n40062, n40063, n40064,
n40065, n40066, n40067, n40068, n40069, n40070, n40071, n40072,
n40073, n40074, n40075, n40076, n40077, n40078, n40079, n40080,
n40081, n40082, n40083, n40084, n40085, n40086, n40087, n40088,
n40089, n40090, n40091, n40092, n40093, n40094, n40095, n40096,
n40097, n40098, n40099, n40100, n40101, n40102, n40103, n40104,
n40105, n40106, n40107, n40108, n40109, n40110, n40111, n40112,
n40113, n40114, n40115, n40116, n40117, n40118, n40119, n40120,
n40121, n40122, n40123, n40124, n40125, n40126, n40127, n40128,
n40129, n40130, n40131, n40132, n40133, n40134, n40135, n40136,
n40137, n40138, n40139, n40140, n40141, n40142, n40143, n40144,
n40145, n40146, n40147, n40148, n40149, n40150, n40151, n40152,
n40153, n40154, n40155, n40156, n40157, n40158, n40159, n40160,
n40161, n40162, n40163, n40164, n40165, n40166, n40167, n40168,
n40169, n40170, n40171, n40172, n40173, n40174, n40175, n40176,
n40177, n40178, n40179, n40180, n40181, n40182, n40183, n40184,
n40185, n40186, n40187, n40188, n40189, n40190, n40191, n40192,
n40193, n40194, n40195, n40196, n40197, n40198, n40199, n40200,
n40201, n40202, n40203, n40204, n40205, n40206, n40207, n40208,
n40209, n40210, n40211, n40212, n40213, n40214, n40215, n40216,
n40217, n40218, n40219, n40220, n40221, n40222, n40223, n40224,
n40225, n40226, n40227, n40228, n40229, n40230, n40231, n40232,
n40233, n40234, n40235, n40236, n40237, n40238, n40239, n40240,
n40241, n40242, n40243, n40244, n40245, n40246, n40247, n40248,
n40249, n40250, n40251, n40252, n40253, n40254, n40255, n40256,
n40257, n40258, n40259, n40260, n40261, n40262, n40263, n40264,
n40265, n40266, n40267, n40268, n40269, n40270, n40271, n40272,
n40273, n40274, n40275, n40276, n40277, n40278, n40279, n40280,
n40281, n40282, n40283, n40284, n40285, n40286, n40287, n40288,
n40289, n40290, n40291, n40292, n40293, n40294, n40295, n40296,
n40297, n40298, n40299, n40300, n40301, n40302, n40303, n40304,
n40305, n40306, n40307, n40308, n40309, n40310, n40311, n40312,
n40313, n40314, n40315, n40316, n40317, n40318, n40319, n40320,
n40321, n40322, n40323, n40324, n40325, n40326, n40327, n40328,
n40329, n40330, n40331, n40332, n40333, n40334, n40335, n40336,
n40337, n40338, n40339, n40340, n40341, n40342, n40343, n40344,
n40345, n40346, n40347, n40348, n40349, n40350, n40351, n40352,
n40353, n40354, n40355, n40356, n40357, n40358, n40359, n40360,
n40361, n40362, n40363, n40364, n40365, n40366, n40367, n40368,
n40369, n40370, n40371, n40372, n40373, n40374, n40375, n40376,
n40377, n40378, n40379, n40380, n40381, n40382, n40383, n40384,
n40385, n40386, n40387, n40388, n40389, n40390, n40391, n40392,
n40393, n40394, n40395, n40396, n40397, n40398, n40399, n40400,
n40401, n40402, n40403, n40404, n40405, n40406, n40407, n40408,
n40409, n40410, n40411, n40412, n40413, n40414, n40415, n40416,
n40417, n40418, n40419, n40420, n40421, n40422, n40423, n40424,
n40425, n40426, n40427, n40428, n40429, n40430, n40431, n40432,
n40433, n40434, n40435, n40436, n40437, n40438, n40439, n40440,
n40441, n40442, n40443, n40444, n40445, n40446, n40447, n40448,
n40449, n40450, n40451, n40452, n40453, n40454, n40455, n40456,
n40457, n40458, n40459, n40460, n40461, n40462, n40463, n40464,
n40465, n40466, n40467, n40468, n40469, n40470, n40471, n40472,
n40473, n40474, n40475, n40476, n40477, n40478, n40479, n40480,
n40481, n40482, n40483, n40484, n40485, n40486, n40487, n40488,
n40489, n40490, n40491, n40492, n40493, n40494, n40495, n40496,
n40497, n40498, n40499, n40500, n40501, n40502, n40503, n40504,
n40505, n40506, n40507, n40508, n40509, n40510, n40511, n40512,
n40513, n40514, n40515, n40516, n40517, n40518, n40519, n40520,
n40521, n40522, n40523, n40524, n40525, n40526, n40527, n40528,
n40529, n40530, n40531, n40532, n40533, n40534, n40535, n40536,
n40537, n40538, n40539, n40540, n40541, n40542, n40543, n40544,
n40545, n40546, n40547, n40548, n40549, n40550, n40551, n40552,
n40553, n40554, n40555, n40556, n40557, n40558, n40559, n40560,
n40561, n40562, n40563, n40564, n40565, n40566, n40567, n40568,
n40569, n40570, n40571, n40572, n40573, n40574, n40575, n40576,
n40577, n40578, n40579, n40580, n40581, n40582, n40583, n40584,
n40585, n40586, n40587, n40588, n40589, n40590, n40591, n40592,
n40593, n40594, n40595, n40596, n40597, n40598, n40599, n40600,
n40601, n40602, n40603, n40604, n40605, n40606, n40607, n40608,
n40609, n40610, n40611, n40612, n40613, n40614, n40615, n40616,
n40617, n40618, n40619, n40620, n40621, n40622, n40623, n40624,
n40625, n40626, n40627, n40628, n40629, n40630, n40631, n40632,
n40633, n40634, n40635, n40636, n40637, n40638, n40639, n40640,
n40641, n40642, n40643, n40644, n40645, n40646, n40647, n40648,
n40649, n40650, n40651, n40652, n40653, n40654, n40655, n40656,
n40657, n40658, n40659, n40660, n40661, n40662, n40663, n40664,
n40665, n40666, n40667, n40668, n40669, n40670, n40671, n40672,
n40673, n40674, n40675, n40676, n40677, n40678, n40679, n40680,
n40681, n40682, n40683, n40684, n40685, n40686, n40687, n40688,
n40689, n40690, n40691, n40692, n40693, n40694, n40695, n40696,
n40697, n40698, n40699, n40700, n40701, n40702, n40703, n40704,
n40705, n40706, n40707, n40708, n40709, n40710, n40711, n40712,
n40713, n40714, n40715, n40716, n40717, n40718, n40719, n40720,
n40721, n40722, n40723, n40724, n40725, n40726, n40727, n40728,
n40729, n40730, n40731, n40732, n40733, n40734, n40735, n40736,
n40737, n40738, n40739, n40740, n40741, n40742, n40743, n40744,
n40745, n40746, n40747, n40748, n40749, n40750, n40751, n40752,
n40753, n40754, n40755, n40756, n40757, n40758, n40759, n40760,
n40761, n40762, n40763, n40764, n40765, n40766, n40767, n40768,
n40769, n40770, n40771, n40772, n40773, n40774, n40775, n40776,
n40777, n40778, n40779, n40780, n40781, n40782, n40783, n40784,
n40785, n40786, n40787, n40788, n40789, n40790, n40791, n40792,
n40793, n40794, n40795, n40796, n40797, n40798, n40799, n40800,
n40801, n40802, n40803, n40804, n40805, n40806, n40807, n40808,
n40809, n40810, n40811, n40812, n40813, n40814, n40815, n40816,
n40817, n40818, n40819, n40820, n40821, n40822, n40823, n40824,
n40825, n40826, n40827, n40828, n40829, n40830, n40831, n40832,
n40833, n40834, n40835, n40836, n40837, n40838, n40839, n40840,
n40841, n40842, n40843, n40844, n40845, n40846, n40847, n40848,
n40849, n40850, n40851, n40852, n40853, n40854, n40855, n40856,
n40857, n40858, n40859, n40860, n40861, n40862, n40863, n40864,
n40865, n40866, n40867, n40868, n40869, n40870, n40871, n40872,
n40873, n40874, n40875, n40876, n40877, n40878, n40879, n40880,
n40881, n40882, n40883, n40884, n40885, n40886, n40887, n40888,
n40889, n40890, n40891, n40892, n40893, n40894, n40895, n40896,
n40897, n40898, n40899, n40900, n40901, n40902, n40903, n40904,
n40905, n40906, n40907, n40908, n40909, n40910, n40911, n40912,
n40913, n40914, n40915, n40916, n40917, n40918, n40919, n40920,
n40921, n40922, n40923, n40924, n40925, n40926, n40927, n40928,
n40929, n40930, n40931, n40932, n40933, n40934, n40935, n40936,
n40937, n40938, n40939, n40940, n40941, n40942, n40943, n40944,
n40945, n40946, n40947, n40948, n40949, n40950, n40951, n40952,
n40953, n40954, n40955, n40956, n40957, n40958, n40959, n40960,
n40961, n40962, n40963, n40964, n40965, n40966, n40967, n40968,
n40969, n40970, n40971, n40972, n40973, n40974, n40975, n40976,
n40977, n40978, n40979, n40980, n40981, n40982, n40983, n40984,
n40985, n40986, n40987, n40988, n40989, n40990, n40991, n40992,
n40993, n40994, n40995, n40996, n40997, n40998, n40999, n41000,
n41001, n41002, n41003, n41004, n41005, n41006, n41007, n41008,
n41009, n41010, n41011, n41012, n41013, n41014, n41015, n41016,
n41017, n41018, n41019, n41020, n41021, n41022, n41023, n41024,
n41025, n41026, n41027, n41028, n41029, n41030, n41031, n41032,
n41033, n41034, n41035, n41036, n41037, n41038, n41039, n41040,
n41041, n41042, n41043, n41044, n41045, n41046, n41047, n41048,
n41049, n41050, n41051, n41052, n41053, n41054, n41055, n41056,
n41057, n41058, n41059, n41060, n41061, n41062, n41063, n41064,
n41065, n41066, n41067, n41068, n41069, n41070, n41071, n41072,
n41073, n41074, n41075, n41076, n41077, n41078, n41079, n41080,
n41081, n41082, n41083, n41084, n41085, n41086, n41087, n41088,
n41089, n41090, n41091, n41092, n41093, n41094, n41095, n41096,
n41097, n41098, n41099, n41100, n41101, n41102, n41103, n41104,
n41105, n41106, n41107, n41108, n41109, n41110, n41111, n41112,
n41113, n41114, n41115, n41116, n41117, n41118, n41119, n41120,
n41121, n41122, n41123, n41124, n41125, n41126, n41127, n41128,
n41129, n41130, n41131, n41132, n41133, n41134, n41135, n41136,
n41137, n41138, n41139, n41140, n41141, n41142, n41143, n41144,
n41145, n41146, n41147, n41148, n41149, n41150, n41151, n41152,
n41153, n41154, n41155, n41156, n41157, n41158, n41159, n41160,
n41161, n41162, n41163, n41164, n41165, n41166, n41167, n41168,
n41169, n41170, n41171, n41172, n41173, n41174, n41175, n41176,
n41177, n41178, n41179, n41180, n41181, n41182, n41183, n41184,
n41185, n41186, n41187, n41188, n41189, n41190, n41191, n41192,
n41193, n41194, n41195, n41196, n41197, n41198, n41199, n41200,
n41201, n41202, n41203, n41204, n41205, n41206, n41207, n41208,
n41209, n41210, n41211, n41212, n41213, n41214, n41215, n41216,
n41217, n41218, n41219, n41220, n41221, n41222, n41223, n41224,
n41225, n41226, n41227, n41228, n41229, n41230, n41231, n41232,
n41233, n41234, n41235, n41236, n41237, n41238, n41239, n41240,
n41241, n41242, n41243, n41244, n41245, n41246, n41247, n41248,
n41249, n41250, n41251, n41252, n41253, n41254, n41255, n41256,
n41257, n41258, n41259, n41260, n41261, n41262, n41263, n41264,
n41265, n41266, n41267, n41268, n41269, n41270, n41271, n41272,
n41273, n41274, n41275, n41276, n41277, n41278, n41279, n41280,
n41281, n41282, n41283, n41284, n41285, n41286, n41287, n41288,
n41289, n41290, n41291, n41292, n41293, n41294, n41295, n41296,
n41297, n41298, n41299, n41300, n41301, n41302, n41303, n41304,
n41305, n41306, n41307, n41308, n41309, n41310, n41311, n41312,
n41313, n41314, n41315, n41316, n41317, n41318, n41319, n41320,
n41321, n41322, n41323, n41324, n41325, n41326, n41327, n41328,
n41329, n41330, n41331, n41332, n41333, n41334, n41335, n41336,
n41337, n41338, n41339, n41340, n41341, n41342, n41343, n41344,
n41345, n41346, n41347, n41348, n41349, n41350, n41351, n41352,
n41353, n41354, n41355, n41356, n41357, n41358, n41359, n41360,
n41361, n41362, n41363, n41364, n41365, n41366, n41367, n41368,
n41369, n41370, n41371, n41372, n41373, n41374, n41375, n41376,
n41377, n41378, n41379, n41380, n41381, n41382, n41383, n41384,
n41385, n41386, n41387, n41388, n41389, n41390, n41391, n41392,
n41393, n41394, n41395, n41396, n41397, n41398, n41399, n41400,
n41401, n41402, n41403, n41404, n41405, n41406, n41407, n41408,
n41409, n41410, n41411, n41412, n41413, n41414, n41415, n41416,
n41417, n41418, n41419, n41420, n41421, n41422, n41423, n41424,
n41425, n41426, n41427, n41428, n41429, n41430, n41431, n41432,
n41433, n41434, n41435, n41436, n41437, n41438, n41439, n41440,
n41441, n41442, n41443, n41444, n41445, n41446, n41447, n41448,
n41449, n41450, n41451, n41452, n41453, n41454, n41455, n41456,
n41457, n41458, n41459, n41460, n41461, n41462, n41463, n41464,
n41465, n41466, n41467, n41468, n41469, n41470, n41471, n41472,
n41473, n41474, n41475, n41476, n41477, n41478, n41479, n41480,
n41481, n41482, n41483, n41484, n41485, n41486, n41487, n41488,
n41489, n41490, n41491, n41492, n41493, n41494, n41495, n41496,
n41497, n41498, n41499, n41500, n41501, n41502, n41503, n41504,
n41505, n41506, n41507, n41508, n41509, n41510, n41511, n41512,
n41513, n41514, n41515, n41516, n41517, n41518, n41519, n41520,
n41521, n41522, n41523, n41524, n41525, n41526, n41527, n41528,
n41529, n41530, n41531, n41532, n41533, n41534, n41535, n41536,
n41537, n41538, n41539, n41540, n41541, n41542, n41543, n41544,
n41545, n41546, n41547, n41548, n41549, n41550, n41551, n41552,
n41553, n41554, n41555, n41556, n41557, n41558, n41559, n41560,
n41561, n41562, n41563, n41564, n41565, n41566, n41567, n41568,
n41569, n41570, n41571, n41572, n41573, n41574, n41575, n41576,
n41577, n41578, n41579, n41580, n41581, n41582, n41583, n41584,
n41585, n41586, n41587, n41588, n41589, n41590, n41591, n41592,
n41593, n41594, n41595, n41596, n41597, n41598, n41599, n41600,
n41601, n41602, n41603, n41604, n41605, n41606, n41607, n41608,
n41609, n41610, n41611, n41612, n41613, n41614, n41615, n41616,
n41617, n41618, n41619, n41620, n41621, n41622, n41623, n41624,
n41625, n41626, n41627, n41628, n41629, n41630, n41631, n41632,
n41633, n41634, n41635, n41636, n41637, n41638, n41639, n41640,
n41641, n41642, n41643, n41644, n41645, n41646, n41647, n41648,
n41649, n41650, n41651, n41652, n41653, n41654, n41655, n41656,
n41657, n41658, n41659, n41660, n41661, n41662, n41663, n41664,
n41665, n41666, n41667, n41668, n41669, n41670, n41671, n41672,
n41673, n41674, n41675, n41676, n41677, n41678, n41679, n41680,
n41681, n41682, n41683, n41684, n41685, n41686, n41687, n41688,
n41689, n41690, n41691, n41692, n41693, n41694, n41695, n41696,
n41697, n41698, n41699, n41700, n41701, n41702, n41703, n41704,
n41705, n41706, n41707, n41708, n41709, n41710, n41711, n41712,
n41713, n41714, n41715, n41716, n41717, n41718, n41719, n41720,
n41721, n41722, n41723, n41724, n41725, n41726, n41727, n41728,
n41729, n41730, n41731, n41732, n41733, n41734, n41735, n41736,
n41737, n41738, n41739, n41740, n41741, n41742, n41743, n41744,
n41745, n41746, n41747, n41748, n41749, n41750, n41751, n41752,
n41753, n41754, n41755, n41756, n41757, n41758, n41759, n41760,
n41761, n41762, n41763, n41764, n41765, n41766, n41767, n41768,
n41769, n41770, n41771, n41772, n41773, n41774, n41775, n41776,
n41777, n41778, n41779, n41780, n41781, n41782, n41783, n41784,
n41785, n41786, n41787, n41788, n41789, n41790, n41791, n41792,
n41793, n41794, n41795, n41796, n41797, n41798, n41799, n41800,
n41801, n41802, n41803, n41804, n41805, n41806, n41807, n41808,
n41809, n41810, n41811, n41812, n41813, n41814, n41815, n41816,
n41817, n41818, n41819, n41820, n41821, n41822, n41823, n41824,
n41825, n41826, n41827, n41828, n41829, n41830, n41831, n41832,
n41833, n41834, n41835, n41836, n41837, n41838, n41839, n41840,
n41841, n41842, n41843, n41844, n41845, n41846, n41847, n41848,
n41849, n41850, n41851, n41852, n41853, n41854, n41855, n41856,
n41857, n41858, n41859, n41860, n41861, n41862, n41863, n41864,
n41865, n41866, n41867, n41868, n41869, n41870, n41871, n41872,
n41873, n41874, n41875, n41876, n41877, n41878, n41879, n41880,
n41881, n41882, n41883, n41884, n41885, n41886, n41887, n41888,
n41889, n41890, n41891, n41892, n41893, n41894, n41895, n41896,
n41897, n41898, n41899, n41900, n41901, n41902, n41903, n41904,
n41905, n41906, n41907, n41908, n41909, n41910, n41911, n41912,
n41913, n41914, n41915, n41916, n41917, n41918, n41919, n41920,
n41921, n41922, n41923, n41924, n41925, n41926, n41927, n41928,
n41929, n41930, n41931, n41932, n41933, n41934, n41935, n41936,
n41937, n41938, n41939, n41940, n41941, n41942, n41943, n41944,
n41945, n41946, n41947, n41948, n41949, n41950, n41951, n41952,
n41953, n41954, n41955, n41956, n41957, n41958, n41959, n41960,
n41961, n41962, n41963, n41964, n41965, n41966, n41967, n41968,
n41969, n41970, n41971, n41972, n41973, n41974, n41975, n41976,
n41977, n41978, n41979, n41980, n41981, n41982, n41983, n41984,
n41985, n41986, n41987, n41988, n41989, n41990, n41991, n41992,
n41993, n41994, n41995, n41996, n41997, n41998, n41999, n42000,
n42001, n42002, n42003, n42004, n42005, n42006, n42007, n42008,
n42009, n42010, n42011, n42012, n42013, n42014, n42015, n42016,
n42017, n42018, n42019, n42020, n42021, n42022, n42023, n42024,
n42025, n42026, n42027, n42028, n42029, n42030, n42031, n42032,
n42033, n42034, n42035, n42036, n42037, n42038, n42039, n42040,
n42041, n42042, n42043, n42044, n42045, n42046, n42047, n42048,
n42049, n42050, n42051, n42052, n42053, n42054, n42055, n42056,
n42057, n42058, n42059, n42060, n42061, n42062, n42063, n42064,
n42065, n42066, n42067, n42068, n42069, n42070, n42071, n42072,
n42073, n42074, n42075, n42076, n42077, n42078, n42079, n42080,
n42081, n42082, n42083, n42084, n42085, n42086, n42087, n42088,
n42089, n42090, n42091, n42092, n42093, n42094, n42095, n42096,
n42097, n42098, n42099, n42100, n42101, n42102, n42103, n42104,
n42105, n42106, n42107, n42108, n42109, n42110, n42111, n42112,
n42113, n42114, n42115, n42116, n42117, n42118, n42119, n42120,
n42121, n42122, n42123, n42124, n42125, n42126, n42127, n42128,
n42129, n42130, n42131, n42132, n42133, n42134, n42135, n42136,
n42137, n42138, n42139, n42140, n42141, n42142, n42143, n42144,
n42145, n42146, n42147, n42148, n42149, n42150, n42151, n42152,
n42153, n42154, n42155, n42156, n42157, n42158, n42159, n42160,
n42161, n42162, n42163, n42164, n42165, n42166, n42167, n42168,
n42169, n42170, n42171, n42172, n42173, n42174, n42175, n42176,
n42177, n42178, n42179, n42180, n42181, n42182, n42183, n42184,
n42185, n42186, n42187, n42188, n42189, n42190, n42191, n42192,
n42193, n42194, n42195, n42196, n42197, n42198, n42199, n42200,
n42201, n42202, n42203, n42204, n42205, n42206, n42207, n42208,
n42209, n42210, n42211, n42212, n42213, n42214, n42215, n42216,
n42217, n42218, n42219, n42220, n42221, n42222, n42223, n42224,
n42225, n42226, n42227, n42228, n42229, n42230, n42231, n42232,
n42233, n42234, n42235, n42236, n42237, n42238, n42239, n42240,
n42241, n42242, n42243, n42244, n42245, n42246, n42247, n42248,
n42249, n42250, n42251, n42252, n42253, n42254, n42255, n42256,
n42257, n42258, n42259, n42260, n42261, n42262, n42263, n42264,
n42265, n42266, n42267, n42268, n42269, n42270, n42271, n42272,
n42273, n42274, n42275, n42276, n42277, n42278, n42279, n42280,
n42281, n42282, n42283, n42284, n42285, n42286, n42287, n42288,
n42289, n42290, n42291, n42292, n42293, n42294, n42295, n42296,
n42297, n42298, n42299, n42300, n42301, n42302, n42303, n42304,
n42305, n42306, n42307, n42308, n42309, n42310, n42311, n42312,
n42313, n42314, n42315, n42316, n42317, n42318, n42319, n42320,
n42321, n42322, n42323, n42324, n42325, n42326, n42327, n42328,
n42329, n42330, n42331, n42332, n42333, n42334, n42335, n42336,
n42337, n42338, n42339, n42340, n42341, n42342, n42343, n42344,
n42345, n42346, n42347, n42348, n42349, n42350, n42351, n42352,
n42353, n42354, n42355, n42356, n42357, n42358, n42359, n42360,
n42361, n42362, n42363, n42364, n42365, n42366, n42367, n42368,
n42369, n42370, n42371, n42372, n42373, n42374, n42375, n42376,
n42377, n42378, n42379, n42380, n42381, n42382, n42383, n42384,
n42385, n42386, n42387, n42388, n42389, n42390, n42391, n42392,
n42393, n42394, n42395, n42396, n42397, n42398, n42399, n42400,
n42401, n42402, n42403, n42404, n42405, n42406, n42407, n42408,
n42409, n42410, n42411, n42412, n42413, n42414, n42415, n42416,
n42417, n42418, n42419, n42420, n42421, n42422, n42423, n42424,
n42425, n42426, n42427, n42428, n42429, n42430, n42431, n42432,
n42433, n42434, n42435, n42436, n42437, n42438, n42439, n42440,
n42441, n42442, n42443, n42444, n42445, n42446, n42447, n42448,
n42449, n42450, n42451, n42452, n42453, n42454, n42455, n42456,
n42457, n42458, n42459, n42460, n42461, n42462, n42463, n42464,
n42465, n42466, n42467, n42468, n42469, n42470, n42471, n42472,
n42473, n42474, n42475, n42476, n42477, n42478, n42479, n42480,
n42481, n42482, n42483, n42484, n42485, n42486, n42487, n42488,
n42489, n42490, n42491, n42492, n42493, n42494, n42495, n42496,
n42497, n42498, n42499, n42500, n42501, n42502, n42503, n42504,
n42505, n42506, n42507, n42508, n42509, n42510, n42511, n42512,
n42513, n42514, n42515, n42516, n42517, n42518, n42519, n42520,
n42521, n42522, n42523, n42524, n42525, n42526, n42527, n42528,
n42529, n42530, n42531, n42532, n42533, n42534, n42535, n42536,
n42537, n42538, n42539, n42540, n42541, n42542, n42543, n42544,
n42545, n42546, n42547, n42548, n42549, n42550, n42551, n42552,
n42553, n42554, n42555, n42556, n42557, n42558, n42559, n42560,
n42561, n42562, n42563, n42564, n42565, n42566, n42567, n42568,
n42569, n42570, n42571, n42572, n42573, n42574, n42575, n42576,
n42577, n42578, n42579, n42580, n42581, n42582, n42583, n42584,
n42585, n42586, n42587, n42588, n42589, n42590, n42591, n42592,
n42593, n42594, n42595, n42596, n42597, n42598, n42599, n42600,
n42601, n42602, n42603, n42604, n42605, n42606, n42607, n42608,
n42609, n42610, n42611, n42612, n42613, n42614, n42615, n42616,
n42617, n42618, n42619, n42620, n42621, n42622, n42623, n42624,
n42625, n42626, n42627, n42628, n42629, n42630, n42631, n42632,
n42633, n42634, n42635, n42636, n42637, n42638, n42639, n42640,
n42641, n42642, n42643, n42644, n42645, n42646, n42647, n42648,
n42649, n42650, n42651, n42652, n42653, n42654, n42655, n42656,
n42657, n42658, n42659, n42660, n42661, n42662, n42663, n42664,
n42665, n42666, n42667, n42668, n42669, n42670, n42671, n42672,
n42673, n42674, n42675, n42676, n42677, n42678, n42679, n42680,
n42681, n42682, n42683, n42684, n42685, n42686, n42687, n42688,
n42689, n42690, n42691, n42692, n42693, n42694, n42695, n42696,
n42697, n42698, n42699, n42700, n42701, n42702, n42703, n42704,
n42705, n42706, n42707, n42708, n42709, n42710, n42711, n42712,
n42713, n42714, n42715, n42716, n42717, n42718, n42719, n42720,
n42721, n42722, n42723, n42724, n42725, n42726, n42727, n42728,
n42729, n42730, n42731, n42732, n42733, n42734, n42735, n42736,
n42737, n42738, n42739, n42740, n42741, n42742, n42743, n42744,
n42745, n42746, n42747, n42748, n42749, n42750, n42751, n42752,
n42753, n42754, n42755, n42756, n42757, n42758, n42759, n42760,
n42761, n42762, n42763, n42764, n42765, n42766, n42767, n42768,
n42769, n42770, n42771, n42772, n42773, n42774, n42775, n42776,
n42777, n42778, n42779, n42780, n42781, n42782, n42783, n42784,
n42785, n42786, n42787, n42788, n42789, n42790, n42791, n42792,
n42793, n42794, n42795, n42796, n42797, n42798, n42799, n42800,
n42801, n42802, n42803, n42804, n42805, n42806, n42807, n42808,
n42809, n42810, n42811, n42812, n42813, n42814, n42815, n42816,
n42817, n42818, n42819, n42820, n42821, n42822, n42823, n42824,
n42825, n42826, n42827, n42828, n42829, n42830, n42831, n42832,
n42833, n42834, n42835, n42836, n42837, n42838, n42839, n42840,
n42841, n42842, n42843, n42844, n42845, n42846, n42847, n42848,
n42849, n42850, n42851, n42852, n42853, n42854, n42855, n42856,
n42857, n42858, n42859, n42860, n42861, n42862, n42863, n42864,
n42865, n42866, n42867, n42868, n42869, n42870, n42871, n42872,
n42873, n42874, n42875, n42876, n42877, n42878, n42879, n42880,
n42881, n42882, n42883, n42884, n42885, n42886, n42887, n42888,
n42889, n42890, n42891, n42892, n42893, n42894, n42895, n42896,
n42897, n42898, n42899, n42900, n42901, n42902, n42903, n42904,
n42905, n42906, n42907, n42908, n42909, n42910, n42911, n42912,
n42913, n42914, n42915, n42916, n42917, n42918, n42919, n42920,
n42921, n42922, n42923, n42924, n42925, n42926, n42927, n42928,
n42929, n42930, n42931, n42932, n42933, n42934, n42935, n42936,
n42937, n42938, n42939, n42940, n42941, n42942, n42943, n42944,
n42945, n42946, n42947, n42948, n42949, n42950, n42951, n42952,
n42953, n42954, n42955, n42956, n42957, n42958, n42959, n42960,
n42961, n42962, n42963, n42964, n42965, n42966, n42967, n42968,
n42969, n42970, n42971, n42972, n42973, n42974, n42975, n42976,
n42977, n42978, n42979, n42980, n42981, n42982, n42983, n42984,
n42985, n42986, n42987, n42988, n42989, n42990, n42991, n42992,
n42993, n42994, n42995, n42996, n42997, n42998, n42999, n43000,
n43001, n43002, n43003, n43004, n43005, n43006, n43007, n43008,
n43009, n43010, n43011, n43012, n43013, n43014, n43015, n43016,
n43017, n43018, n43019, n43020, n43021, n43022, n43023, n43024,
n43025, n43026, n43027, n43028, n43029, n43030, n43031, n43032,
n43033, n43034, n43035, n43036, n43037, n43038, n43039, n43040,
n43041, n43042, n43043, n43044, n43045, n43046, n43047, n43048,
n43049, n43050, n43051, n43052, n43053, n43054, n43055, n43056,
n43057, n43058, n43059, n43060, n43061, n43062, n43063, n43064,
n43065, n43066, n43067, n43068, n43069, n43070, n43071, n43072,
n43073, n43074, n43075, n43076, n43077, n43078, n43079, n43080,
n43081, n43082, n43083, n43084, n43085, n43086, n43087, n43088,
n43089, n43090, n43091, n43092, n43093, n43094, n43095, n43096,
n43097, n43098, n43099, n43100, n43101, n43102, n43103, n43104,
n43105, n43106, n43107, n43108, n43109, n43110, n43111, n43112,
n43113, n43114, n43115, n43116, n43117, n43118, n43119, n43120,
n43121, n43122, n43123, n43124, n43125, n43126, n43127, n43128,
n43129, n43130, n43131, n43132, n43133, n43134, n43135, n43136,
n43137, n43138, n43139, n43140, n43141, n43142, n43143, n43144,
n43145, n43146, n43147, n43148, n43149, n43150, n43151, n43152,
n43153, n43154, n43155, n43156, n43157, n43158, n43159, n43160,
n43161, n43162, n43163, n43164, n43165, n43166, n43167, n43168,
n43169, n43170, n43171, n43172, n43173, n43174, n43175, n43176,
n43177, n43178, n43179, n43180, n43181, n43182, n43183, n43184,
n43185, n43186, n43187, n43188, n43189, n43190, n43191, n43192,
n43193, n43194, n43195, n43196, n43197, n43198, n43199, n43200,
n43201, n43202, n43203, n43204, n43205, n43206, n43207, n43208,
n43209, n43210, n43211, n43212, n43213, n43214, n43215, n43216,
n43217, n43218, n43219, n43220, n43221, n43222, n43223, n43224,
n43225, n43226, n43227, n43228, n43229, n43230, n43231, n43232,
n43233, n43234, n43235, n43236, n43237, n43238, n43239, n43240,
n43241, n43242, n43243, n43244, n43245, n43246, n43247, n43248,
n43249, n43250, n43251, n43252, n43253, n43254, n43255, n43256,
n43257, n43258, n43259, n43260, n43261, n43262, n43263, n43264,
n43265, n43266, n43267, n43268, n43269, n43270, n43271, n43272,
n43273, n43274, n43275, n43276, n43277, n43278, n43279, n43280,
n43281, n43282, n43283, n43284, n43285, n43286, n43287, n43288,
n43289, n43290, n43291, n43292, n43293, n43294, n43295, n43296,
n43297, n43298, n43299, n43300, n43301, n43302, n43303, n43304,
n43305, n43306, n43307, n43308, n43309, n43310, n43311, n43312,
n43313, n43314, n43315, n43316, n43317, n43318, n43319, n43320,
n43321, n43322, n43323, n43324, n43325, n43326, n43327, n43328,
n43329, n43330, n43331, n43332, n43333, n43334, n43335, n43336,
n43337, n43338, n43339, n43340, n43341, n43342, n43343, n43344,
n43345, n43346, n43347, n43348, n43349, n43350, n43351, n43352,
n43353, n43354, n43355, n43356, n43357, n43358, n43359, n43360,
n43361, n43362, n43363, n43364, n43365, n43366, n43367, n43368,
n43369, n43370, n43371, n43372, n43373, n43374, n43375, n43376,
n43377, n43378, n43379, n43380, n43381, n43382, n43383, n43384,
n43385, n43386, n43387, n43388, n43389, n43390, n43391, n43392,
n43393, n43394, n43395, n43396, n43397, n43398, n43399, n43400,
n43401, n43402, n43403, n43404, n43405, n43406, n43407, n43408,
n43409, n43410, n43411, n43412, n43413, n43414, n43415, n43416,
n43417, n43418, n43419, n43420, n43421, n43422, n43423, n43424,
n43425, n43426, n43427, n43428, n43429, n43430, n43431, n43432,
n43433, n43434, n43435, n43436, n43437, n43438, n43439, n43440,
n43441, n43442, n43443, n43444, n43445, n43446, n43447, n43448,
n43449, n43450, n43451, n43452, n43453, n43454, n43455, n43456,
n43457, n43458, n43459, n43460, n43461, n43462, n43463, n43464,
n43465, n43466, n43467, n43468, n43469, n43470, n43471, n43472,
n43473, n43474, n43475, n43476, n43477, n43478, n43479, n43480,
n43481, n43482, n43483, n43484, n43485, n43486, n43487, n43488,
n43489, n43490, n43491, n43492, n43493, n43494, n43495, n43496,
n43497, n43498, n43499, n43500, n43501, n43502, n43503, n43504,
n43505, n43506, n43507, n43508, n43509, n43510, n43511, n43512,
n43513, n43514, n43515, n43516, n43517, n43518, n43519, n43520,
n43521, n43522, n43523, n43524, n43525, n43526, n43527, n43528,
n43529, n43530, n43531, n43532, n43533, n43534, n43535, n43536,
n43537, n43538, n43539, n43540, n43541, n43542, n43543, n43544,
n43545, n43546, n43547, n43548, n43549, n43550, n43551, n43552,
n43553, n43554, n43555, n43556, n43557, n43558, n43559, n43560,
n43561, n43562, n43563, n43564, n43565, n43566, n43567, n43568,
n43569, n43570, n43571, n43572, n43573, n43574, n43575, n43576,
n43577, n43578, n43579, n43580, n43581, n43582, n43583, n43584,
n43585, n43586, n43587, n43588, n43589, n43590, n43591, n43592,
n43593, n43594, n43595, n43596, n43597, n43598, n43599, n43600,
n43601, n43602, n43603, n43604, n43605, n43606, n43607, n43608,
n43609, n43610, n43611, n43612, n43613, n43614, n43615, n43616,
n43617, n43618, n43619, n43620, n43621, n43622, n43623, n43624,
n43625, n43626, n43627, n43628, n43629, n43630, n43631, n43632,
n43633, n43634, n43635, n43636, n43637, n43638, n43639, n43640,
n43641, n43642, n43643, n43644, n43645, n43646, n43647, n43648,
n43649, n43650, n43651, n43652, n43653, n43654, n43655, n43656,
n43657, n43658, n43659, n43660, n43661, n43662, n43663, n43664,
n43665, n43666, n43667, n43668, n43669, n43670, n43671, n43672,
n43673, n43674, n43675, n43676, n43677, n43678, n43679, n43680,
n43681, n43682, n43683, n43684, n43685, n43686, n43687, n43688,
n43689, n43690, n43691, n43692, n43693, n43694, n43695, n43696,
n43697, n43698, n43699, n43700, n43701, n43702, n43703, n43704,
n43705, n43706, n43707, n43708, n43709, n43710, n43711, n43712,
n43713, n43714, n43715, n43716, n43717, n43718, n43719, n43720,
n43721, n43722, n43723, n43724, n43725, n43726, n43727, n43728,
n43729, n43730, n43731, n43732, n43733, n43734, n43735, n43736,
n43737, n43738, n43739, n43740, n43741, n43742, n43743, n43744,
n43745, n43746, n43747, n43748, n43749, n43750, n43751, n43752,
n43753, n43754, n43755, n43756, n43757, n43758, n43759, n43760,
n43761, n43762, n43763, n43764, n43765, n43766, n43767, n43768,
n43769, n43770, n43771, n43772, n43773, n43774, n43775, n43776,
n43777, n43778, n43779, n43780, n43781, n43782, n43783, n43784,
n43785, n43786, n43787, n43788, n43789, n43790, n43791, n43792,
n43793, n43794, n43795, n43796, n43797, n43798, n43799, n43800,
n43801, n43802, n43803, n43804, n43805, n43806, n43807, n43808,
n43809, n43810, n43811, n43812, n43813, n43814, n43815, n43816,
n43817, n43818, n43819, n43820, n43821, n43822, n43823, n43824,
n43825, n43826, n43827, n43828, n43829, n43830, n43831, n43832,
n43833, n43834, n43835, n43836, n43837, n43838, n43839, n43840,
n43841, n43842, n43843, n43844, n43845, n43846, n43847, n43848,
n43849, n43850, n43851, n43852, n43853, n43854, n43855, n43856,
n43857, n43858, n43859, n43860, n43861, n43862, n43863, n43864,
n43865, n43866, n43867, n43868, n43869, n43870, n43871, n43872,
n43873, n43874, n43875, n43876, n43877, n43878, n43879, n43880,
n43881, n43882, n43883, n43884, n43885, n43886, n43887, n43888,
n43889, n43890, n43891, n43892, n43893, n43894, n43895, n43896,
n43897, n43898, n43899, n43900, n43901, n43902, n43903, n43904,
n43905, n43906, n43907, n43908, n43909, n43910, n43911, n43912,
n43913, n43914, n43915, n43916, n43917, n43918, n43919, n43920,
n43921, n43922, n43923, n43924, n43925, n43926, n43927, n43928,
n43929, n43930, n43931, n43932, n43933, n43934, n43935, n43936,
n43937, n43938, n43939, n43940, n43941, n43942, n43943, n43944,
n43945, n43946, n43947, n43948, n43949, n43950, n43951, n43952,
n43953, n43954, n43955, n43956, n43957, n43958, n43959, n43960,
n43961, n43962, n43963, n43964, n43965, n43966, n43967, n43968,
n43969, n43970, n43971, n43972, n43973, n43974, n43975, n43976,
n43977, n43978, n43979, n43980, n43981, n43982, n43983, n43984,
n43985, n43986, n43987, n43988, n43989, n43990, n43991, n43992,
n43993, n43994, n43995, n43996, n43997, n43998, n43999, n44000,
n44001, n44002, n44003, n44004, n44005, n44006, n44007, n44008,
n44009, n44010, n44011, n44012, n44013, n44014, n44015, n44016,
n44017, n44018, n44019, n44020, n44021, n44022, n44023, n44024,
n44025, n44026, n44027, n44028, n44029, n44030, n44031, n44032,
n44033, n44034, n44035, n44036, n44037, n44038, n44039, n44040,
n44041, n44042, n44043, n44044, n44045, n44046, n44047, n44048,
n44049, n44050, n44051, n44052, n44053, n44054, n44055, n44056,
n44057, n44058, n44059, n44060, n44061, n44062, n44063, n44064,
n44065, n44066, n44067, n44068, n44069, n44070, n44071, n44072,
n44073, n44074, n44075, n44076, n44077, n44078, n44079, n44080,
n44081, n44082, n44083, n44084, n44085, n44086, n44087, n44088,
n44089, n44090, n44091, n44092, n44093, n44094, n44095, n44096,
n44097, n44098, n44099, n44100, n44101, n44102, n44103, n44104,
n44105, n44106, n44107, n44108, n44109, n44110, n44111, n44112,
n44113, n44114, n44115, n44116, n44117, n44118, n44119, n44120,
n44121, n44122, n44123, n44124, n44125, n44126, n44127, n44128,
n44129, n44130, n44131, n44132, n44133, n44134, n44135, n44136,
n44137, n44138, n44139, n44140, n44141, n44142, n44143, n44144,
n44145, n44146, n44147, n44148, n44149, n44150, n44151, n44152,
n44153, n44154, n44155, n44156, n44157, n44158, n44159, n44160,
n44161, n44162, n44163, n44164, n44165, n44166, n44167, n44168,
n44169, n44170, n44171, n44172, n44173, n44174, n44175, n44176,
n44177, n44178, n44179, n44180, n44181, n44182, n44183, n44184,
n44185, n44186, n44187, n44188, n44189, n44190, n44191, n44192,
n44193, n44194, n44195, n44196, n44197, n44198, n44199, n44200,
n44201, n44202, n44203, n44204, n44205, n44206, n44207, n44208,
n44209, n44210, n44211, n44212, n44213, n44214, n44215, n44216,
n44217, n44218, n44219, n44220, n44221, n44222, n44223, n44224,
n44225, n44226, n44227, n44228, n44229, n44230, n44231, n44232,
n44233, n44234, n44235, n44236, n44237, n44238, n44239, n44240,
n44241, n44242, n44243, n44244, n44245, n44246, n44247, n44248,
n44249, n44250, n44251, n44252, n44253, n44254, n44255, n44256,
n44257, n44258, n44259, n44260, n44261, n44262, n44263, n44264,
n44265, n44266, n44267, n44268, n44269, n44270, n44271, n44272,
n44273, n44274, n44275, n44276, n44277, n44278, n44279, n44280,
n44281, n44282, n44283, n44284, n44285, n44286, n44287, n44288,
n44289, n44290, n44291, n44292, n44293, n44294, n44295, n44296,
n44297, n44298, n44299, n44300, n44301, n44302, n44303, n44304,
n44305, n44306, n44307, n44308, n44309, n44310, n44311, n44312,
n44313, n44314, n44315, n44316, n44317, n44318, n44319, n44320,
n44321, n44322, n44323, n44324, n44325, n44326, n44327, n44328,
n44329, n44330, n44331, n44332, n44333, n44334, n44335, n44336,
n44337, n44338, n44339, n44340, n44341, n44342, n44343, n44344,
n44345, n44346, n44347, n44348, n44349, n44350, n44351, n44352,
n44353, n44354, n44355, n44356, n44357, n44358, n44359, n44360,
n44361, n44362, n44363, n44364, n44365, n44366, n44367, n44368,
n44369, n44370, n44371, n44372, n44373, n44374, n44375, n44376,
n44377, n44378, n44379, n44380, n44381, n44382, n44383, n44384,
n44385, n44386, n44387, n44388, n44389, n44390, n44391, n44392,
n44393, n44394, n44395, n44396, n44397, n44398, n44399, n44400,
n44401, n44402, n44403, n44404, n44405, n44406, n44407, n44408,
n44409, n44410, n44411, n44412, n44413, n44414, n44415, n44416,
n44417, n44418, n44419, n44420, n44421, n44422, n44423, n44424,
n44425, n44426, n44427, n44428, n44429, n44430, n44431, n44432,
n44433, n44434, n44435, n44436, n44437, n44438, n44439, n44440,
n44441, n44442, n44443, n44444, n44445, n44446, n44447, n44448,
n44449, n44450, n44451, n44452, n44453, n44454, n44455, n44456,
n44457, n44458, n44459, n44460, n44461, n44462, n44463, n44464,
n44465, n44466, n44467, n44468, n44469, n44470, n44471, n44472,
n44473, n44474, n44475, n44476, n44477, n44478, n44479, n44480,
n44481, n44482, n44483, n44484, n44485, n44486, n44487, n44488,
n44489, n44490, n44491, n44492, n44493, n44494, n44495, n44496,
n44497, n44498, n44499, n44500, n44501, n44502, n44503, n44504,
n44505, n44506, n44507, n44508, n44509, n44510, n44511, n44512,
n44513, n44514, n44515, n44516, n44517, n44518, n44519, n44520,
n44521, n44522, n44523, n44524, n44525, n44526, n44527, n44528,
n44529, n44530, n44531, n44532, n44533, n44534, n44535, n44536,
n44537, n44538, n44539, n44540, n44541, n44542, n44543, n44544,
n44545, n44546, n44547, n44548, n44549, n44550, n44551, n44552,
n44553, n44554, n44555, n44556, n44557, n44558, n44559, n44560,
n44561, n44562, n44563, n44564, n44565, n44566, n44567, n44568,
n44569, n44570, n44571, n44572, n44573, n44574, n44575, n44576,
n44577, n44578, n44579, n44580, n44581, n44582, n44583, n44584,
n44585, n44586, n44587, n44588, n44589, n44590, n44591, n44592,
n44593, n44594, n44595, n44596, n44597, n44598, n44599, n44600,
n44601, n44602, n44603, n44604, n44605, n44606, n44607, n44608,
n44609, n44610, n44611, n44612, n44613, n44614, n44615, n44616,
n44617, n44618, n44619, n44620, n44621, n44622, n44623, n44624,
n44625, n44626, n44627, n44628, n44629, n44630, n44631, n44632,
n44633, n44634, n44635, n44636, n44637, n44638, n44639, n44640,
n44641, n44642, n44643, n44644, n44645, n44646, n44647, n44648,
n44649, n44650, n44651, n44652, n44653, n44654, n44655, n44656,
n44657, n44658, n44659, n44660, n44661, n44662, n44663, n44664,
n44665, n44666, n44667, n44668, n44669, n44670, n44671, n44672,
n44673, n44674, n44675, n44676, n44677, n44678, n44679, n44680,
n44681, n44682, n44683, n44684, n44685, n44686, n44687, n44688,
n44689, n44690, n44691, n44692, n44693, n44694, n44695, n44696,
n44697, n44698, n44699, n44700, n44701, n44702, n44703, n44704,
n44705, n44706, n44707, n44708, n44709, n44710, n44711, n44712,
n44713, n44714, n44715, n44716, n44717, n44718, n44719, n44720,
n44721, n44722, n44723, n44724, n44725, n44726, n44727, n44728,
n44729, n44730, n44731, n44732, n44733, n44734, n44735, n44736,
n44737, n44738, n44739, n44740, n44741, n44742, n44743, n44744,
n44745, n44746, n44747, n44748, n44749, n44750, n44751, n44752,
n44753, n44754, n44755, n44756, n44757, n44758, n44759, n44760,
n44761, n44762, n44763, n44764, n44765, n44766, n44767, n44768,
n44769, n44770, n44771, n44772, n44773, n44774, n44775, n44776,
n44777, n44778, n44779, n44780, n44781, n44782, n44783, n44784,
n44785, n44786, n44787, n44788, n44789, n44790, n44791, n44792,
n44793, n44794, n44795, n44796, n44797, n44798, n44799, n44800,
n44801, n44802, n44803, n44804, n44805, n44806, n44807, n44808,
n44809, n44810, n44811, n44812, n44813, n44814, n44815, n44816,
n44817, n44818, n44819, n44820, n44821, n44822, n44823, n44824,
n44825, n44826, n44827, n44828, n44829, n44830, n44831, n44832,
n44833, n44834, n44835, n44836, n44837, n44838, n44839, n44840,
n44841, n44842, n44843, n44844, n44845, n44846, n44847, n44848,
n44849, n44850, n44851, n44852, n44853, n44854, n44855, n44856,
n44857, n44858, n44859, n44860, n44861, n44862, n44863, n44864,
n44865, n44866, n44867, n44868, n44869, n44870, n44871, n44872,
n44873, n44874, n44875, n44876, n44877, n44878, n44879, n44880,
n44881, n44882, n44883, n44884, n44885, n44886, n44887, n44888,
n44889, n44890, n44891, n44892, n44893, n44894, n44895, n44896,
n44897, n44898, n44899, n44900, n44901, n44902, n44903, n44904,
n44905, n44906, n44907, n44908, n44909, n44910, n44911, n44912,
n44913, n44914, n44915, n44916, n44917, n44918, n44919, n44920,
n44921, n44922, n44923, n44924, n44925, n44926, n44927, n44928,
n44929, n44930, n44931, n44932, n44933, n44934, n44935, n44936,
n44937, n44938, n44939, n44940, n44941, n44942, n44943, n44944,
n44945, n44946, n44947, n44948, n44949, n44950, n44951, n44952,
n44953, n44954, n44955, n44956, n44957, n44958, n44959, n44960,
n44961, n44962, n44963, n44964, n44965, n44966, n44967, n44968,
n44969, n44970, n44971, n44972, n44973, n44974, n44975, n44976,
n44977, n44978, n44979, n44980, n44981, n44982, n44983, n44984,
n44985, n44986, n44987, n44988, n44989, n44990, n44991, n44992,
n44993, n44994, n44995, n44996, n44997, n44998, n44999, n45000,
n45001, n45002, n45003, n45004, n45005, n45006, n45007, n45008,
n45009, n45010, n45011, n45012, n45013, n45014, n45015, n45016,
n45017, n45018, n45019, n45020, n45021, n45022, n45023, n45024,
n45025, n45026, n45027, n45028, n45029, n45030, n45031, n45032,
n45033, n45034, n45035, n45036, n45037, n45038, n45039, n45040,
n45041, n45042, n45043, n45044, n45045, n45046, n45047, n45048,
n45049, n45050, n45051, n45052, n45053, n45054, n45055, n45056,
n45057, n45058, n45059, n45060, n45061, n45062, n45063, n45064,
n45065, n45066, n45067, n45068, n45069, n45070, n45071, n45072,
n45073, n45074, n45075, n45076, n45077, n45078, n45079, n45080,
n45081, n45082, n45083, n45084, n45085, n45086, n45087, n45088,
n45089, n45090, n45091, n45092, n45093, n45094, n45095, n45096,
n45097, n45098, n45099, n45100, n45101, n45102, n45103, n45104,
n45105, n45106, n45107, n45108, n45109, n45110, n45111, n45112,
n45113, n45114, n45115, n45116, n45117, n45118, n45119, n45120,
n45121, n45122, n45123, n45124, n45125, n45126, n45127, n45128,
n45129, n45130, n45131, n45132, n45133, n45134, n45135, n45136,
n45137, n45138, n45139, n45140, n45141, n45142, n45143, n45144,
n45145, n45146, n45147, n45148, n45149, n45150, n45151, n45152,
n45153, n45154, n45155, n45156, n45157, n45158, n45159, n45160,
n45161, n45162, n45163, n45164, n45165, n45166, n45167, n45168,
n45169, n45170, n45171, n45172, n45173, n45174, n45175, n45176,
n45177, n45178, n45179, n45180, n45181, n45182, n45183, n45184,
n45185, n45186, n45187, n45188, n45189, n45190, n45191, n45192,
n45193, n45194, n45195, n45196, n45197, n45198, n45199, n45200,
n45201, n45202, n45203, n45204, n45205, n45206, n45207, n45208,
n45209, n45210, n45211, n45212, n45213, n45214, n45215, n45216,
n45217, n45218, n45219, n45220, n45221, n45222, n45223, n45224,
n45225, n45226, n45227, n45228, n45229, n45230, n45231, n45232,
n45233, n45234, n45235, n45236, n45237, n45238, n45239, n45240,
n45241, n45242, n45243, n45244, n45245, n45246, n45247, n45248,
n45249, n45250, n45251, n45252, n45253, n45254, n45255, n45256,
n45257, n45258, n45259, n45260, n45261, n45262, n45263, n45264,
n45265, n45266, n45267, n45268, n45269, n45270, n45271, n45272,
n45273, n45274, n45275, n45276, n45277, n45278, n45279, n45280,
n45281, n45282, n45283, n45284, n45285, n45286, n45287, n45288,
n45289, n45290, n45291, n45292, n45293, n45294, n45295, n45296,
n45297, n45298, n45299, n45300, n45301, n45302, n45303, n45304,
n45305, n45306, n45307, n45308, n45309, n45310, n45311, n45312,
n45313, n45314, n45315, n45316, n45317, n45318, n45319, n45320,
n45321, n45322, n45323, n45324, n45325, n45326, n45327, n45328,
n45329, n45330, n45331, n45332, n45333, n45334, n45335, n45336,
n45337, n45338, n45339, n45340, n45341, n45342, n45343, n45344,
n45345, n45346, n45347, n45348, n45349, n45350, n45351, n45352,
n45353, n45354, n45355, n45356, n45357, n45358, n45359, n45360,
n45361, n45362, n45363, n45364, n45365, n45366, n45367, n45368,
n45369, n45370, n45371, n45372, n45373, n45374, n45375, n45376,
n45377, n45378, n45379, n45380, n45381, n45382, n45383, n45384,
n45385, n45386, n45387, n45388, n45389, n45390, n45391, n45392,
n45393, n45394, n45395, n45396, n45397, n45398, n45399, n45400,
n45401, n45402, n45403, n45404, n45405, n45406, n45407, n45408,
n45409, n45410, n45411, n45412, n45413, n45414, n45415, n45416,
n45417, n45418, n45419, n45420, n45421, n45422, n45423, n45424,
n45425, n45426, n45427, n45428, n45429, n45430, n45431, n45432,
n45433, n45434, n45435, n45436, n45437, n45438, n45439, n45440,
n45441, n45442, n45443, n45444, n45445, n45446, n45447, n45448,
n45449, n45450, n45451, n45452, n45453, n45454, n45455, n45456,
n45457, n45458, n45459, n45460, n45461, n45462, n45463, n45464,
n45465, n45466, n45467, n45468, n45469, n45470, n45471, n45472,
n45473, n45474, n45475, n45476, n45477, n45478, n45479, n45480,
n45481, n45482, n45483, n45484, n45485, n45486, n45487, n45488,
n45489, n45490, n45491, n45492, n45493, n45494, n45495, n45496,
n45497, n45498, n45499, n45500, n45501, n45502, n45503, n45504,
n45505, n45506, n45507, n45508, n45509, n45510, n45511, n45512,
n45513, n45514, n45515, n45516, n45517, n45518, n45519, n45520,
n45521, n45522, n45523, n45524, n45525, n45526, n45527, n45528,
n45529, n45530, n45531, n45532, n45533, n45534, n45535, n45536,
n45537, n45538, n45539, n45540, n45541, n45542, n45543, n45544,
n45545, n45546, n45547, n45548, n45549, n45550, n45551, n45552,
n45553, n45554, n45555, n45556, n45557, n45558, n45559, n45560,
n45561, n45562, n45563, n45564, n45565, n45566, n45567, n45568,
n45569, n45570, n45571, n45572, n45573, n45574, n45575, n45576,
n45577, n45578, n45579, n45580, n45581, n45582, n45583, n45584,
n45585, n45586, n45587, n45588, n45589, n45590, n45591, n45592,
n45593, n45594, n45595, n45596, n45597, n45598, n45599, n45600,
n45601, n45602, n45603, n45604, n45605, n45606, n45607, n45608,
n45609, n45610, n45611, n45612, n45613, n45614, n45615, n45616,
n45617, n45618, n45619, n45620, n45621, n45622, n45623, n45624,
n45625, n45626, n45627, n45628, n45629, n45630, n45631, n45632,
n45633, n45634, n45635, n45636, n45637, n45638, n45639, n45640,
n45641, n45642, n45643, n45644, n45645, n45646, n45647, n45648,
n45649, n45650, n45651, n45652, n45653, n45654, n45655, n45656,
n45657, n45658, n45659, n45660, n45661, n45662, n45663, n45664,
n45665, n45666, n45667, n45668, n45669, n45670, n45671, n45672,
n45673, n45674, n45675, n45676, n45677, n45678, n45679, n45680,
n45681, n45682, n45683, n45684, n45685, n45686, n45687, n45688,
n45689, n45690, n45691, n45692, n45693, n45694, n45695, n45696,
n45697, n45698, n45699, n45700, n45701, n45702, n45703, n45704,
n45705, n45706, n45707, n45708, n45709, n45710, n45711, n45712,
n45713, n45714, n45715, n45716, n45717, n45718, n45719, n45720,
n45721, n45722, n45723, n45724, n45725, n45726, n45727, n45728,
n45729, n45730, n45731, n45732, n45733, n45734, n45735, n45736,
n45737, n45738, n45739, n45740, n45741, n45742, n45743, n45744,
n45745, n45746, n45747, n45748, n45749, n45750, n45751, n45752,
n45753, n45754, n45755, n45756, n45757, n45758, n45759, n45760,
n45761, n45762, n45763, n45764, n45765, n45766, n45767, n45768,
n45769, n45770, n45771, n45772, n45773, n45774, n45775, n45776,
n45777, n45778, n45779, n45780, n45781, n45782, n45783, n45784,
n45785, n45786, n45787, n45788, n45789, n45790, n45791, n45792,
n45793, n45794, n45795, n45796, n45797, n45798, n45799, n45800,
n45801, n45802, n45803, n45804, n45805, n45806, n45807, n45808,
n45809, n45810, n45811, n45812, n45813, n45814, n45815, n45816,
n45817, n45818, n45819, n45820, n45821, n45822, n45823, n45824,
n45825, n45826, n45827, n45828, n45829, n45830, n45831, n45832,
n45833, n45834, n45835, n45836, n45837, n45838, n45839, n45840,
n45841, n45842, n45843, n45844, n45845, n45846, n45847, n45848,
n45849, n45850, n45851, n45852, n45853, n45854, n45855, n45856,
n45857, n45858, n45859, n45860, n45861, n45862, n45863, n45864,
n45865, n45866, n45867, n45868, n45869, n45870, n45871, n45872,
n45873, n45874, n45875, n45876, n45877, n45878, n45879, n45880,
n45881, n45882, n45883, n45884, n45885, n45886, n45887, n45888,
n45889, n45890, n45891, n45892, n45893, n45894, n45895, n45896,
n45897, n45898, n45899, n45900, n45901, n45902, n45903, n45904,
n45905, n45906, n45907, n45908, n45909, n45910, n45911, n45912,
n45913, n45914, n45915, n45916, n45917, n45918, n45919, n45920,
n45921, n45922, n45923, n45924, n45925, n45926, n45927, n45928,
n45929, n45930, n45931, n45932, n45933, n45934, n45935, n45936,
n45937, n45938, n45939, n45940, n45941, n45942, n45943, n45944,
n45945, n45946, n45947, n45948, n45949, n45950, n45951, n45952,
n45953, n45954, n45955, n45956, n45957, n45958, n45959, n45960,
n45961, n45962, n45963, n45964, n45965, n45966, n45967, n45968,
n45969, n45970, n45971, n45972, n45973, n45974, n45975, n45976,
n45977, n45978, n45979, n45980, n45981, n45982, n45983, n45984,
n45985, n45986, n45987, n45988, n45989, n45990, n45991, n45992,
n45993, n45994, n45995, n45996, n45997, n45998, n45999, n46000,
n46001, n46002, n46003, n46004, n46005, n46006, n46007, n46008,
n46009, n46010, n46011, n46012, n46013, n46014, n46015, n46016,
n46017, n46018, n46019, n46020, n46021, n46022, n46023, n46024,
n46025, n46026, n46027, n46028, n46029, n46030, n46031, n46032,
n46033, n46034, n46035, n46036, n46037, n46038, n46039, n46040,
n46041, n46042, n46043, n46044, n46045, n46046, n46047, n46048,
n46049, n46050, n46051, n46052, n46053, n46054, n46055, n46056,
n46057, n46058, n46059, n46060, n46061, n46062, n46063, n46064,
n46065, n46066, n46067, n46068, n46069, n46070, n46071, n46072,
n46073, n46074, n46075, n46076, n46077, n46078, n46079, n46080,
n46081, n46082, n46083, n46084, n46085, n46086, n46087, n46088,
n46089, n46090, n46091, n46092, n46093, n46094, n46095, n46096,
n46097, n46098, n46099, n46100, n46101, n46102, n46103, n46104,
n46105, n46106, n46107, n46108, n46109, n46110, n46111, n46112,
n46113, n46114, n46115, n46116, n46117, n46118, n46119, n46120,
n46121, n46122, n46123, n46124, n46125, n46126, n46127, n46128,
n46129, n46130, n46131, n46132, n46133, n46134, n46135, n46136,
n46137, n46138, n46139, n46140, n46141, n46142, n46143, n46144,
n46145, n46146, n46147, n46148, n46149, n46150, n46151, n46152,
n46153, n46154, n46155, n46156, n46157, n46158, n46159, n46160,
n46161, n46162, n46163, n46164, n46165, n46166, n46167, n46168,
n46169, n46170, n46171, n46172, n46173, n46174, n46175, n46176,
n46177, n46178, n46179, n46180, n46181, n46182, n46183, n46184,
n46185, n46186, n46187, n46188, n46189, n46190, n46191, n46192,
n46193, n46194, n46195, n46196, n46197, n46198, n46199, n46200,
n46201, n46202, n46203, n46204, n46205, n46206, n46207, n46208,
n46209, n46210, n46211, n46212, n46213, n46214, n46215, n46216,
n46217, n46218, n46219, n46220, n46221, n46222, n46223, n46224,
n46225, n46226, n46227, n46228, n46229, n46230, n46231, n46232,
n46233, n46234, n46235, n46236, n46237, n46238, n46239, n46240,
n46241, n46242, n46243, n46244, n46245, n46246, n46247, n46248,
n46249, n46250, n46251, n46252, n46253, n46254, n46255, n46256,
n46257, n46258, n46259, n46260, n46261, n46262, n46263, n46264,
n46265, n46266, n46267, n46268, n46269, n46270, n46271, n46272,
n46273, n46274, n46275, n46276, n46277, n46278, n46279, n46280,
n46281, n46282, n46283, n46284, n46285, n46286, n46287, n46288,
n46289, n46290, n46291, n46292, n46293, n46294, n46295, n46296,
n46297, n46298, n46299, n46300, n46301, n46302, n46303, n46304,
n46305, n46306, n46307, n46308, n46309, n46310, n46311, n46312,
n46313, n46314, n46315, n46316, n46317, n46318, n46319, n46320,
n46321, n46322, n46323, n46324, n46325, n46326, n46327, n46328,
n46329, n46330, n46331, n46332, n46333, n46334, n46335, n46336,
n46337, n46338, n46339, n46340, n46341, n46342, n46343, n46344,
n46345, n46346, n46347, n46348, n46349, n46350, n46351, n46352,
n46353, n46354, n46355, n46356, n46357, n46358, n46359, n46360,
n46361, n46362, n46363, n46364, n46365, n46366, n46367, n46368,
n46369, n46370, n46371, n46372, n46373, n46374, n46375, n46376,
n46377, n46378, n46379, n46380, n46381, n46382, n46383, n46384,
n46385, n46386, n46387, n46388, n46389, n46390, n46391, n46392,
n46393, n46394, n46395, n46396, n46397, n46398, n46399, n46400,
n46401, n46402, n46403, n46404, n46405, n46406, n46407, n46408,
n46409, n46410, n46411, n46412, n46413, n46414, n46415, n46416,
n46417, n46418, n46419, n46420, n46421, n46422, n46423, n46424,
n46425, n46426, n46427, n46428, n46429, n46430, n46431, n46432,
n46433, n46434, n46435, n46436, n46437, n46438, n46439, n46440,
n46441, n46442, n46443, n46444, n46445, n46446, n46447, n46448,
n46449, n46450, n46451, n46452, n46453, n46454, n46455, n46456,
n46457, n46458, n46459, n46460, n46461, n46462, n46463, n46464,
n46465, n46466, n46467, n46468, n46469, n46470, n46471, n46472,
n46473, n46474, n46475, n46476, n46477, n46478, n46479, n46480,
n46481, n46482, n46483, n46484, n46485, n46486, n46487, n46488,
n46489, n46490, n46491, n46492, n46493, n46494, n46495, n46496,
n46497, n46498, n46499, n46500, n46501, n46502, n46503, n46504,
n46505, n46506, n46507, n46508, n46509, n46510, n46511, n46512,
n46513, n46514, n46515, n46516, n46517, n46518, n46519, n46520,
n46521, n46522, n46523, n46524, n46525, n46526, n46527, n46528,
n46529, n46530, n46531, n46532, n46533, n46534, n46535, n46536,
n46537, n46538, n46539, n46540, n46541, n46542, n46543, n46544,
n46545, n46546, n46547, n46548, n46549, n46550, n46551, n46552,
n46553, n46554, n46555, n46556, n46557, n46558, n46559, n46560,
n46561, n46562, n46563, n46564, n46565, n46566, n46567, n46568,
n46569, n46570, n46571, n46572, n46573, n46574, n46575, n46576,
n46577, n46578, n46579, n46580, n46581, n46582, n46583, n46584,
n46585, n46586, n46587, n46588, n46589, n46590, n46591, n46592,
n46593, n46594, n46595, n46596, n46597, n46598, n46599, n46600,
n46601, n46602, n46603, n46604, n46605, n46606, n46607, n46608,
n46609, n46610, n46611, n46612, n46613, n46614, n46615, n46616,
n46617, n46618, n46619, n46620, n46621, n46622, n46623, n46624,
n46625, n46626, n46627, n46628, n46629, n46630, n46631, n46632,
n46633, n46634, n46635, n46636, n46637, n46638, n46639, n46640,
n46641, n46642, n46643, n46644, n46645, n46646, n46647, n46648,
n46649, n46650, n46651, n46652, n46653, n46654, n46655, n46656,
n46657, n46658, n46659, n46660, n46661, n46662, n46663, n46664,
n46665, n46666, n46667, n46668, n46669, n46670, n46671, n46672,
n46673, n46674, n46675, n46676, n46677, n46678, n46679, n46680,
n46681, n46682, n46683, n46684, n46685, n46686, n46687, n46688,
n46689, n46690, n46691, n46692, n46693, n46694, n46695, n46696,
n46697, n46698, n46699, n46700, n46701, n46702, n46703, n46704,
n46705, n46706, n46707, n46708, n46709, n46710, n46711, n46712,
n46713, n46714, n46715, n46716, n46717, n46718, n46719, n46720,
n46721, n46722, n46723, n46724, n46725, n46726, n46727, n46728,
n46729, n46730, n46731, n46732, n46733, n46734, n46735, n46736,
n46737, n46738, n46739, n46740, n46741, n46742, n46743, n46744,
n46745, n46746, n46747, n46748, n46749, n46750, n46751, n46752,
n46753, n46754, n46755, n46756, n46757, n46758, n46759, n46760,
n46761, n46762, n46763, n46764, n46765, n46766, n46767, n46768,
n46769, n46770, n46771, n46772, n46773, n46774, n46775, n46776,
n46777, n46778, n46779, n46780, n46781, n46782, n46783, n46784,
n46785, n46786, n46787, n46788, n46789, n46790, n46791, n46792,
n46793, n46794, n46795, n46796, n46797, n46798, n46799, n46800,
n46801, n46802, n46803, n46804, n46805, n46806, n46807, n46808,
n46809, n46810, n46811, n46812, n46813, n46814, n46815, n46816,
n46817, n46818, n46819, n46820, n46821, n46822, n46823, n46824,
n46825, n46826, n46827, n46828, n46829, n46830, n46831, n46832,
n46833, n46834, n46835, n46836, n46837, n46838, n46839, n46840,
n46841, n46842, n46843, n46844, n46845, n46846, n46847, n46848,
n46849, n46850, n46851, n46852, n46853, n46854, n46855, n46856,
n46857, n46858, n46859, n46860, n46861, n46862, n46863, n46864,
n46865, n46866, n46867, n46868, n46869, n46870, n46871, n46872,
n46873, n46874, n46875, n46876, n46877, n46878, n46879, n46880,
n46881, n46882, n46883, n46884, n46885, n46886, n46887, n46888,
n46889, n46890, n46891, n46892, n46893, n46894, n46895, n46896,
n46897, n46898, n46899, n46900, n46901, n46902, n46903, n46904,
n46905, n46906, n46907, n46908, n46909, n46910, n46911, n46912,
n46913, n46914, n46915, n46916, n46917, n46918, n46919, n46920,
n46921, n46922, n46923, n46924, n46925, n46926, n46927, n46928,
n46929, n46930, n46931, n46932, n46933, n46934, n46935, n46936,
n46937, n46938, n46939, n46940, n46941, n46942, n46943, n46944,
n46945, n46946, n46947, n46948, n46949, n46950, n46951, n46952,
n46953, n46954, n46955, n46956, n46957, n46958, n46959, n46960,
n46961, n46962, n46963, n46964, n46965, n46966, n46967, n46968,
n46969, n46970, n46971, n46972, n46973, n46974, n46975, n46976,
n46977, n46978, n46979, n46980, n46981, n46982, n46983, n46984,
n46985, n46986, n46987, n46988, n46989, n46990, n46991, n46992,
n46993, n46994, n46995, n46996, n46997, n46998, n46999, n47000,
n47001, n47002, n47003, n47004, n47005, n47006, n47007, n47008,
n47009, n47010, n47011, n47012, n47013, n47014, n47015, n47016,
n47017, n47018, n47019, n47020, n47021, n47022, n47023, n47024,
n47025, n47026, n47027, n47028, n47029, n47030, n47031, n47032,
n47033, n47034, n47035, n47036, n47037, n47038, n47039, n47040,
n47041, n47042, n47043, n47044, n47045, n47046, n47047, n47048,
n47049, n47050, n47051, n47052, n47053, n47054, n47055, n47056,
n47057, n47058, n47059, n47060, n47061, n47062, n47063, n47064,
n47065, n47066, n47067, n47068, n47069, n47070, n47071, n47072,
n47073, n47074, n47075, n47076, n47077, n47078, n47079, n47080,
n47081, n47082, n47083, n47084, n47085, n47086, n47087, n47088,
n47089, n47090, n47091, n47092, n47093, n47094, n47095, n47096,
n47097, n47098, n47099, n47100, n47101, n47102, n47103, n47104,
n47105, n47106, n47107, n47108, n47109, n47110, n47111, n47112,
n47113, n47114, n47115, n47116, n47117, n47118, n47119, n47120,
n47121, n47122, n47123, n47124, n47125, n47126, n47127, n47128,
n47129, n47130, n47131, n47132, n47133, n47134, n47135, n47136,
n47137, n47138, n47139, n47140, n47141, n47142, n47143, n47144,
n47145, n47146, n47147, n47148, n47149, n47150, n47151, n47152,
n47153, n47154, n47155, n47156, n47157, n47158, n47159, n47160,
n47161, n47162, n47163, n47164, n47165, n47166, n47167, n47168,
n47169, n47170, n47171, n47172, n47173, n47174, n47175, n47176,
n47177, n47178, n47179, n47180, n47181, n47182, n47183, n47184,
n47185, n47186, n47187, n47188, n47189, n47190, n47191, n47192,
n47193, n47194, n47195, n47196, n47197, n47198, n47199, n47200,
n47201, n47202, n47203, n47204, n47205, n47206, n47207, n47208,
n47209, n47210, n47211, n47212, n47213, n47214, n47215, n47216,
n47217, n47218, n47219, n47220, n47221, n47222, n47223, n47224,
n47225, n47226, n47227, n47228, n47229, n47230, n47231, n47232,
n47233, n47234, n47235, n47236, n47237, n47238, n47239, n47240,
n47241, n47242, n47243, n47244, n47245, n47246, n47247, n47248,
n47249, n47250, n47251, n47252, n47253, n47254, n47255, n47256,
n47257, n47258, n47259, n47260, n47261, n47262, n47263, n47264,
n47265, n47266, n47267, n47268, n47269, n47270, n47271, n47272,
n47273, n47274, n47275, n47276, n47277, n47278, n47279, n47280,
n47281, n47282, n47283, n47284, n47285, n47286, n47287, n47288,
n47289, n47290, n47291, n47292, n47293, n47294, n47295, n47296,
n47297, n47298, n47299, n47300, n47301, n47302, n47303, n47304,
n47305, n47306, n47307, n47308, n47309, n47310, n47311, n47312,
n47313, n47314, n47315, n47316, n47317, n47318, n47319, n47320,
n47321, n47322, n47323, n47324, n47325, n47326, n47327, n47328,
n47329, n47330, n47331, n47332, n47333, n47334, n47335, n47336,
n47337, n47338, n47339, n47340, n47341, n47342, n47343, n47344,
n47345, n47346, n47347, n47348, n47349, n47350, n47351, n47352,
n47353, n47354, n47355, n47356, n47357, n47358, n47359, n47360,
n47361, n47362, n47363, n47364, n47365, n47366, n47367, n47368,
n47369, n47370, n47371, n47372, n47373, n47374, n47375, n47376,
n47377, n47378, n47379, n47380, n47381, n47382, n47383, n47384,
n47385, n47386, n47387, n47388, n47389, n47390, n47391, n47392,
n47393, n47394, n47395, n47396, n47397, n47398, n47399, n47400,
n47401, n47402, n47403, n47404, n47405, n47406, n47407, n47408,
n47409, n47410, n47411, n47412, n47413, n47414, n47415, n47416,
n47417, n47418, n47419, n47420, n47421, n47422, n47423, n47424,
n47425, n47426, n47427, n47428, n47429, n47430, n47431, n47432,
n47433, n47434, n47435, n47436, n47437, n47438, n47439, n47440,
n47441, n47442, n47443, n47444, n47445, n47446, n47447, n47448,
n47449, n47450, n47451, n47452, n47453, n47454, n47455, n47456,
n47457, n47458, n47459, n47460, n47461, n47462, n47463, n47464,
n47465, n47466, n47467, n47468, n47469, n47470, n47471, n47472,
n47473, n47474, n47475, n47476, n47477, n47478, n47479, n47480,
n47481, n47482, n47483, n47484, n47485, n47486, n47487, n47488,
n47489, n47490, n47491, n47492, n47493, n47494, n47495, n47496,
n47497, n47498, n47499, n47500, n47501, n47502, n47503, n47504,
n47505, n47506, n47507, n47508, n47509, n47510, n47511, n47512,
n47513, n47514, n47515, n47516, n47517, n47518, n47519, n47520,
n47521, n47522, n47523, n47524, n47525, n47526, n47527, n47528,
n47529, n47530, n47531, n47532, n47533, n47534, n47535, n47536,
n47537, n47538, n47539, n47540, n47541, n47542, n47543, n47544,
n47545, n47546, n47547, n47548, n47549, n47550, n47551, n47552,
n47553, n47554, n47555, n47556, n47557, n47558, n47559, n47560,
n47561, n47562, n47563, n47564, n47565, n47566, n47567, n47568,
n47569, n47570, n47571, n47572, n47573, n47574, n47575, n47576,
n47577, n47578, n47579, n47580, n47581, n47582, n47583, n47584,
n47585, n47586, n47587, n47588, n47589, n47590, n47591, n47592,
n47593, n47594, n47595, n47596, n47597, n47598, n47599, n47600,
n47601, n47602, n47603, n47604, n47605, n47606, n47607, n47608,
n47609, n47610, n47611, n47612, n47613, n47614, n47615, n47616,
n47617, n47618, n47619, n47620, n47621, n47622, n47623, n47624,
n47625, n47626, n47627, n47628, n47629, n47630, n47631, n47632,
n47633, n47634, n47635, n47636, n47637, n47638, n47639, n47640,
n47641, n47642, n47643, n47644, n47645, n47646, n47647, n47648,
n47649, n47650, n47651, n47652, n47653, n47654, n47655, n47656,
n47657, n47658, n47659, n47660, n47661, n47662, n47663, n47664,
n47665, n47666, n47667, n47668, n47669, n47670, n47671, n47672,
n47673, n47674, n47675, n47676, n47677, n47678, n47679, n47680,
n47681, n47682, n47683, n47684, n47685, n47686, n47687, n47688,
n47689, n47690, n47691, n47692, n47693, n47694, n47695, n47696,
n47697, n47698, n47699, n47700, n47701, n47702, n47703, n47704,
n47705, n47706, n47707, n47708, n47709, n47710, n47711, n47712,
n47713, n47714, n47715, n47716, n47717, n47718, n47719, n47720,
n47721, n47722, n47723, n47724, n47725, n47726, n47727, n47728,
n47729, n47730, n47731, n47732, n47733, n47734, n47735, n47736,
n47737, n47738, n47739, n47740, n47741, n47742, n47743, n47744,
n47745, n47746, n47747, n47748, n47749, n47750, n47751, n47752,
n47753, n47754, n47755, n47756, n47757, n47758, n47759, n47760,
n47761, n47762, n47763, n47764, n47765, n47766, n47767, n47768,
n47769, n47770, n47771, n47772, n47773, n47774, n47775, n47776,
n47777, n47778, n47779, n47780, n47781, n47782, n47783, n47784,
n47785, n47786, n47787, n47788, n47789, n47790, n47791, n47792,
n47793, n47794, n47795, n47796, n47797, n47798, n47799, n47800,
n47801, n47802, n47803, n47804, n47805, n47806, n47807, n47808,
n47809, n47810, n47811, n47812, n47813, n47814, n47815, n47816,
n47817, n47818, n47819, n47820, n47821, n47822, n47823, n47824,
n47825, n47826, n47827, n47828, n47829, n47830, n47831, n47832,
n47833, n47834, n47835, n47836, n47837, n47838, n47839, n47840,
n47841, n47842, n47843, n47844, n47845, n47846, n47847, n47848,
n47849, n47850, n47851, n47852, n47853, n47854, n47855, n47856,
n47857, n47858, n47859, n47860, n47861, n47862, n47863, n47864,
n47865, n47866, n47867, n47868, n47869, n47870, n47871, n47872,
n47873, n47874, n47875, n47876, n47877, n47878, n47879, n47880,
n47881, n47882, n47883, n47884, n47885, n47886, n47887, n47888,
n47889, n47890, n47891, n47892, n47893, n47894, n47895, n47896,
n47897, n47898, n47899, n47900, n47901, n47902, n47903, n47904,
n47905, n47906, n47907, n47908, n47909, n47910, n47911, n47912,
n47913, n47914, n47915, n47916, n47917, n47918, n47919, n47920,
n47921, n47922, n47923, n47924, n47925, n47926, n47927, n47928,
n47929, n47930, n47931, n47932, n47933, n47934, n47935, n47936,
n47937, n47938, n47939, n47940, n47941, n47942, n47943, n47944,
n47945, n47946, n47947, n47948, n47949, n47950, n47951, n47952,
n47953, n47954, n47955, n47956, n47957, n47958, n47959, n47960,
n47961, n47962, n47963, n47964, n47965, n47966, n47967, n47968,
n47969, n47970, n47971, n47972, n47973, n47974, n47975, n47976,
n47977, n47978, n47979, n47980, n47981, n47982, n47983, n47984,
n47985, n47986, n47987, n47988, n47989, n47990, n47991, n47992,
n47993, n47994, n47995, n47996, n47997, n47998, n47999, n48000,
n48001, n48002, n48003, n48004, n48005, n48006, n48007, n48008,
n48009, n48010, n48011, n48012, n48013, n48014, n48015, n48016,
n48017, n48018, n48019, n48020, n48021, n48022, n48023, n48024,
n48025, n48026, n48027, n48028, n48029, n48030, n48031, n48032,
n48033, n48034, n48035, n48036, n48037, n48038, n48039, n48040,
n48041, n48042, n48043, n48044, n48045, n48046, n48047, n48048,
n48049, n48050, n48051, n48052, n48053, n48054, n48055, n48056,
n48057, n48058, n48059, n48060, n48061, n48062, n48063, n48064,
n48065, n48066, n48067, n48068, n48069, n48070, n48071, n48072,
n48073, n48074, n48075, n48076, n48077, n48078, n48079, n48080,
n48081, n48082, n48083, n48084, n48085, n48086, n48087, n48088,
n48089, n48090, n48091, n48092, n48093, n48094, n48095, n48096,
n48097, n48098, n48099, n48100, n48101, n48102, n48103, n48104,
n48105, n48106, n48107, n48108, n48109, n48110, n48111, n48112,
n48113, n48114, n48115, n48116, n48117, n48118, n48119, n48120,
n48121, n48122, n48123, n48124, n48125, n48126, n48127, n48128,
n48129, n48130, n48131, n48132, n48133, n48134, n48135, n48136,
n48137, n48138, n48139, n48140, n48141, n48142, n48143, n48144,
n48145, n48146, n48147, n48148, n48149, n48150, n48151, n48152,
n48153, n48154, n48155, n48156, n48157, n48158, n48159, n48160,
n48161, n48162, n48163, n48164, n48165, n48166, n48167, n48168,
n48169, n48170, n48171, n48172, n48173, n48174, n48175, n48176,
n48177, n48178, n48179, n48180, n48181, n48182, n48183, n48184,
n48185, n48186, n48187, n48188, n48189, n48190, n48191, n48192,
n48193, n48194, n48195, n48196, n48197, n48198, n48199, n48200,
n48201, n48202, n48203, n48204, n48205, n48206, n48207, n48208,
n48209, n48210, n48211, n48212, n48213, n48214, n48215, n48216,
n48217, n48218, n48219, n48220, n48221, n48222, n48223, n48224,
n48225, n48226, n48227, n48228, n48229, n48230, n48231, n48232,
n48233, n48234, n48235, n48236, n48237, n48238, n48239, n48240,
n48241, n48242, n48243, n48244, n48245, n48246, n48247, n48248,
n48249, n48250, n48251, n48252, n48253, n48254, n48255, n48256,
n48257, n48258, n48259, n48260, n48261, n48262, n48263, n48264,
n48265, n48266, n48267, n48268, n48269, n48270, n48271, n48272,
n48273, n48274, n48275, n48276, n48277, n48278, n48279, n48280,
n48281, n48282, n48283, n48284, n48285, n48286, n48287, n48288,
n48289, n48290, n48291, n48292, n48293, n48294, n48295, n48296,
n48297, n48298, n48299, n48300, n48301, n48302, n48303, n48304,
n48305, n48306, n48307, n48308, n48309, n48310, n48311, n48312,
n48313, n48314, n48315, n48316, n48317, n48318, n48319, n48320,
n48321, n48322, n48323, n48324, n48325, n48326, n48327, n48328,
n48329, n48330, n48331, n48332, n48333, n48334, n48335, n48336,
n48337, n48338, n48339, n48340, n48341, n48342, n48343, n48344,
n48345, n48346, n48347, n48348, n48349, n48350, n48351, n48352,
n48353, n48354, n48355, n48356, n48357, n48358, n48359, n48360,
n48361, n48362, n48363, n48364, n48365, n48366, n48367, n48368,
n48369, n48370, n48371, n48372, n48373, n48374, n48375, n48376,
n48377, n48378, n48379, n48380, n48381, n48382, n48383, n48384,
n48385, n48386, n48387, n48388, n48389, n48390, n48391, n48392,
n48393, n48394, n48395, n48396, n48397, n48398, n48399, n48400,
n48401, n48402, n48403, n48404, n48405, n48406, n48407, n48408,
n48409, n48410, n48411, n48412, n48413, n48414, n48415, n48416,
n48417, n48418, n48419, n48420, n48421, n48422, n48423, n48424,
n48425, n48426, n48427, n48428, n48429, n48430, n48431, n48432,
n48433, n48434, n48435, n48436, n48437, n48438, n48439, n48440,
n48441, n48442, n48443, n48444, n48445, n48446, n48447, n48448,
n48449, n48450, n48451, n48452, n48453, n48454, n48455, n48456,
n48457, n48458, n48459, n48460, n48461, n48462, n48463, n48464,
n48465, n48466, n48467, n48468, n48469, n48470, n48471, n48472,
n48473, n48474, n48475, n48476, n48477, n48478, n48479, n48480,
n48481, n48482, n48483, n48484, n48485, n48486, n48487, n48488,
n48489, n48490, n48491, n48492, n48493, n48494, n48495, n48496,
n48497, n48498, n48499, n48500, n48501, n48502, n48503, n48504,
n48505, n48506, n48507, n48508, n48509, n48510, n48511, n48512,
n48513, n48514, n48515, n48516, n48517, n48518, n48519, n48520,
n48521, n48522, n48523, n48524, n48525, n48526, n48527, n48528,
n48529, n48530, n48531, n48532, n48533, n48534, n48535, n48536,
n48537, n48538, n48539, n48540, n48541, n48542, n48543, n48544,
n48545, n48546, n48547, n48548, n48549, n48550, n48551, n48552,
n48553, n48554, n48555, n48556, n48557, n48558, n48559, n48560,
n48561, n48562, n48563, n48564, n48565, n48566, n48567, n48568,
n48569, n48570, n48571, n48572, n48573, n48574, n48575, n48576,
n48577, n48578, n48579, n48580, n48581, n48582, n48583, n48584,
n48585, n48586, n48587, n48588, n48589, n48590, n48591, n48592,
n48593, n48594, n48595, n48596, n48597, n48598, n48599, n48600,
n48601, n48602, n48603, n48604, n48605, n48606, n48607, n48608,
n48609, n48610, n48611, n48612, n48613, n48614, n48615, n48616,
n48617, n48618, n48619, n48620, n48621, n48622, n48623, n48624,
n48625, n48626, n48627, n48628, n48629, n48630, n48631, n48632,
n48633, n48634, n48635, n48636, n48637, n48638, n48639, n48640,
n48641, n48642, n48643, n48644, n48645, n48646, n48647, n48648,
n48649, n48650, n48651, n48652, n48653, n48654, n48655, n48656,
n48657, n48658, n48659, n48660, n48661, n48662, n48663, n48664,
n48665, n48666, n48667, n48668, n48669, n48670, n48671, n48672,
n48673, n48674, n48675, n48676, n48677, n48678, n48679, n48680,
n48681, n48682, n48683, n48684, n48685, n48686, n48687, n48688,
n48689, n48690, n48691, n48692, n48693, n48694, n48695, n48696,
n48697, n48698, n48699, n48700, n48701, n48702, n48703, n48704,
n48705, n48706, n48707, n48708, n48709, n48710, n48711, n48712,
n48713, n48714, n48715, n48716, n48717, n48718, n48719, n48720,
n48721, n48722, n48723, n48724, n48725, n48726, n48727, n48728,
n48729, n48730, n48731, n48732, n48733, n48734, n48735, n48736,
n48737, n48738, n48739, n48740, n48741, n48742, n48743, n48744,
n48745, n48746, n48747, n48748, n48749, n48750, n48751, n48752,
n48753, n48754, n48755, n48756, n48757, n48758, n48759, n48760,
n48761, n48762, n48763, n48764, n48765, n48766, n48767, n48768,
n48769, n48770, n48771, n48772, n48773, n48774, n48775, n48776,
n48777, n48778, n48779, n48780, n48781, n48782, n48783, n48784,
n48785, n48786, n48787, n48788, n48789, n48790, n48791, n48792,
n48793, n48794, n48795, n48796, n48797, n48798, n48799, n48800,
n48801, n48802, n48803, n48804, n48805, n48806, n48807, n48808,
n48809, n48810, n48811, n48812, n48813, n48814, n48815, n48816,
n48817, n48818, n48819, n48820, n48821, n48822, n48823, n48824,
n48825, n48826, n48827, n48828, n48829, n48830, n48831, n48832,
n48833, n48834, n48835, n48836, n48837, n48838, n48839, n48840,
n48841, n48842, n48843, n48844, n48845, n48846, n48847, n48848,
n48849, n48850, n48851, n48852, n48853, n48854, n48855, n48856,
n48857, n48858, n48859, n48860, n48861, n48862, n48863, n48864,
n48865, n48866, n48867, n48868, n48869, n48870, n48871, n48872,
n48873, n48874, n48875, n48876, n48877, n48878, n48879, n48880,
n48881, n48882, n48883, n48884, n48885, n48886, n48887, n48888,
n48889, n48890, n48891, n48892, n48893, n48894, n48895, n48896,
n48897, n48898, n48899, n48900, n48901, n48902, n48903, n48904,
n48905, n48906, n48907, n48908, n48909, n48910, n48911, n48912,
n48913, n48914, n48915, n48916, n48917, n48918, n48919, n48920,
n48921, n48922, n48923, n48924, n48925, n48926, n48927, n48928,
n48929, n48930, n48931, n48932, n48933, n48934, n48935, n48936,
n48937, n48938, n48939, n48940, n48941, n48942, n48943, n48944,
n48945, n48946, n48947, n48948, n48949, n48950, n48951, n48952,
n48953, n48954, n48955, n48956, n48957, n48958, n48959, n48960,
n48961, n48962, n48963, n48964, n48965, n48966, n48967, n48968,
n48969, n48970, n48971, n48972, n48973, n48974, n48975, n48976,
n48977, n48978, n48979, n48980, n48981, n48982, n48983, n48984,
n48985, n48986, n48987, n48988, n48989, n48990, n48991, n48992,
n48993, n48994, n48995, n48996, n48997, n48998, n48999, n49000,
n49001, n49002, n49003, n49004, n49005, n49006, n49007, n49008,
n49009, n49010, n49011, n49012, n49013, n49014, n49015, n49016,
n49017, n49018, n49019, n49020, n49021, n49022, n49023, n49024,
n49025, n49026, n49027, n49028, n49029, n49030, n49031, n49032,
n49033, n49034, n49035, n49036, n49037, n49038, n49039, n49040,
n49041, n49042, n49043, n49044, n49045, n49046, n49047, n49048,
n49049, n49050, n49051, n49052, n49053, n49054, n49055, n49056,
n49057, n49058, n49059, n49060, n49061, n49062, n49063, n49064,
n49065, n49066, n49067, n49068, n49069, n49070, n49071, n49072,
n49073, n49074, n49075, n49076, n49077, n49078, n49079, n49080,
n49081, n49082, n49083, n49084, n49085, n49086, n49087, n49088,
n49089, n49090, n49091, n49092, n49093, n49094, n49095, n49096,
n49097, n49098, n49099, n49100, n49101, n49102, n49103, n49104,
n49105, n49106, n49107, n49108, n49109, n49110, n49111, n49112,
n49113, n49114, n49115, n49116, n49117, n49118, n49119, n49120,
n49121, n49122, n49123, n49124, n49125, n49126, n49127, n49128,
n49129, n49130, n49131, n49132, n49133, n49134, n49135, n49136,
n49137, n49138, n49139, n49140, n49141, n49142, n49143, n49144,
n49145, n49146, n49147, n49148, n49149, n49150, n49151, n49152,
n49153, n49154, n49155, n49156, n49157, n49158, n49159, n49160,
n49161, n49162, n49163, n49164, n49165, n49166, n49167, n49168,
n49169, n49170, n49171, n49172, n49173, n49174, n49175, n49176,
n49177, n49178, n49179, n49180, n49181, n49182, n49183, n49184,
n49185, n49186, n49187, n49188, n49189, n49190, n49191, n49192,
n49193, n49194, n49195, n49196, n49197, n49198, n49199, n49200,
n49201, n49202, n49203, n49204, n49205, n49206, n49207, n49208,
n49209, n49210, n49211, n49212, n49213, n49214, n49215, n49216,
n49217, n49218, n49219, n49220, n49221, n49222, n49223, n49224,
n49225, n49226, n49227, n49228, n49229, n49230, n49231, n49232,
n49233, n49234, n49235, n49236, n49237, n49238, n49239, n49240,
n49241, n49242, n49243, n49244, n49245, n49246, n49247, n49248,
n49249, n49250, n49251, n49252, n49253, n49254, n49255, n49256,
n49257, n49258, n49259, n49260, n49261, n49262, n49263, n49264,
n49265, n49266, n49267, n49268, n49269, n49270, n49271, n49272,
n49273, n49274, n49275, n49276, n49277, n49278, n49279, n49280,
n49281, n49282, n49283, n49284, n49285, n49286, n49287, n49288,
n49289, n49290, n49291, n49292, n49293, n49294, n49295, n49296,
n49297, n49298, n49299, n49300, n49301, n49302, n49303, n49304,
n49305, n49306, n49307, n49308, n49309, n49310, n49311, n49312,
n49313, n49314, n49315, n49316, n49317, n49318, n49319, n49320,
n49321, n49322, n49323, n49324, n49325, n49326, n49327, n49328,
n49329, n49330, n49331, n49332, n49333, n49334, n49335, n49336,
n49337, n49338, n49339, n49340, n49341, n49342, n49343, n49344,
n49345, n49346, n49347, n49348, n49349, n49350, n49351, n49352,
n49353, n49354, n49355, n49356, n49357, n49358, n49359, n49360,
n49361, n49362, n49363, n49364, n49365, n49366, n49367, n49368,
n49369, n49370, n49371, n49372, n49373, n49374, n49375, n49376,
n49377, n49378, n49379, n49380, n49381, n49382, n49383, n49384,
n49385, n49386, n49387, n49388, n49389, n49390, n49391, n49392,
n49393, n49394, n49395, n49396, n49397, n49398, n49399, n49400,
n49401, n49402, n49403, n49404, n49405, n49406, n49407, n49408,
n49409, n49410, n49411, n49412, n49413, n49414, n49415, n49416,
n49417, n49418, n49419, n49420, n49421, n49422, n49423, n49424,
n49425, n49426, n49427, n49428, n49429, n49430, n49431, n49432,
n49433, n49434, n49435, n49436, n49437, n49438, n49439, n49440,
n49441, n49442, n49443, n49444, n49445, n49446, n49447, n49448,
n49449, n49450, n49451, n49452, n49453, n49454, n49455, n49456,
n49457, n49458, n49459, n49460, n49461, n49462, n49463, n49464,
n49465, n49466, n49467, n49468, n49469, n49470, n49471, n49472,
n49473, n49474, n49475, n49476, n49477, n49478, n49479, n49480,
n49481, n49482, n49483, n49484, n49485, n49486, n49487, n49488,
n49489, n49490, n49491, n49492, n49493, n49494, n49495, n49496,
n49497, n49498, n49499, n49500, n49501, n49502, n49503, n49504,
n49505, n49506, n49507, n49508, n49509, n49510, n49511, n49512,
n49513, n49514, n49515, n49516, n49517, n49518, n49519, n49520,
n49521, n49522, n49523, n49524, n49525, n49526, n49527, n49528,
n49529, n49530, n49531, n49532, n49533, n49534, n49535, n49536,
n49537, n49538, n49539, n49540, n49541, n49542, n49543, n49544,
n49545, n49546, n49547, n49548, n49549, n49550, n49551, n49552,
n49553, n49554, n49555, n49556, n49557, n49558, n49559, n49560,
n49561, n49562, n49563, n49564, n49565, n49566, n49567, n49568,
n49569, n49570, n49571, n49572, n49573, n49574, n49575, n49576,
n49577, n49578, n49579, n49580, n49581, n49582, n49583, n49584,
n49585, n49586, n49587, n49588, n49589, n49590, n49591, n49592,
n49593, n49594, n49595, n49596, n49597, n49598, n49599, n49600,
n49601, n49602, n49603, n49604, n49605, n49606, n49607, n49608,
n49609, n49610, n49611, n49612, n49613, n49614, n49615, n49616,
n49617, n49618, n49619, n49620, n49621, n49622, n49623, n49624,
n49625, n49626, n49627, n49628, n49629, n49630, n49631, n49632,
n49633, n49634, n49635, n49636, n49637, n49638, n49639, n49640,
n49641, n49642, n49643, n49644, n49645, n49646, n49647, n49648,
n49649, n49650, n49651, n49652, n49653, n49654, n49655, n49656,
n49657, n49658, n49659, n49660, n49661, n49662, n49663, n49664,
n49665, n49666, n49667, n49668, n49669, n49670, n49671, n49672,
n49673, n49674, n49675, n49676, n49677, n49678, n49679, n49680,
n49681, n49682, n49683, n49684, n49685, n49686, n49687, n49688,
n49689, n49690, n49691, n49692, n49693, n49694, n49695, n49696,
n49697, n49698, n49699, n49700, n49701, n49702, n49703, n49704,
n49705, n49706, n49707, n49708, n49709, n49710, n49711, n49712,
n49713, n49714, n49715, n49716, n49717, n49718, n49719, n49720,
n49721, n49722, n49723, n49724, n49725, n49726, n49727, n49728,
n49729, n49730, n49731, n49732, n49733, n49734, n49735, n49736,
n49737, n49738, n49739, n49740, n49741, n49742, n49743, n49744,
n49745, n49746, n49747, n49748, n49749, n49750, n49751, n49752,
n49753, n49754, n49755, n49756, n49757, n49758, n49759, n49760,
n49761, n49762, n49763, n49764, n49765, n49766, n49767, n49768,
n49769, n49770, n49771, n49772, n49773, n49774, n49775, n49776,
n49777, n49778, n49779, n49780, n49781, n49782, n49783, n49784,
n49785, n49786, n49787, n49788, n49789, n49790, n49791, n49792,
n49793, n49794, n49795, n49796, n49797, n49798, n49799, n49800,
n49801, n49802, n49803, n49804, n49805, n49806, n49807, n49808,
n49809, n49810, n49811, n49812, n49813, n49814, n49815, n49816,
n49817, n49818, n49819, n49820, n49821, n49822, n49823, n49824,
n49825, n49826, n49827, n49828, n49829, n49830, n49831, n49832,
n49833, n49834, n49835, n49836, n49837, n49838, n49839, n49840,
n49841, n49842, n49843, n49844, n49845, n49846, n49847, n49848,
n49849, n49850, n49851, n49852, n49853, n49854, n49855, n49856,
n49857, n49858, n49859, n49860, n49861, n49862, n49863, n49864,
n49865, n49866, n49867, n49868, n49869, n49870, n49871, n49872,
n49873, n49874, n49875, n49876, n49877, n49878, n49879, n49880,
n49881, n49882, n49883, n49884, n49885, n49886, n49887, n49888,
n49889, n49890, n49891, n49892, n49893, n49894, n49895, n49896,
n49897, n49898, n49899, n49900, n49901, n49902, n49903, n49904,
n49905, n49906, n49907, n49908, n49909, n49910, n49911, n49912,
n49913, n49914, n49915, n49916, n49917, n49918, n49919, n49920,
n49921, n49922, n49923, n49924, n49925, n49926, n49927, n49928,
n49929, n49930, n49931, n49932, n49933, n49934, n49935, n49936,
n49937, n49938, n49939, n49940, n49941, n49942, n49943, n49944,
n49945, n49946, n49947, n49948, n49949, n49950, n49951, n49952,
n49953, n49954, n49955, n49956, n49957, n49958, n49959, n49960,
n49961, n49962, n49963, n49964, n49965, n49966, n49967, n49968,
n49969, n49970, n49971, n49972, n49973, n49974, n49975, n49976,
n49977, n49978, n49979, n49980, n49981, n49982, n49983, n49984,
n49985, n49986, n49987, n49988, n49989, n49990, n49991, n49992,
n49993, n49994, n49995, n49996, n49997, n49998, n49999, n50000,
n50001, n50002, n50003, n50004, n50005, n50006, n50007, n50008,
n50009, n50010, n50011, n50012, n50013, n50014, n50015, n50016,
n50017, n50018, n50019, n50020, n50021, n50022, n50023, n50024,
n50025, n50026, n50027, n50028, n50029, n50030, n50031, n50032,
n50033, n50034, n50035, n50036, n50037, n50038, n50039, n50040,
n50041, n50042, n50043, n50044, n50045, n50046, n50047, n50048,
n50049, n50050, n50051, n50052, n50053, n50054, n50055, n50056,
n50057, n50058, n50059, n50060, n50061, n50062, n50063, n50064,
n50065, n50066, n50067, n50068, n50069, n50070, n50071, n50072,
n50073, n50074, n50075, n50076, n50077, n50078, n50079, n50080,
n50081, n50082, n50083, n50084, n50085, n50086, n50087, n50088,
n50089, n50090, n50091, n50092, n50093, n50094, n50095, n50096,
n50097, n50098, n50099, n50100, n50101, n50102, n50103, n50104,
n50105, n50106, n50107, n50108, n50109, n50110, n50111, n50112,
n50113, n50114, n50115, n50116, n50117, n50118, n50119, n50120,
n50121, n50122, n50123, n50124, n50125, n50126, n50127, n50128,
n50129, n50130, n50131, n50132, n50133, n50134, n50135, n50136,
n50137, n50138, n50139, n50140, n50141, n50142, n50143, n50144,
n50145, n50146, n50147, n50148, n50149, n50150, n50151, n50152,
n50153, n50154, n50155, n50156, n50157, n50158, n50159, n50160,
n50161, n50162, n50163, n50164, n50165, n50166, n50167, n50168,
n50169, n50170, n50171, n50172, n50173, n50174, n50175, n50176,
n50177, n50178, n50179, n50180, n50181, n50182, n50183, n50184,
n50185, n50186, n50187, n50188, n50189, n50190, n50191, n50192,
n50193, n50194, n50195, n50196, n50197, n50198, n50199, n50200,
n50201, n50202, n50203, n50204, n50205, n50206, n50207, n50208,
n50209, n50210, n50211, n50212, n50213, n50214, n50215, n50216,
n50217, n50218, n50219, n50220, n50221, n50222, n50223, n50224,
n50225, n50226, n50227, n50228, n50229, n50230, n50231, n50232,
n50233, n50234, n50235, n50236, n50237, n50238, n50239, n50240,
n50241, n50242, n50243, n50244, n50245, n50246, n50247, n50248,
n50249, n50250, n50251, n50252, n50253, n50254, n50255, n50256,
n50257, n50258, n50259, n50260, n50261, n50262, n50263, n50264,
n50265, n50266, n50267, n50268, n50269, n50270, n50271, n50272,
n50273, n50274, n50275, n50276, n50277, n50278, n50279, n50280,
n50281, n50282, n50283, n50284, n50285, n50286, n50287, n50288,
n50289, n50290, n50291, n50292, n50293, n50294, n50295, n50296,
n50297, n50298, n50299, n50300, n50301, n50302, n50303, n50304,
n50305, n50306, n50307, n50308, n50309, n50310, n50311, n50312,
n50313, n50314, n50315, n50316, n50317, n50318, n50319, n50320,
n50321, n50322, n50323, n50324, n50325, n50326, n50327, n50328,
n50329, n50330, n50331, n50332, n50333, n50334, n50335, n50336,
n50337, n50338, n50339, n50340, n50341, n50342, n50343, n50344,
n50345, n50346, n50347, n50348, n50349, n50350, n50351, n50352,
n50353, n50354, n50355, n50356, n50357, n50358, n50359, n50360,
n50361, n50362, n50363, n50364, n50365, n50366, n50367, n50368,
n50369, n50370, n50371, n50372, n50373, n50374, n50375, n50376,
n50377, n50378, n50379, n50380, n50381, n50382, n50383, n50384,
n50385, n50386, n50387, n50388, n50389, n50390, n50391, n50392,
n50393, n50394, n50395, n50396, n50397, n50398, n50399, n50400,
n50401, n50402, n50403, n50404, n50405, n50406, n50407, n50408,
n50409, n50410, n50411, n50412, n50413, n50414, n50415, n50416,
n50417, n50418, n50419, n50420, n50421, n50422, n50423, n50424,
n50425, n50426, n50427, n50428, n50429, n50430, n50431, n50432,
n50433, n50434, n50435, n50436, n50437, n50438, n50439, n50440,
n50441, n50442, n50443, n50444, n50445, n50446, n50447, n50448,
n50449, n50450, n50451, n50452, n50453, n50454, n50455, n50456,
n50457, n50458, n50459, n50460, n50461, n50462, n50463, n50464,
n50465, n50466, n50467, n50468, n50469, n50470, n50471, n50472,
n50473, n50474, n50475, n50476, n50477, n50478, n50479, n50480,
n50481, n50482, n50483, n50484, n50485, n50486, n50487, n50488,
n50489, n50490, n50491, n50492, n50493, n50494, n50495, n50496,
n50497, n50498, n50499, n50500, n50501, n50502, n50503, n50504,
n50505, n50506, n50507, n50508, n50509, n50510, n50511, n50512,
n50513, n50514, n50515, n50516, n50517, n50518, n50519, n50520,
n50521, n50522, n50523, n50524, n50525, n50526, n50527, n50528,
n50529, n50530, n50531, n50532, n50533, n50534, n50535, n50536,
n50537, n50538, n50539, n50540, n50541, n50542, n50543, n50544,
n50545, n50546, n50547, n50548, n50549, n50550, n50551, n50552,
n50553, n50554, n50555, n50556, n50557, n50558, n50559, n50560,
n50561, n50562, n50563, n50564, n50565, n50566, n50567, n50568,
n50569, n50570, n50571, n50572, n50573, n50574, n50575, n50576,
n50577, n50578, n50579, n50580, n50581, n50582, n50583, n50584,
n50585, n50586, n50587, n50588, n50589, n50590, n50591, n50592,
n50593, n50594, n50595, n50596, n50597, n50598, n50599, n50600,
n50601, n50602, n50603, n50604, n50605, n50606, n50607, n50608,
n50609, n50610, n50611, n50612, n50613, n50614, n50615, n50616,
n50617, n50618, n50619, n50620, n50621, n50622, n50623, n50624,
n50625, n50626, n50627, n50628, n50629, n50630, n50631, n50632,
n50633, n50634, n50635, n50636, n50637, n50638, n50639, n50640,
n50641, n50642, n50643, n50644, n50645, n50646, n50647, n50648,
n50649, n50650, n50651, n50652, n50653, n50654, n50655, n50656,
n50657, n50658, n50659, n50660, n50661, n50662, n50663, n50664,
n50665, n50666, n50667, n50668, n50669, n50670, n50671, n50672,
n50673, n50674, n50675, n50676, n50677, n50678, n50679, n50680,
n50681, n50682, n50683, n50684, n50685, n50686, n50687, n50688,
n50689, n50690, n50691, n50692, n50693, n50694, n50695, n50696,
n50697, n50698, n50699, n50700, n50701, n50702, n50703, n50704,
n50705, n50706, n50707, n50708, n50709, n50710, n50711, n50712,
n50713, n50714, n50715, n50716, n50717, n50718, n50719, n50720,
n50721, n50722, n50723, n50724, n50725, n50726, n50727, n50728,
n50729, n50730, n50731, n50732, n50733, n50734, n50735, n50736,
n50737, n50738, n50739, n50740, n50741, n50742, n50743, n50744,
n50745, n50746, n50747, n50748, n50749, n50750, n50751, n50752,
n50753, n50754, n50755, n50756, n50757, n50758, n50759, n50760,
n50761, n50762, n50763, n50764, n50765, n50766, n50767, n50768,
n50769, n50770, n50771, n50772, n50773, n50774, n50775, n50776,
n50777, n50778, n50779, n50780, n50781, n50782, n50783, n50784,
n50785, n50786, n50787, n50788, n50789, n50790, n50791, n50792,
n50793, n50794, n50795, n50796, n50797, n50798, n50799, n50800,
n50801, n50802, n50803, n50804, n50805, n50806, n50807, n50808,
n50809, n50810, n50811, n50812, n50813, n50814, n50815, n50816,
n50817, n50818, n50819, n50820, n50821, n50822, n50823, n50824,
n50825, n50826, n50827, n50828, n50829, n50830, n50831, n50832,
n50833, n50834, n50835, n50836, n50837, n50838, n50839, n50840,
n50841, n50842, n50843, n50844, n50845, n50846, n50847, n50848,
n50849, n50850, n50851, n50852, n50853, n50854, n50855, n50856,
n50857, n50858, n50859, n50860, n50861, n50862, n50863, n50864,
n50865, n50866, n50867, n50868, n50869, n50870, n50871, n50872,
n50873, n50874, n50875, n50876, n50877, n50878, n50879, n50880,
n50881, n50882, n50883, n50884, n50885, n50886, n50887, n50888,
n50889, n50890, n50891, n50892, n50893, n50894, n50895, n50896,
n50897, n50898, n50899, n50900, n50901, n50902, n50903, n50904,
n50905, n50906, n50907, n50908, n50909, n50910, n50911, n50912,
n50913, n50914, n50915, n50916, n50917, n50918, n50919, n50920,
n50921, n50922, n50923, n50924, n50925, n50926, n50927, n50928,
n50929, n50930, n50931, n50932, n50933, n50934, n50935, n50936,
n50937, n50938, n50939, n50940, n50941, n50942, n50943, n50944,
n50945, n50946, n50947, n50948, n50949, n50950, n50951, n50952,
n50953, n50954, n50955, n50956, n50957, n50958, n50959, n50960,
n50961, n50962, n50963, n50964, n50965, n50966, n50967, n50968,
n50969, n50970, n50971, n50972, n50973, n50974, n50975, n50976,
n50977, n50978, n50979, n50980, n50981, n50982, n50983, n50984,
n50985, n50986, n50987, n50988, n50989, n50990, n50991, n50992,
n50993, n50994, n50995, n50996, n50997, n50998, n50999, n51000,
n51001, n51002, n51003, n51004, n51005, n51006, n51007, n51008,
n51009, n51010, n51011, n51012, n51013, n51014, n51015, n51016,
n51017, n51018, n51019, n51020, n51021, n51022, n51023, n51024,
n51025, n51026, n51027, n51028, n51029, n51030, n51031, n51032,
n51033, n51034, n51035, n51036, n51037, n51038, n51039, n51040,
n51041, n51042, n51043, n51044, n51045, n51046, n51047, n51048,
n51049, n51050, n51051, n51052, n51053, n51054, n51055, n51056,
n51057, n51058, n51059, n51060, n51061, n51062, n51063, n51064,
n51065, n51066, n51067, n51068, n51069, n51070, n51071, n51072,
n51073, n51074, n51075, n51076, n51077, n51078, n51079, n51080,
n51081, n51082, n51083, n51084, n51085, n51086, n51087, n51088,
n51089, n51090, n51091, n51092, n51093, n51094, n51095, n51096,
n51097, n51098, n51099, n51100, n51101, n51102, n51103, n51104,
n51105, n51106, n51107, n51108, n51109, n51110, n51111, n51112,
n51113, n51114, n51115, n51116, n51117, n51118, n51119, n51120,
n51121, n51122, n51123, n51124, n51125, n51126, n51127, n51128,
n51129, n51130, n51131, n51132, n51133, n51134, n51135, n51136,
n51137, n51138, n51139, n51140, n51141, n51142, n51143, n51144,
n51145, n51146, n51147, n51148, n51149, n51150, n51151, n51152,
n51153, n51154, n51155, n51156, n51157, n51158, n51159, n51160,
n51161, n51162, n51163, n51164, n51165, n51166, n51167, n51168,
n51169, n51170, n51171, n51172, n51173, n51174, n51175, n51176,
n51177, n51178, n51179, n51180, n51181, n51182, n51183, n51184,
n51185, n51186, n51187, n51188, n51189, n51190, n51191, n51192,
n51193, n51194, n51195, n51196, n51197, n51198, n51199, n51200,
n51201, n51202, n51203, n51204, n51205, n51206, n51207, n51208,
n51209, n51210, n51211, n51212, n51213, n51214, n51215, n51216,
n51217, n51218, n51219, n51220, n51221, n51222, n51223, n51224,
n51225, n51226, n51227, n51228, n51229, n51230, n51231, n51232,
n51233, n51234, n51235, n51236, n51237, n51238, n51239, n51240,
n51241, n51242, n51243, n51244, n51245, n51246, n51247, n51248,
n51249, n51250, n51251, n51252, n51253, n51254, n51255, n51256,
n51257, n51258, n51259, n51260, n51261, n51262, n51263, n51264,
n51265, n51266, n51267, n51268, n51269, n51270, n51271, n51272,
n51273, n51274, n51275, n51276, n51277, n51278, n51279, n51280,
n51281, n51282, n51283, n51284, n51285, n51286, n51287, n51288,
n51289, n51290, n51291, n51292, n51293, n51294, n51295, n51296,
n51297, n51298, n51299, n51300, n51301, n51302, n51303, n51304,
n51305, n51306, n51307, n51308, n51309, n51310, n51311, n51312,
n51313, n51314, n51315, n51316, n51317, n51318, n51319, n51320,
n51321, n51322, n51323, n51324, n51325, n51326, n51327, n51328,
n51329, n51330, n51331, n51332, n51333, n51334, n51335, n51336,
n51337, n51338, n51339, n51340, n51341, n51342, n51343, n51344,
n51345, n51346, n51347, n51348, n51349, n51350, n51351, n51352,
n51353, n51354, n51355, n51356, n51357, n51358, n51359, n51360,
n51361, n51362, n51363, n51364, n51365, n51366, n51367, n51368,
n51369, n51370, n51371, n51372, n51373, n51374, n51375, n51376,
n51377, n51378, n51379, n51380, n51381, n51382, n51383, n51384,
n51385, n51386, n51387, n51388, n51389, n51390, n51391, n51392,
n51393, n51394, n51395, n51396, n51397, n51398, n51399, n51400,
n51401, n51402, n51403, n51404, n51405, n51406, n51407, n51408,
n51409, n51410, n51411, n51412, n51413, n51414, n51415, n51416,
n51417, n51418, n51419, n51420, n51421, n51422, n51423, n51424,
n51425, n51426, n51427, n51428, n51429, n51430, n51431, n51432,
n51433, n51434, n51435, n51436, n51437, n51438, n51439, n51440,
n51441, n51442, n51443, n51444, n51445, n51446, n51447, n51448,
n51449, n51450, n51451, n51452, n51453, n51454, n51455, n51456,
n51457, n51458, n51459, n51460, n51461, n51462, n51463, n51464,
n51465, n51466, n51467, n51468, n51469, n51470, n51471, n51472,
n51473, n51474, n51475, n51476, n51477, n51478, n51479, n51480,
n51481, n51482, n51483, n51484, n51485, n51486, n51487, n51488,
n51489, n51490, n51491, n51492, n51493, n51494, n51495, n51496,
n51497, n51498, n51499, n51500, n51501, n51502, n51503, n51504,
n51505, n51506, n51507, n51508, n51509, n51510, n51511, n51512,
n51513, n51514, n51515, n51516, n51517, n51518, n51519, n51520,
n51521, n51522, n51523, n51524, n51525, n51526, n51527, n51528,
n51529, n51530, n51531, n51532, n51533, n51534, n51535, n51536,
n51537, n51538, n51539, n51540, n51541, n51542, n51543, n51544,
n51545, n51546, n51547, n51548, n51549, n51550, n51551, n51552,
n51553, n51554, n51555, n51556, n51557, n51558, n51559, n51560,
n51561, n51562, n51563, n51564, n51565, n51566, n51567, n51568,
n51569, n51570, n51571, n51572, n51573, n51574, n51575, n51576,
n51577, n51578, n51579, n51580, n51581, n51582, n51583, n51584,
n51585, n51586, n51587, n51588, n51589, n51590, n51591, n51592,
n51593, n51594, n51595, n51596, n51597, n51598, n51599, n51600,
n51601, n51602, n51603, n51604, n51605, n51606, n51607, n51608,
n51609, n51610, n51611, n51612, n51613, n51614, n51615, n51616,
n51617, n51618, n51619, n51620, n51621, n51622, n51623, n51624,
n51625, n51626, n51627, n51628, n51629, n51630, n51631, n51632,
n51633, n51634, n51635, n51636, n51637, n51638, n51639, n51640,
n51641, n51642, n51643, n51644, n51645, n51646, n51647, n51648,
n51649, n51650, n51651, n51652, n51653, n51654, n51655, n51656,
n51657, n51658, n51659, n51660, n51661, n51662, n51663, n51664,
n51665, n51666, n51667, n51668, n51669, n51670, n51671, n51672,
n51673, n51674, n51675, n51676, n51677, n51678, n51679, n51680,
n51681, n51682, n51683, n51684, n51685, n51686, n51687, n51688,
n51689, n51690, n51691, n51692, n51693, n51694, n51695, n51696,
n51697, n51698, n51699, n51700, n51701, n51702, n51703, n51704,
n51705, n51706, n51707, n51708, n51709, n51710, n51711, n51712,
n51713, n51714, n51715, n51716, n51717, n51718, n51719, n51720,
n51721, n51722, n51723, n51724, n51725, n51726, n51727, n51728,
n51729, n51730, n51731, n51732, n51733, n51734, n51735, n51736,
n51737, n51738, n51739, n51740, n51741, n51742, n51743, n51744,
n51745, n51746, n51747, n51748, n51749, n51750, n51751, n51752,
n51753, n51754, n51755, n51756, n51757, n51758, n51759, n51760,
n51761, n51762, n51763, n51764, n51765, n51766, n51767, n51768,
n51769, n51770, n51771, n51772, n51773, n51774, n51775, n51776,
n51777, n51778, n51779, n51780, n51781, n51782, n51783, n51784,
n51785, n51786, n51787, n51788, n51789, n51790, n51791, n51792,
n51793, n51794, n51795, n51796, n51797, n51798, n51799, n51800,
n51801, n51802, n51803, n51804, n51805, n51806, n51807, n51808,
n51809, n51810, n51811, n51812, n51813, n51814, n51815, n51816,
n51817, n51818, n51819, n51820, n51821, n51822, n51823, n51824,
n51825, n51826, n51827, n51828, n51829, n51830, n51831, n51832,
n51833, n51834, n51835, n51836, n51837, n51838, n51839, n51840,
n51841, n51842, n51843, n51844, n51845, n51846, n51847, n51848,
n51849, n51850, n51851, n51852, n51853, n51854, n51855, n51856,
n51857, n51858, n51859, n51860, n51861, n51862, n51863, n51864,
n51865, n51866, n51867, n51868, n51869, n51870, n51871, n51872,
n51873, n51874, n51875, n51876, n51877, n51878, n51879, n51880,
n51881, n51882, n51883, n51884, n51885, n51886, n51887, n51888,
n51889, n51890, n51891, n51892, n51893, n51894, n51895, n51896,
n51897, n51898, n51899, n51900, n51901, n51902, n51903, n51904,
n51905, n51906, n51907, n51908, n51909, n51910, n51911, n51912,
n51913, n51914, n51915, n51916, n51917, n51918, n51919, n51920,
n51921, n51922, n51923, n51924, n51925, n51926, n51927, n51928,
n51929, n51930, n51931, n51932, n51933, n51934, n51935, n51936,
n51937, n51938, n51939, n51940, n51941, n51942, n51943, n51944,
n51945, n51946, n51947, n51948, n51949, n51950, n51951, n51952,
n51953, n51954, n51955, n51956, n51957, n51958, n51959, n51960,
n51961, n51962, n51963, n51964, n51965, n51966, n51967, n51968,
n51969, n51970, n51971, n51972, n51973, n51974, n51975, n51976,
n51977, n51978, n51979, n51980, n51981, n51982, n51983, n51984,
n51985, n51986, n51987, n51988, n51989, n51990, n51991, n51992,
n51993, n51994, n51995, n51996, n51997, n51998, n51999, n52000,
n52001, n52002, n52003, n52004, n52005, n52006, n52007, n52008,
n52009, n52010, n52011, n52012, n52013, n52014, n52015, n52016,
n52017, n52018, n52019, n52020, n52021, n52022, n52023, n52024,
n52025, n52026, n52027, n52028, n52029, n52030, n52031, n52032,
n52033, n52034, n52035, n52036, n52037, n52038, n52039, n52040,
n52041, n52042, n52043, n52044, n52045, n52046, n52047, n52048,
n52049, n52050, n52051, n52052, n52053, n52054, n52055, n52056,
n52057, n52058, n52059, n52060, n52061, n52062, n52063, n52064,
n52065, n52066, n52067, n52068, n52069, n52070, n52071, n52072,
n52073, n52074, n52075, n52076, n52077, n52078, n52079, n52080,
n52081, n52082, n52083, n52084, n52085, n52086, n52087, n52088,
n52089, n52090, n52091, n52092, n52093, n52094, n52095, n52096,
n52097, n52098, n52099, n52100, n52101, n52102, n52103, n52104,
n52105, n52106, n52107, n52108, n52109, n52110, n52111, n52112,
n52113, n52114, n52115, n52116, n52117, n52118, n52119, n52120,
n52121, n52122, n52123, n52124, n52125, n52126, n52127, n52128,
n52129, n52130, n52131, n52132, n52133, n52134, n52135, n52136,
n52137, n52138, n52139, n52140, n52141, n52142, n52143, n52144,
n52145, n52146, n52147, n52148, n52149, n52150, n52151, n52152,
n52153, n52154, n52155, n52156, n52157, n52158, n52159, n52160,
n52161, n52162, n52163, n52164, n52165, n52166, n52167, n52168,
n52169, n52170, n52171, n52172, n52173, n52174, n52175, n52176,
n52177, n52178, n52179, n52180, n52181, n52182, n52183, n52184,
n52185, n52186, n52187, n52188, n52189, n52190, n52191, n52192,
n52193, n52194, n52195, n52196, n52197, n52198, n52199, n52200,
n52201, n52202, n52203, n52204, n52205, n52206, n52207, n52208,
n52209, n52210, n52211, n52212, n52213, n52214, n52215, n52216,
n52217, n52218, n52219, n52220, n52221, n52222, n52223, n52224,
n52225, n52226, n52227, n52228, n52229, n52230, n52231, n52232,
n52233, n52234, n52235, n52236, n52237, n52238, n52239, n52240,
n52241, n52242, n52243, n52244, n52245, n52246, n52247, n52248,
n52249, n52250, n52251, n52252, n52253, n52254, n52255, n52256,
n52257, n52258, n52259, n52260, n52261, n52262, n52263, n52264,
n52265, n52266, n52267, n52268, n52269, n52270, n52271, n52272,
n52273, n52274, n52275, n52276, n52277, n52278, n52279, n52280,
n52281, n52282, n52283, n52284, n52285, n52286, n52287, n52288,
n52289, n52290, n52291, n52292, n52293, n52294, n52295, n52296,
n52297, n52298, n52299, n52300, n52301, n52302, n52303, n52304,
n52305, n52306, n52307, n52308, n52309, n52310, n52311, n52312,
n52313, n52314, n52315, n52316, n52317, n52318, n52319, n52320,
n52321, n52322, n52323, n52324, n52325, n52326, n52327, n52328,
n52329, n52330, n52331, n52332, n52333, n52334, n52335, n52336,
n52337, n52338, n52339, n52340, n52341, n52342, n52343, n52344,
n52345, n52346, n52347, n52348, n52349, n52350, n52351, n52352,
n52353, n52354, n52355, n52356, n52357, n52358, n52359, n52360,
n52361, n52362, n52363, n52364, n52365, n52366, n52367, n52368,
n52369, n52370, n52371, n52372, n52373, n52374, n52375, n52376,
n52377, n52378, n52379, n52380, n52381, n52382, n52383, n52384,
n52385, n52386, n52387, n52388, n52389, n52390, n52391, n52392,
n52393, n52394, n52395, n52396, n52397, n52398, n52399, n52400,
n52401, n52402, n52403, n52404, n52405, n52406, n52407, n52408,
n52409, n52410, n52411, n52412, n52413, n52414, n52415, n52416,
n52417, n52418, n52419, n52420, n52421, n52422, n52423, n52424,
n52425, n52426, n52427, n52428, n52429, n52430, n52431, n52432,
n52433, n52434, n52435, n52436, n52437, n52438, n52439, n52440,
n52441, n52442, n52443, n52444, n52445, n52446, n52447, n52448,
n52449, n52450, n52451, n52452, n52453, n52454, n52455, n52456,
n52457, n52458, n52459, n52460, n52461, n52462, n52463, n52464,
n52465, n52466, n52467, n52468, n52469, n52470, n52471, n52472,
n52473, n52474, n52475, n52476, n52477, n52478, n52479, n52480,
n52481, n52482, n52483, n52484, n52485, n52486, n52487, n52488,
n52489, n52490, n52491, n52492, n52493, n52494, n52495, n52496,
n52497, n52498, n52499, n52500, n52501, n52502, n52503, n52504,
n52505, n52506, n52507, n52508, n52509, n52510, n52511, n52512,
n52513, n52514, n52515, n52516, n52517, n52518, n52519, n52520,
n52521, n52522, n52523, n52524, n52525, n52526, n52527, n52528,
n52529, n52530, n52531, n52532, n52533, n52534, n52535, n52536,
n52537, n52538, n52539, n52540, n52541, n52542, n52543, n52544,
n52545, n52546, n52547, n52548, n52549, n52550, n52551, n52552,
n52553, n52554, n52555, n52556, n52557, n52558, n52559, n52560,
n52561, n52562, n52563, n52564, n52565, n52566, n52567, n52568,
n52569, n52570, n52571, n52572, n52573, n52574, n52575, n52576,
n52577, n52578, n52579, n52580, n52581, n52582, n52583, n52584,
n52585, n52586, n52587, n52588, n52589, n52590, n52591, n52592,
n52593, n52594, n52595, n52596, n52597, n52598, n52599, n52600,
n52601, n52602, n52603, n52604, n52605, n52606, n52607, n52608,
n52609, n52610, n52611, n52612, n52613, n52614, n52615, n52616,
n52617, n52618, n52619, n52620, n52621, n52622, n52623, n52624,
n52625, n52626, n52627, n52628, n52629, n52630, n52631, n52632,
n52633, n52634, n52635, n52636, n52637, n52638, n52639, n52640,
n52641, n52642, n52643, n52644, n52645, n52646, n52647, n52648,
n52649, n52650, n52651, n52652, n52653, n52654, n52655, n52656,
n52657, n52658, n52659, n52660, n52661, n52662, n52663, n52664,
n52665, n52666, n52667, n52668, n52669, n52670, n52671, n52672,
n52673, n52674, n52675, n52676, n52677, n52678, n52679, n52680,
n52681, n52682, n52683, n52684, n52685, n52686, n52687, n52688,
n52689, n52690, n52691, n52692, n52693, n52694, n52695, n52696,
n52697, n52698, n52699, n52700, n52701, n52702, n52703, n52704,
n52705, n52706, n52707, n52708, n52709, n52710, n52711, n52712,
n52713, n52714, n52715, n52716, n52717, n52718, n52719, n52720,
n52721, n52722, n52723, n52724, n52725, n52726, n52727, n52728,
n52729, n52730, n52731, n52732, n52733, n52734, n52735, n52736,
n52737, n52738, n52739, n52740, n52741, n52742, n52743, n52744,
n52745, n52746, n52747, n52748, n52749, n52750, n52751, n52752,
n52753, n52754, n52755, n52756, n52757, n52758, n52759, n52760,
n52761, n52762, n52763, n52764, n52765, n52766, n52767, n52768,
n52769, n52770, n52771, n52772, n52773, n52774, n52775, n52776,
n52777, n52778, n52779, n52780, n52781, n52782, n52783, n52784,
n52785, n52786, n52787, n52788, n52789, n52790, n52791, n52792,
n52793, n52794, n52795, n52796, n52797, n52798, n52799, n52800,
n52801, n52802, n52803, n52804, n52805, n52806, n52807, n52808,
n52809, n52810, n52811, n52812, n52813, n52814, n52815, n52816,
n52817, n52818, n52819, n52820, n52821, n52822, n52823, n52824,
n52825, n52826, n52827, n52828, n52829, n52830, n52831, n52832,
n52833, n52834, n52835, n52836, n52837, n52838, n52839, n52840,
n52841, n52842, n52843, n52844, n52845, n52846, n52847, n52848,
n52849, n52850, n52851, n52852, n52853, n52854, n52855, n52856,
n52857, n52858, n52859, n52860, n52861, n52862, n52863, n52864,
n52865, n52866, n52867, n52868, n52869, n52870, n52871, n52872,
n52873, n52874, n52875, n52876, n52877, n52878, n52879, n52880,
n52881, n52882, n52883, n52884, n52885, n52886, n52887, n52888,
n52889, n52890, n52891, n52892, n52893, n52894, n52895, n52896,
n52897, n52898, n52899, n52900, n52901, n52902, n52903, n52904,
n52905, n52906, n52907, n52908, n52909, n52910, n52911, n52912,
n52913, n52914, n52915, n52916, n52917, n52918, n52919, n52920,
n52921, n52922, n52923, n52924, n52925, n52926, n52927, n52928,
n52929, n52930, n52931, n52932, n52933, n52934, n52935, n52936,
n52937, n52938, n52939, n52940, n52941, n52942, n52943, n52944,
n52945, n52946, n52947, n52948, n52949, n52950, n52951, n52952,
n52953, n52954, n52955, n52956, n52957, n52958, n52959, n52960,
n52961, n52962, n52963, n52964, n52965, n52966, n52967, n52968,
n52969, n52970, n52971, n52972, n52973, n52974, n52975, n52976,
n52977, n52978, n52979, n52980, n52981, n52982, n52983, n52984,
n52985, n52986, n52987, n52988, n52989, n52990, n52991, n52992,
n52993, n52994, n52995, n52996, n52997, n52998, n52999, n53000,
n53001, n53002, n53003, n53004, n53005, n53006, n53007, n53008,
n53009, n53010, n53011, n53012, n53013, n53014, n53015, n53016,
n53017, n53018, n53019, n53020, n53021, n53022, n53023, n53024,
n53025, n53026, n53027, n53028, n53029, n53030, n53031, n53032,
n53033, n53034, n53035, n53036, n53037, n53038, n53039, n53040,
n53041, n53042, n53043, n53044, n53045, n53046, n53047, n53048,
n53049, n53050, n53051, n53052, n53053, n53054, n53055, n53056,
n53057, n53058, n53059, n53060, n53061, n53062, n53063, n53064,
n53065, n53066, n53067, n53068, n53069, n53070, n53071, n53072,
n53073, n53074, n53075, n53076, n53077, n53078, n53079, n53080,
n53081, n53082, n53083, n53084, n53085, n53086, n53087, n53088,
n53089, n53090, n53091, n53092, n53093, n53094, n53095, n53096,
n53097, n53098, n53099, n53100, n53101, n53102, n53103, n53104,
n53105, n53106, n53107, n53108, n53109, n53110, n53111, n53112,
n53113;


   and U26626 ( n25181,n28132,n28738 );
   and U26627 ( n25182,n28094,n49328 );
   and U26628 ( n25183,n41032,n27896 );
   and U26629 ( n25184,n41847,n41848 );
   not U26630 ( p2_u2874,n25184 );
   and U26631 ( n25186,n41802,n41803 );
   not U26632 ( p2_u2880,n25186 );
   nand U26633 ( n25188,p1_instqueuewr_addr_reg_4_,n45384 );
   not U26634 ( p1_u3032,n25188 );
   nand U26635 ( n25190,p2_instqueuewr_addr_reg_4_,n36665 );
   not U26636 ( p2_u3047,n25190 );
   and U26637 ( n25192,n34231,n34232 );
   not U26638 ( p3_u2703,n25192 );
   and U26639 ( n25194,n41816,n41817 );
   not U26640 ( p2_u2878,n25194 );
   and U26641 ( n25196,n41772,n41773 );
   not U26642 ( p2_u2885,n25196 );
   and U26643 ( n25198,n41833,n41834 );
   not U26644 ( p2_u2876,n25198 );
   and U26645 ( n25200,n41866,n41867 );
   not U26646 ( p2_u2872,n25200 );
   and U26647 ( n25202,n41782,n41783 );
   not U26648 ( p2_u2883,n25202 );
   and U26649 ( n25204,n34389,n34390 );
   not U26650 ( p3_u2693,n25204 );
   and U26651 ( n25206,n34543,n34544 );
   not U26652 ( p3_u2689,n25206 );
   and U26653 ( n25208,n34633,n34634 );
   not U26654 ( p3_u2687,n25208 );
   and U26655 ( n25210,n34279,n34280 );
   not U26656 ( p3_u2697,n25210 );
   and U26657 ( n25212,n34246,n34247 );
   not U26658 ( p3_u2701,n25212 );
   and U26659 ( n25214,n34262,n34263 );
   not U26660 ( p3_u2699,n25214 );
   and U26661 ( n25216,n41875,n41876 );
   not U26662 ( p2_u2871,n25216 );
   and U26663 ( n25218,n41840,n41841 );
   not U26664 ( p2_u2875,n25218 );
   and U26665 ( n25220,n41794,n41795 );
   not U26666 ( p2_u2881,n25220 );
   and U26667 ( n25222,n41759,n41760 );
   not U26668 ( p2_u2887,n25222 );
   and U26669 ( n25224,n34296,n34297 );
   not U26670 ( p3_u2695,n25224 );
   and U26671 ( n25226,n41777,n41778 );
   not U26672 ( p2_u2884,n25226 );
   and U26673 ( n25228,n34990,n34991 );
   not U26674 ( p3_u2674,n25228 );
   and U26675 ( n25230,n34999,n35000 );
   not U26676 ( p3_u2673,n25230 );
   and U26677 ( n25232,n41767,n41768 );
   not U26678 ( p2_u2886,n25232 );
   and U26679 ( n25234,n41809,n41810 );
   not U26680 ( p2_u2879,n25234 );
   and U26681 ( n25236,n41858,n41859 );
   not U26682 ( p2_u2873,n25236 );
   and U26683 ( n25238,n41826,n41827 );
   not U26684 ( p2_u2877,n25238 );
   and U26685 ( n25240,n34272,n34273 );
   not U26686 ( p3_u2698,n25240 );
   and U26687 ( n25242,n34255,n34256 );
   not U26688 ( p3_u2700,n25242 );
   and U26689 ( n25244,n34352,n34353 );
   not U26690 ( p3_u2694,n25244 );
   and U26691 ( n25246,n34289,n34290 );
   not U26692 ( p3_u2696,n25246 );
   and U26693 ( n25248,n34429,n34430 );
   not U26694 ( p3_u2692,n25248 );
   and U26695 ( n25250,n34583,n34584 );
   not U26696 ( p3_u2688,n25250 );
   and U26697 ( n25252,n49044,n49045 );
   not U26698 ( p1_u2963,n25252 );
   and U26699 ( n25254,n49054,n49055 );
   not U26700 ( p1_u2961,n25254 );
   and U26701 ( n25256,n49039,n49040 );
   not U26702 ( p1_u2964,n25256 );
   and U26703 ( n25258,n49049,n49050 );
   not U26704 ( p1_u2962,n25258 );
   and U26705 ( n25260,n28893,n28894 );
   not U26706 ( p3_u3281,n25260 );
   and U26707 ( n25262,n45504,n45505 );
   not U26708 ( p1_u3465,n25262 );
   and U26709 ( n25264,n49029,n49030 );
   not U26710 ( p1_u2966,n25264 );
   and U26711 ( n25266,n49079,n49080 );
   not U26712 ( p1_u2956,n25266 );
   and U26713 ( n25268,n49104,n49105 );
   not U26714 ( p1_u2951,n25268 );
   and U26715 ( n25270,n49094,n49095 );
   not U26716 ( p1_u2953,n25270 );
   and U26717 ( n25272,n49089,n49090 );
   not U26718 ( p1_u2954,n25272 );
   and U26719 ( n25274,n49069,n49070 );
   not U26720 ( p1_u2958,n25274 );
   and U26721 ( n25276,n49099,n49100 );
   not U26722 ( p1_u2952,n25276 );
   and U26723 ( n25278,n49074,n49075 );
   not U26724 ( p1_u2957,n25278 );
   and U26725 ( n25280,n49059,n49060 );
   not U26726 ( p1_u2960,n25280 );
   and U26727 ( n25282,n49084,n49085 );
   not U26728 ( p1_u2955,n25282 );
   and U26729 ( n25284,n49034,n49035 );
   not U26730 ( p1_u2965,n25284 );
   and U26731 ( n25286,n49064,n49065 );
   not U26732 ( p1_u2959,n25286 );
   and U26733 ( n25288,n49352,n49353 );
   not U26734 ( p1_u2901,n25288 );
   and U26735 ( n25290,n49400,n49401 );
   not U26736 ( p1_u2893,n25290 );
   and U26737 ( n25292,n49376,n49377 );
   not U26738 ( p1_u2897,n25292 );
   and U26739 ( n25294,n49370,n49371 );
   not U26740 ( p1_u2898,n25294 );
   and U26741 ( n25296,n33399,n33400 );
   not U26742 ( p3_u2737,n25296 );
   and U26743 ( n25298,n28749,n27891 );
   not U26744 ( u212,n25298 );
   and U26745 ( n25300,n49424,n49425 );
   not U26746 ( p1_u2889,n25300 );
   and U26747 ( n25302,n49394,n49395 );
   not U26748 ( p1_u2894,n25302 );
   and U26749 ( n25304,n49333,n49334 );
   not U26750 ( p1_u2904,n25304 );
   and U26751 ( n25306,n49388,n49389 );
   not U26752 ( p1_u2895,n25306 );
   and U26753 ( n25308,n49418,n49419 );
   not U26754 ( p1_u2890,n25308 );
   and U26755 ( n25310,n49358,n49359 );
   not U26756 ( p1_u2900,n25310 );
   and U26757 ( n25312,n49318,n49319 );
   not U26758 ( p1_u2907,n25312 );
   and U26759 ( n25314,n49263,n49264 );
   not U26760 ( p1_u2918,n25314 );
   and U26761 ( n25316,n49288,n49289 );
   not U26762 ( p1_u2913,n25316 );
   and U26763 ( n25318,n49181,n49182 );
   not U26764 ( p1_u2935,n25318 );
   and U26765 ( n25320,n49278,n49279 );
   not U26766 ( p1_u2915,n25320 );
   and U26767 ( n25322,n49293,n49294 );
   not U26768 ( p1_u2912,n25322 );
   and U26769 ( n25324,n49268,n49269 );
   not U26770 ( p1_u2917,n25324 );
   and U26771 ( n25326,n49308,n49309 );
   not U26772 ( p1_u2909,n25326 );
   and U26773 ( n25328,n49273,n49274 );
   not U26774 ( p1_u2916,n25328 );
   and U26775 ( n25330,n49174,n49175 );
   not U26776 ( p1_u2936,n25330 );
   and U26777 ( n25332,n49313,n49314 );
   not U26778 ( p1_u2908,n25332 );
   and U26779 ( n25334,n49258,n49259 );
   not U26780 ( p1_u2919,n25334 );
   and U26781 ( n25336,n41061,n41062 );
   not U26782 ( p2_u2947,n25336 );
   and U26783 ( n25338,n49303,n49304 );
   not U26784 ( p1_u2910,n25338 );
   and U26785 ( n25340,n49298,n49299 );
   not U26786 ( p1_u2911,n25340 );
   and U26787 ( n25342,n49283,n49284 );
   not U26788 ( p1_u2914,n25342 );
   and U26789 ( n25344,n49252,n49253 );
   not U26790 ( p1_u2920,n25344 );
   and U26791 ( n25346,n49323,n49324 );
   not U26792 ( p1_u2906,n25346 );
   and U26793 ( n25348,n41056,n41057 );
   not U26794 ( p2_u2948,n25348 );
   and U26795 ( n25350,n41051,n41052 );
   not U26796 ( p2_u2949,n25350 );
   and U26797 ( n25352,n41066,n41067 );
   not U26798 ( p2_u2946,n25352 );
   and U26799 ( n25354,n41076,n41077 );
   not U26800 ( p2_u2944,n25354 );
   and U26801 ( n25356,n41111,n41112 );
   not U26802 ( p2_u2937,n25356 );
   and U26803 ( n25358,n41046,n41047 );
   not U26804 ( p2_u2950,n25358 );
   and U26805 ( n25360,n41116,n41117 );
   not U26806 ( p2_u2936,n25360 );
   and U26807 ( n25362,n41071,n41072 );
   not U26808 ( p2_u2945,n25362 );
   and U26809 ( n25364,n41122,n41123 );
   not U26810 ( p2_u2935,n25364 );
   and U26811 ( n25366,n41106,n41107 );
   not U26812 ( p2_u2938,n25366 );
   and U26813 ( n25368,n41096,n41097 );
   not U26814 ( p2_u2940,n25368 );
   and U26815 ( n25370,n41101,n41102 );
   not U26816 ( p2_u2939,n25370 );
   and U26817 ( n25372,n30779,n30780 );
   not U26818 ( p3_u2864,n25372 );
   and U26819 ( n25374,n36313,n36314 );
   not U26820 ( p3_u2636,n25374 );
   and U26821 ( n25376,n36317,n36314 );
   not U26822 ( p3_u2635,n25376 );
   and U26823 ( n25378,n41091,n41092 );
   not U26824 ( p2_u2941,n25378 );
   and U26825 ( n25380,n41081,n41082 );
   not U26826 ( p2_u2943,n25380 );
   and U26827 ( n25382,n41086,n41087 );
   not U26828 ( p2_u2942,n25382 );
   and U26829 ( n25384,n49205,n49206 );
   not U26830 ( p1_u2930,n25384 );
   and U26831 ( n25386,n49234,n49235 );
   not U26832 ( p1_u2924,n25386 );
   and U26833 ( n25388,n49225,n49226 );
   not U26834 ( p1_u2926,n25388 );
   and U26835 ( n25390,n49229,n49230 );
   not U26836 ( p1_u2925,n25390 );
   and U26837 ( n25392,n49186,n49187 );
   not U26838 ( p1_u2934,n25392 );
   and U26839 ( n25394,n34199,n34200 );
   not U26840 ( p3_u2704,n25394 );
   and U26841 ( n25396,n49248,n49249 );
   not U26842 ( p1_u2921,n25396 );
   and U26843 ( n25398,n49191,n49192 );
   not U26844 ( p1_u2933,n25398 );
   and U26845 ( n25400,n49201,n49202 );
   not U26846 ( p1_u2931,n25400 );
   and U26847 ( n25402,n49196,n49197 );
   not U26848 ( p1_u2932,n25402 );
   and U26849 ( n25404,n49244,n49245 );
   not U26850 ( p1_u2922,n25404 );
   and U26851 ( n25406,n49239,n49240 );
   not U26852 ( p1_u2923,n25406 );
   and U26853 ( n25408,n41929,n41930 );
   not U26854 ( p2_u2864,n25408 );
   and U26855 ( n25410,n41899,n41900 );
   not U26856 ( p2_u2868,n25410 );
   and U26857 ( n25412,n41914,n41915 );
   not U26858 ( p2_u2866,n25412 );
   and U26859 ( n25414,n49210,n49211 );
   not U26860 ( p1_u2929,n25414 );
   and U26861 ( n25416,n49215,n49216 );
   not U26862 ( p1_u2928,n25416 );
   and U26863 ( n25418,n49220,n49221 );
   not U26864 ( p1_u2927,n25418 );
   and U26865 ( n25420,n49109,n49110 );
   not U26866 ( p1_u2950,n25420 );
   and U26867 ( n25422,n49155,n49156 );
   not U26868 ( p1_u2940,n25422 );
   and U26869 ( n25424,n49143,n49144 );
   not U26870 ( p1_u2943,n25424 );
   and U26871 ( n25426,n49119,n49120 );
   not U26872 ( p1_u2948,n25426 );
   and U26873 ( n25428,n49021,n49022 );
   not U26874 ( p1_u2967,n25428 );
   and U26875 ( n25430,n49114,n49115 );
   not U26876 ( p1_u2949,n25430 );
   and U26877 ( n25432,n49163,n49164 );
   not U26878 ( p1_u2938,n25432 );
   and U26879 ( n25434,n49147,n49148 );
   not U26880 ( p1_u2942,n25434 );
   and U26881 ( n25436,n49151,n49152 );
   not U26882 ( p1_u2941,n25436 );
   and U26883 ( n25438,n49124,n49125 );
   not U26884 ( p1_u2947,n25438 );
   and U26885 ( n25440,n49134,n49135 );
   not U26886 ( p1_u2945,n25440 );
   and U26887 ( n25442,n49139,n49140 );
   not U26888 ( p1_u2944,n25442 );
   and U26889 ( n25444,n41163,n41164 );
   not U26890 ( p2_u2927,n25444 );
   and U26891 ( n25446,n41148,n41149 );
   not U26892 ( p2_u2930,n25446 );
   and U26893 ( n25448,n49821,n49822 );
   not U26894 ( p1_u2841,n25448 );
   and U26895 ( n25450,n49159,n49160 );
   not U26896 ( p1_u2939,n25450 );
   and U26897 ( n25452,n49167,n49168 );
   not U26898 ( p1_u2937,n25452 );
   and U26899 ( n25454,n49129,n49130 );
   not U26900 ( p1_u2946,n25454 );
   and U26901 ( n25456,n41138,n41139 );
   not U26902 ( p2_u2932,n25456 );
   and U26903 ( n25458,n41128,n41129 );
   not U26904 ( p2_u2934,n25458 );
   and U26905 ( n25460,n41133,n41134 );
   not U26906 ( p2_u2933,n25460 );
   and U26907 ( n25462,n41168,n41169 );
   not U26908 ( p2_u2926,n25462 );
   and U26909 ( n25464,n41038,n41039 );
   not U26910 ( p2_u2951,n25464 );
   and U26911 ( n25466,n41153,n41154 );
   not U26912 ( p2_u2929,n25466 );
   and U26913 ( n25468,n41158,n41159 );
   not U26914 ( p2_u2928,n25468 );
   and U26915 ( n25470,n41193,n41194 );
   not U26916 ( p2_u2921,n25470 );
   and U26917 ( n25472,n41173,n41174 );
   not U26918 ( p2_u2925,n25472 );
   and U26919 ( n25474,n41178,n41179 );
   not U26920 ( p2_u2924,n25474 );
   and U26921 ( n25476,n41188,n41189 );
   not U26922 ( p2_u2922,n25476 );
   and U26923 ( n25478,n41143,n41144 );
   not U26924 ( p2_u2931,n25478 );
   and U26925 ( n25480,n41999,n42000 );
   not U26926 ( p2_u2858,n25480 );
   and U26927 ( n25482,n41920,n41921 );
   not U26928 ( p2_u2865,n25482 );
   and U26929 ( n25484,n41940,n41941 );
   not U26930 ( p2_u2863,n25484 );
   and U26931 ( n25486,n42006,n42007 );
   not U26932 ( p2_u2857,n25486 );
   and U26933 ( n25488,n41884,n41885 );
   not U26934 ( p2_u2870,n25488 );
   and U26935 ( n25490,n41183,n41184 );
   not U26936 ( p2_u2923,n25490 );
   and U26937 ( n25492,n41987,n41988 );
   not U26938 ( p2_u2859,n25492 );
   and U26939 ( n25494,n41976,n41977 );
   not U26940 ( p2_u2860,n25494 );
   and U26941 ( n25496,n41964,n41965 );
   not U26942 ( p2_u2861,n25496 );
   and U26943 ( n25498,n41890,n41891 );
   not U26944 ( p2_u2869,n25498 );
   and U26945 ( n25500,n41905,n41906 );
   not U26946 ( p2_u2867,n25500 );
   and U26947 ( n25502,n41953,n41954 );
   not U26948 ( p2_u2862,n25502 );
   and U26949 ( n25504,n34880,n34881 );
   not U26950 ( p3_u2681,n25504 );
   and U26951 ( n25506,n34803,n34804 );
   not U26952 ( p3_u2683,n25506 );
   and U26953 ( n25508,n34466,n34467 );
   not U26954 ( p3_u2691,n25508 );
   and U26955 ( n25510,n34929,n34930 );
   not U26956 ( p3_u2679,n25510 );
   and U26957 ( n25512,n34920,n34921 );
   not U26958 ( p3_u2680,n25512 );
   and U26959 ( n25514,n36980,n36981 );
   not U26960 ( p2_u3210,n25514 );
   and U26961 ( n25516,n34843,n34844 );
   not U26962 ( p3_u2682,n25516 );
   and U26963 ( n25518,n34766,n34767 );
   not U26964 ( p3_u2684,n25518 );
   and U26965 ( n25520,n34978,n34979 );
   not U26966 ( p3_u2675,n25520 );
   and U26967 ( n25522,n34506,n34507 );
   not U26968 ( p3_u2690,n25522 );
   and U26969 ( n25524,n34955,n34956 );
   not U26970 ( p3_u2677,n25524 );
   and U26971 ( n25526,n34689,n34690 );
   not U26972 ( p3_u2686,n25526 );
   and U26973 ( n25528,n28427,n28428 );
   not U26974 ( u369,n25528 );
   and U26975 ( n25530,n28433,n28434 );
   not U26976 ( u366,n25530 );
   and U26977 ( n25532,n28455,n28456 );
   not U26978 ( u355,n25532 );
   and U26979 ( n25534,n28447,n28448 );
   not U26980 ( u359,n25534 );
   and U26981 ( n25536,n28421,n28422 );
   not U26982 ( u372,n25536 );
   and U26983 ( n25538,n34726,n34727 );
   not U26984 ( p3_u2685,n25538 );
   and U26985 ( n25540,n28423,n28424 );
   not U26986 ( u371,n25540 );
   and U26987 ( n25542,n28429,n28430 );
   not U26988 ( u368,n25542 );
   and U26989 ( n25544,n28435,n28436 );
   not U26990 ( u365,n25544 );
   and U26991 ( n25546,n28425,n28426 );
   not U26992 ( u370,n25546 );
   and U26993 ( n25548,n28439,n28440 );
   not U26994 ( u363,n25548 );
   and U26995 ( n25550,n28417,n28418 );
   not U26996 ( u374,n25550 );
   and U26997 ( n25552,n28437,n28438 );
   not U26998 ( u364,n25552 );
   and U26999 ( n25554,n28449,n28450 );
   not U27000 ( u358,n25554 );
   and U27001 ( n25556,n28445,n28446 );
   not U27002 ( u360,n25556 );
   and U27003 ( n25558,n28443,n28444 );
   not U27004 ( u361,n25558 );
   and U27005 ( n25560,n28453,n28454 );
   not U27006 ( u356,n25560 );
   and U27007 ( n25562,n28419,n28420 );
   not U27008 ( u373,n25562 );
   and U27009 ( n25564,n52744,n52741 );
   not U27010 ( p1_u2804,n25564 );
   and U27011 ( n25566,n42616,n42617 );
   not U27012 ( p2_u2856,n25566 );
   and U27013 ( n25568,n28431,n28432 );
   not U27014 ( u367,n25568 );
   and U27015 ( n25570,n28451,n28452 );
   not U27016 ( u357,n25570 );
   and U27017 ( n25572,n28457,n28458 );
   not U27018 ( u354,n25572 );
   and U27019 ( n25574,n28441,n28442 );
   not U27020 ( u362,n25574 );
   and U27021 ( n25576,n49732,n49733 );
   not U27022 ( p1_u2857,n25576 );
   and U27023 ( n25578,n49701,n49702 );
   not U27024 ( p1_u2864,n25578 );
   and U27025 ( n25580,n49710,n49711 );
   not U27026 ( p1_u2862,n25580 );
   and U27027 ( n25582,n52740,n52741 );
   not U27028 ( p1_u2805,n25582 );
   and U27029 ( n25584,n44721,n44722 );
   not U27030 ( p2_u2818,n25584 );
   and U27031 ( n25586,n44725,n44722 );
   not U27032 ( p2_u2817,n25586 );
   and U27033 ( n25588,n49728,n49729 );
   not U27034 ( p1_u2858,n25588 );
   and U27035 ( n25590,n49696,n49697 );
   not U27036 ( p1_u2865,n25590 );
   and U27037 ( n25592,n49737,n49738 );
   not U27038 ( p1_u2856,n25592 );
   and U27039 ( n25594,n49742,n49743 );
   not U27040 ( p1_u2855,n25594 );
   and U27041 ( n25596,n49673,n49674 );
   not U27042 ( p1_u2870,n25596 );
   and U27043 ( n25598,n49714,n49715 );
   not U27044 ( p1_u2861,n25598 );
   and U27045 ( n25600,n49723,n49724 );
   not U27046 ( p1_u2859,n25600 );
   and U27047 ( n25602,n49687,n49688 );
   not U27048 ( p1_u2867,n25602 );
   and U27049 ( n25604,n49683,n49684 );
   not U27050 ( p1_u2868,n25604 );
   and U27051 ( n25606,n49705,n49706 );
   not U27052 ( p1_u2863,n25606 );
   and U27053 ( n25608,n49692,n49693 );
   not U27054 ( p1_u2866,n25608 );
   and U27055 ( n25610,n49719,n49720 );
   not U27056 ( p1_u2860,n25610 );
   and U27057 ( n25612,n33284,n33285 );
   not U27058 ( p3_u2760,n25612 );
   and U27059 ( n25614,n33294,n33295 );
   not U27060 ( p3_u2758,n25614 );
   and U27061 ( n25616,n33299,n33300 );
   not U27062 ( p3_u2757,n25616 );
   and U27063 ( n25618,n33269,n33270 );
   not U27064 ( p3_u2763,n25618 );
   and U27065 ( n25620,n45510,n45511 );
   not U27066 ( p1_u3464,n25620 );
   and U27067 ( n25622,n28900,n28901 );
   not U27068 ( p3_u3280,n25622 );
   and U27069 ( n25624,n33289,n33290 );
   not U27070 ( p3_u2759,n25624 );
   and U27071 ( n25626,n33314,n33315 );
   not U27072 ( p3_u2754,n25626 );
   and U27073 ( n25628,n33279,n33280 );
   not U27074 ( p3_u2761,n25628 );
   and U27075 ( n25630,n33349,n33350 );
   not U27076 ( p3_u2747,n25630 );
   and U27077 ( n25632,n33324,n33325 );
   not U27078 ( p3_u2752,n25632 );
   and U27079 ( n25634,n33359,n33360 );
   not U27080 ( p3_u2745,n25634 );
   and U27081 ( n25636,n33344,n33345 );
   not U27082 ( p3_u2748,n25636 );
   and U27083 ( n25638,n33259,n33260 );
   not U27084 ( p3_u2765,n25638 );
   and U27085 ( n25640,n33334,n33335 );
   not U27086 ( p3_u2750,n25640 );
   and U27087 ( n25642,n33319,n33320 );
   not U27088 ( p3_u2753,n25642 );
   and U27089 ( n25644,n33364,n33365 );
   not U27090 ( p3_u2744,n25644 );
   and U27091 ( n25646,n33304,n33305 );
   not U27092 ( p3_u2756,n25646 );
   and U27093 ( n25648,n33264,n33265 );
   not U27094 ( p3_u2764,n25648 );
   and U27095 ( n25650,n33274,n33275 );
   not U27096 ( p3_u2762,n25650 );
   and U27097 ( n25652,n33329,n33330 );
   not U27098 ( p3_u2751,n25652 );
   and U27099 ( n25654,n33309,n33310 );
   not U27100 ( p3_u2755,n25654 );
   and U27101 ( n25656,n33339,n33340 );
   not U27102 ( p3_u2749,n25656 );
   and U27103 ( n25658,n33354,n33355 );
   not U27104 ( p3_u2746,n25658 );
   and U27105 ( n25660,n36871,n36872 );
   not U27106 ( p2_u3229,n25660 );
   and U27107 ( n25662,n36881,n36882 );
   not U27108 ( p2_u3227,n25662 );
   and U27109 ( n25664,n36876,n36877 );
   not U27110 ( p2_u3228,n25664 );
   and U27111 ( n25666,n36931,n36932 );
   not U27112 ( p2_u3217,n25666 );
   and U27113 ( n25668,n36886,n36887 );
   not U27114 ( p2_u3226,n25668 );
   and U27115 ( n25670,n29010,n29011 );
   not U27116 ( p3_u3042,n25670 );
   and U27117 ( n25672,n29005,n29006 );
   not U27118 ( p3_u3043,n25672 );
   and U27119 ( n25674,n28950,n28951 );
   not U27120 ( p3_u3054,n25674 );
   and U27121 ( n25676,n28975,n28976 );
   not U27122 ( p3_u3049,n25676 );
   and U27123 ( n25678,n36846,n36847 );
   not U27124 ( p2_u3234,n25678 );
   and U27125 ( n25680,n36861,n36862 );
   not U27126 ( p2_u3231,n25680 );
   and U27127 ( n25682,n36851,n36852 );
   not U27128 ( p2_u3233,n25682 );
   and U27129 ( n25684,n36906,n36907 );
   not U27130 ( p2_u3222,n25684 );
   and U27131 ( n25686,n28930,n28931 );
   not U27132 ( p3_u3058,n25686 );
   and U27133 ( n25688,n36921,n36922 );
   not U27134 ( p2_u3219,n25688 );
   and U27135 ( n25690,n28965,n28966 );
   not U27136 ( p3_u3051,n25690 );
   and U27137 ( n25692,n36901,n36902 );
   not U27138 ( p2_u3223,n25692 );
   and U27139 ( n25694,n36826,n36827 );
   not U27140 ( p2_u3238,n25694 );
   and U27141 ( n25696,n36816,n36817 );
   not U27142 ( p2_u3240,n25696 );
   and U27143 ( n25698,n28910,n28911 );
   not U27144 ( p3_u3274,n25698 );
   and U27145 ( n25700,n36804,n36805 );
   not U27146 ( p2_u3586,n25700 );
   and U27147 ( n25702,n28980,n28981 );
   not U27148 ( p3_u3048,n25702 );
   and U27149 ( n25704,n36831,n36832 );
   not U27150 ( p2_u3237,n25704 );
   and U27151 ( n25706,n36836,n36837 );
   not U27152 ( p2_u3236,n25706 );
   and U27153 ( n25708,n45595,n45596 );
   not U27154 ( p1_u3212,n25708 );
   and U27155 ( n25710,n45645,n45646 );
   not U27156 ( p1_u3202,n25710 );
   and U27157 ( n25712,n45522,n45523 );
   not U27158 ( p1_u3226,n25712 );
   and U27159 ( n25714,n45330,n45331 );
   not U27160 ( p1_u3486,n25714 );
   and U27161 ( n25716,n45605,n45606 );
   not U27162 ( p1_u3210,n25716 );
   and U27163 ( n25718,n28908,n28909 );
   not U27164 ( p3_u3275,n25718 );
   and U27165 ( n25720,n36951,n36952 );
   not U27166 ( p2_u3213,n25720 );
   and U27167 ( n25722,n45620,n45621 );
   not U27168 ( p1_u3207,n25722 );
   and U27169 ( n25724,n29055,n29056 );
   not U27170 ( p3_u3033,n25724 );
   and U27171 ( n25726,n28778,n28779 );
   not U27172 ( p3_u3297,n25726 );
   and U27173 ( n25728,n36806,n36807 );
   not U27174 ( p2_u3585,n25728 );
   and U27175 ( n25730,n29035,n29036 );
   not U27176 ( p3_u3037,n25730 );
   and U27177 ( n25732,n45530,n45531 );
   not U27178 ( p1_u3225,n25732 );
   and U27179 ( n25734,n45518,n45519 );
   not U27180 ( p1_u3459,n25734 );
   and U27181 ( n25736,n45565,n45566 );
   not U27182 ( p1_u3218,n25736 );
   and U27183 ( n25738,n45635,n45636 );
   not U27184 ( p1_u3204,n25738 );
   and U27185 ( n25740,n45665,n45666 );
   not U27186 ( p1_u3198,n25740 );
   and U27187 ( n25742,n29025,n29026 );
   not U27188 ( p3_u3039,n25742 );
   and U27189 ( n25744,n28945,n28946 );
   not U27190 ( p3_u3055,n25744 );
   and U27191 ( n25746,n45615,n45616 );
   not U27192 ( p1_u3208,n25746 );
   and U27193 ( n25748,n28920,n28921 );
   not U27194 ( p3_u3060,n25748 );
   and U27195 ( n25750,n28990,n28991 );
   not U27196 ( p3_u3046,n25750 );
   and U27197 ( n25752,n28912,n28913 );
   not U27198 ( p3_u3061,n25752 );
   and U27199 ( n25754,n28935,n28936 );
   not U27200 ( p3_u3057,n25754 );
   and U27201 ( n25756,n45585,n45586 );
   not U27202 ( p1_u3214,n25756 );
   and U27203 ( n25758,n45600,n45601 );
   not U27204 ( p1_u3211,n25758 );
   and U27205 ( n25760,n45540,n45541 );
   not U27206 ( p1_u3223,n25760 );
   and U27207 ( n25762,n36617,n36618 );
   not U27208 ( p2_u3611,n25762 );
   and U27209 ( n25764,n45560,n45561 );
   not U27210 ( p1_u3219,n25764 );
   and U27211 ( n25766,n28955,n28956 );
   not U27212 ( p3_u3053,n25766 );
   and U27213 ( n25768,n28995,n28996 );
   not U27214 ( p3_u3045,n25768 );
   and U27215 ( n25770,n45550,n45551 );
   not U27216 ( p1_u3221,n25770 );
   and U27217 ( n25772,n36808,n36809 );
   not U27218 ( p2_u3241,n25772 );
   and U27219 ( n25774,n36841,n36842 );
   not U27220 ( p2_u3235,n25774 );
   and U27221 ( n25776,n28940,n28941 );
   not U27222 ( p3_u3056,n25776 );
   and U27223 ( n25778,n28985,n28986 );
   not U27224 ( p3_u3047,n25778 );
   and U27225 ( n25780,n45520,n45521 );
   not U27226 ( p1_u3458,n25780 );
   and U27227 ( n25782,n45555,n45556 );
   not U27228 ( p1_u3220,n25782 );
   and U27229 ( n25784,n45545,n45546 );
   not U27230 ( p1_u3222,n25784 );
   and U27231 ( n25786,n45575,n45576 );
   not U27232 ( p1_u3216,n25786 );
   and U27233 ( n25788,n45590,n45591 );
   not U27234 ( p1_u3213,n25788 );
   and U27235 ( n25790,n36891,n36892 );
   not U27236 ( p2_u3225,n25790 );
   and U27237 ( n25792,n36941,n36942 );
   not U27238 ( p2_u3215,n25792 );
   and U27239 ( n25794,n36936,n36937 );
   not U27240 ( p2_u3216,n25794 );
   and U27241 ( n25796,n36916,n36917 );
   not U27242 ( p2_u3220,n25796 );
   and U27243 ( n25798,n29045,n29046 );
   not U27244 ( p3_u3035,n25798 );
   and U27245 ( n25800,n36946,n36947 );
   not U27246 ( p2_u3214,n25800 );
   and U27247 ( n25802,n28970,n28971 );
   not U27248 ( p3_u3050,n25802 );
   and U27249 ( n25804,n29020,n29021 );
   not U27250 ( p3_u3040,n25804 );
   and U27251 ( n25806,n36896,n36897 );
   not U27252 ( p2_u3224,n25806 );
   and U27253 ( n25808,n29060,n29061 );
   not U27254 ( p3_u3032,n25808 );
   and U27255 ( n25810,n29030,n29031 );
   not U27256 ( p3_u3038,n25810 );
   and U27257 ( n25812,n29050,n29051 );
   not U27258 ( p3_u3034,n25812 );
   and U27259 ( n25814,n36956,n36957 );
   not U27260 ( p2_u3212,n25814 );
   and U27261 ( n25816,n29015,n29016 );
   not U27262 ( p3_u3041,n25816 );
   and U27263 ( n25818,n28960,n28961 );
   not U27264 ( p3_u3052,n25818 );
   and U27265 ( n25820,n29000,n29001 );
   not U27266 ( p3_u3044,n25820 );
   and U27267 ( n25822,n36856,n36857 );
   not U27268 ( p2_u3232,n25822 );
   and U27269 ( n25824,n36911,n36912 );
   not U27270 ( p2_u3221,n25824 );
   and U27271 ( n25826,n45660,n45661 );
   not U27272 ( p1_u3199,n25826 );
   and U27273 ( n25828,n45535,n45536 );
   not U27274 ( p1_u3224,n25828 );
   and U27275 ( n25830,n36821,n36822 );
   not U27276 ( p2_u3239,n25830 );
   and U27277 ( n25832,n45516,n45517 );
   not U27278 ( p1_u3460,n25832 );
   and U27279 ( n25834,n45630,n45631 );
   not U27280 ( p1_u3205,n25834 );
   and U27281 ( n25836,n45570,n45571 );
   not U27282 ( p1_u3217,n25836 );
   and U27283 ( n25838,n45650,n45651 );
   not U27284 ( p1_u3201,n25838 );
   and U27285 ( n25840,n36802,n36803 );
   not U27286 ( p2_u3587,n25840 );
   and U27287 ( n25842,n36800,n36801 );
   not U27288 ( p2_u3588,n25842 );
   and U27289 ( n25844,n28925,n28926 );
   not U27290 ( p3_u3059,n25844 );
   and U27291 ( n25846,n28906,n28907 );
   not U27292 ( p3_u3276,n25846 );
   and U27293 ( n25848,n36866,n36867 );
   not U27294 ( p2_u3230,n25848 );
   and U27295 ( n25850,n45514,n45515 );
   not U27296 ( p1_u3461,n25850 );
   and U27297 ( n25852,n45655,n45656 );
   not U27298 ( p1_u3200,n25852 );
   and U27299 ( n25854,n29040,n29041 );
   not U27300 ( p3_u3036,n25854 );
   and U27301 ( n25856,n45610,n45611 );
   not U27302 ( p1_u3209,n25856 );
   and U27303 ( n25858,n45640,n45641 );
   not U27304 ( p1_u3203,n25858 );
   and U27305 ( n25860,n45625,n45626 );
   not U27306 ( p1_u3206,n25860 );
   and U27307 ( n25862,n45670,n45671 );
   not U27308 ( p1_u3197,n25862 );
   and U27309 ( n25864,n40955,n40956 );
   not U27310 ( p2_u2968,n25864 );
   and U27311 ( n25866,n40975,n40976 );
   not U27312 ( p2_u2964,n25866 );
   and U27313 ( n25868,n40945,n40946 );
   not U27314 ( p2_u2970,n25868 );
   and U27315 ( n25870,n36926,n36927 );
   not U27316 ( p2_u3218,n25870 );
   and U27317 ( n25872,n28904,n28905 );
   not U27318 ( p3_u3277,n25872 );
   and U27319 ( n25874,n45580,n45581 );
   not U27320 ( p1_u3215,n25874 );
   and U27321 ( n25876,n40970,n40971 );
   not U27322 ( p2_u2965,n25876 );
   and U27323 ( n25878,n40900,n40901 );
   not U27324 ( p2_u2979,n25878 );
   and U27325 ( n25880,n40980,n40981 );
   not U27326 ( p2_u2963,n25880 );
   and U27327 ( n25882,n40915,n40916 );
   not U27328 ( p2_u2976,n25882 );
   and U27329 ( n25884,n40965,n40966 );
   not U27330 ( p2_u2966,n25884 );
   and U27331 ( n25886,n40960,n40961 );
   not U27332 ( p2_u2967,n25886 );
   and U27333 ( n25888,n40905,n40906 );
   not U27334 ( p2_u2978,n25888 );
   and U27335 ( n25890,n40985,n40986 );
   not U27336 ( p2_u2962,n25890 );
   and U27337 ( n25892,n40940,n40941 );
   not U27338 ( p2_u2971,n25892 );
   and U27339 ( n25894,n40920,n40921 );
   not U27340 ( p2_u2975,n25894 );
   and U27341 ( n25896,n40930,n40931 );
   not U27342 ( p2_u2973,n25896 );
   and U27343 ( n25898,n40935,n40936 );
   not U27344 ( p2_u2972,n25898 );
   and U27345 ( n25900,n33184,n33185 );
   not U27346 ( p3_u2780,n25900 );
   and U27347 ( n25902,n33159,n33160 );
   not U27348 ( p3_u2785,n25902 );
   and U27349 ( n25904,n40925,n40926 );
   not U27350 ( p2_u2974,n25904 );
   and U27351 ( n25906,n40950,n40951 );
   not U27352 ( p2_u2969,n25906 );
   and U27353 ( n25908,n40895,n40896 );
   not U27354 ( p2_u2980,n25908 );
   and U27355 ( n25910,n40910,n40911 );
   not U27356 ( p2_u2977,n25910 );
   and U27357 ( n25912,n33174,n33175 );
   not U27358 ( p3_u2782,n25912 );
   and U27359 ( n25914,n33119,n33120 );
   not U27360 ( p3_u2793,n25914 );
   and U27361 ( n25916,n33164,n33165 );
   not U27362 ( p3_u2784,n25916 );
   and U27363 ( n25918,n33139,n33140 );
   not U27364 ( p3_u2789,n25918 );
   and U27365 ( n25920,n33189,n33190 );
   not U27366 ( p3_u2779,n25920 );
   and U27367 ( n25922,n33104,n33105 );
   not U27368 ( p3_u2796,n25922 );
   and U27369 ( n25924,n33149,n33150 );
   not U27370 ( p3_u2787,n25924 );
   and U27371 ( n25926,n33154,n33155 );
   not U27372 ( p3_u2786,n25926 );
   and U27373 ( n25928,n33109,n33110 );
   not U27374 ( p3_u2795,n25928 );
   and U27375 ( n25930,n33169,n33170 );
   not U27376 ( p3_u2783,n25930 );
   and U27377 ( n25932,n33194,n33195 );
   not U27378 ( p3_u2778,n25932 );
   and U27379 ( n25934,n33124,n33125 );
   not U27380 ( p3_u2792,n25934 );
   and U27381 ( n25936,n36796,n36797 );
   not U27382 ( p2_u3591,n25936 );
   and U27383 ( n25938,n33114,n33115 );
   not U27384 ( p3_u2794,n25938 );
   and U27385 ( n25940,n33129,n33130 );
   not U27386 ( p3_u2791,n25940 );
   and U27387 ( n25942,n33134,n33135 );
   not U27388 ( p3_u2790,n25942 );
   and U27389 ( n25944,n33144,n33145 );
   not U27390 ( p3_u2788,n25944 );
   and U27391 ( n25946,n33179,n33180 );
   not U27392 ( p3_u2781,n25946 );
   and U27393 ( n25948,n28613,n28614 );
   not U27394 ( u236,n25948 );
   and U27395 ( n25950,n28637,n28638 );
   not U27396 ( u232,n25950 );
   and U27397 ( n25952,n28661,n28662 );
   not U27398 ( u228,n25952 );
   and U27399 ( n25954,n28655,n28656 );
   not U27400 ( u229,n25954 );
   and U27401 ( n25956,n28583,n28584 );
   not U27402 ( u241,n25956 );
   and U27403 ( n25958,n28619,n28620 );
   not U27404 ( u235,n25958 );
   and U27405 ( n25960,n28571,n28572 );
   not U27406 ( u243,n25960 );
   and U27407 ( n25962,n28643,n28644 );
   not U27408 ( u231,n25962 );
   and U27409 ( n25964,n28631,n28632 );
   not U27410 ( u233,n25964 );
   and U27411 ( n25966,n28559,n28560 );
   not U27412 ( u245,n25966 );
   and U27413 ( n25968,n28732,n28733 );
   not U27414 ( u216,n25968 );
   and U27415 ( n25970,n28607,n28608 );
   not U27416 ( u237,n25970 );
   and U27417 ( n25972,n28625,n28626 );
   not U27418 ( u234,n25972 );
   and U27419 ( n25974,n28667,n28668 );
   not U27420 ( u227,n25974 );
   and U27421 ( n25976,n28601,n28602 );
   not U27422 ( u238,n25976 );
   and U27423 ( n25978,n28649,n28650 );
   not U27424 ( u230,n25978 );
   and U27425 ( n25980,n28595,n28596 );
   not U27426 ( u239,n25980 );
   and U27427 ( n25982,n28577,n28578 );
   not U27428 ( u242,n25982 );
   and U27429 ( n25984,n41322,n41323 );
   not U27430 ( p2_u2905,n25984 );
   and U27431 ( n25986,n41300,n41301 );
   not U27432 ( p2_u2910,n25986 );
   and U27433 ( n25988,n41293,n41294 );
   not U27434 ( p2_u2911,n25988 );
   and U27435 ( n25990,n41327,n41328 );
   not U27436 ( p2_u2904,n25990 );
   and U27437 ( n25992,n41312,n41313 );
   not U27438 ( p2_u2907,n25992 );
   and U27439 ( n25994,n28589,n28590 );
   not U27440 ( u240,n25994 );
   and U27441 ( n25996,n41788,n41789 );
   not U27442 ( p2_u2882,n25996 );
   and U27443 ( n25998,n29103,n29104 );
   not U27444 ( p3_u3029,n25998 );
   and U27445 ( n26000,n45712,n45713 );
   not U27446 ( p1_u3194,n26000 );
   and U27447 ( n26002,n41304,n41305 );
   not U27448 ( p2_u2909,n26002 );
   and U27449 ( n26004,n41308,n41309 );
   not U27450 ( p2_u2908,n26004 );
   and U27451 ( n26006,n41317,n41318 );
   not U27452 ( p2_u2906,n26006 );
   and U27453 ( n26008,n36252,n36253 );
   not U27454 ( p3_u2638,n26008 );
   and U27455 ( n26010,n52695,n52696 );
   not U27456 ( p1_u2807,n26010 );
   and U27457 ( n26012,n44673,n44674 );
   not U27458 ( p2_u2819,n26012 );
   and U27459 ( n26014,n34967,n34968 );
   not U27460 ( p3_u2676,n26014 );
   and U27461 ( n26016,n34945,n34946 );
   not U27462 ( p3_u2678,n26016 );
   and U27463 ( n26018,n28772,n28773 );
   not U27464 ( p3_u3298,n26018 );
   and U27465 ( n26020,n49759,n49760 );
   not U27466 ( p1_u2852,n26020 );
   and U27467 ( n26022,n49797,n49798 );
   not U27468 ( p1_u2845,n26022 );
   and U27469 ( n26024,n49781,n49782 );
   not U27470 ( p1_u2848,n26024 );
   and U27471 ( n26026,n49748,n49749 );
   not U27472 ( p1_u2854,n26026 );
   and U27473 ( n26028,n49764,n49765 );
   not U27474 ( p1_u2851,n26028 );
   and U27475 ( n26030,n49678,n49679 );
   not U27476 ( p1_u2869,n26030 );
   and U27477 ( n26032,n49668,n49669 );
   not U27478 ( p1_u2871,n26032 );
   and U27479 ( n26034,n49792,n49793 );
   not U27480 ( p1_u2846,n26034 );
   and U27481 ( n26036,n49753,n49754 );
   not U27482 ( p1_u2853,n26036 );
   and U27483 ( n26038,n49786,n49787 );
   not U27484 ( p1_u2847,n26038 );
   and U27485 ( n26040,n49808,n49809 );
   not U27486 ( p1_u2843,n26040 );
   and U27487 ( n26042,n49803,n49804 );
   not U27488 ( p1_u2844,n26042 );
   and U27489 ( n26044,n45320,n45321 );
   not U27490 ( p1_u3487,n26044 );
   and U27491 ( n26046,n36656,n36657 );
   not U27492 ( p2_u3609,n26046 );
   and U27493 ( n26048,n49661,n49662 );
   not U27494 ( p1_u2872,n26048 );
   and U27495 ( n26050,n49775,n49776 );
   not U27496 ( p1_u2849,n26050 );
   and U27497 ( n26052,n49770,n49771 );
   not U27498 ( p1_u2850,n26052 );
   and U27499 ( n26054,n49814,n49815 );
   not U27500 ( p1_u2842,n26054 );
   and U27501 ( n26056,n49406,n49407 );
   not U27502 ( p1_u2892,n26056 );
   and U27503 ( n26058,n49364,n49365 );
   not U27504 ( p1_u2899,n26058 );
   and U27505 ( n26060,n49346,n49347 );
   not U27506 ( p1_u2902,n26060 );
   and U27507 ( n26062,n49412,n49413 );
   not U27508 ( p1_u2891,n26062 );
   and U27509 ( n26064,n45374,n45375 );
   not U27510 ( p1_u3481,n26064 );
   and U27511 ( n26066,n28824,n28825 );
   not U27512 ( p3_u3292,n26066 );
   and U27513 ( n26068,n28766,n28767 );
   not U27514 ( p3_u3299,n26068 );
   and U27515 ( n26070,n44640,n44632 );
   not U27516 ( p2_u2820,n26070 );
   and U27517 ( n26072,n36247,n36248 );
   not U27518 ( p3_u2639,n26072 );
   and U27519 ( n26074,n52690,n52691 );
   not U27520 ( p1_u2808,n26074 );
   and U27521 ( n26076,n49382,n49383 );
   not U27522 ( p1_u2896,n26076 );
   and U27523 ( n26078,n49341,n49342 );
   not U27524 ( p1_u2903,n26078 );
   and U27525 ( n26080,n30089,n30090 );
   not U27526 ( p3_u2928,n26080 );
   and U27527 ( n26082,n30060,n30061 );
   not U27528 ( p3_u2931,n26082 );
   and U27529 ( n26084,n30105,n30106 );
   not U27530 ( p3_u2926,n26084 );
   and U27531 ( n26086,n30931,n30932 );
   not U27532 ( p3_u2857,n26086 );
   and U27533 ( n26088,n30878,n30879 );
   not U27534 ( p3_u2859,n26088 );
   and U27535 ( n26090,n30954,n30955 );
   not U27536 ( p3_u2856,n26090 );
   and U27537 ( n26092,n29851,n29852 );
   not U27538 ( p3_u2953,n26092 );
   and U27539 ( n26094,n30097,n30098 );
   not U27540 ( p3_u2927,n26094 );
   and U27541 ( n26096,n30113,n30114 );
   not U27542 ( p3_u2925,n26096 );
   and U27543 ( n26098,n30073,n30074 );
   not U27544 ( p3_u2930,n26098 );
   and U27545 ( n26100,n30121,n30122 );
   not U27546 ( p3_u2924,n26100 );
   and U27547 ( n26102,n30081,n30082 );
   not U27548 ( p3_u2929,n26102 );
   and U27549 ( n26104,n30160,n30161 );
   not U27550 ( p3_u2921,n26104 );
   and U27551 ( n26106,n29920,n29921 );
   not U27552 ( p3_u2946,n26106 );
   and U27553 ( n26108,n29801,n29802 );
   not U27554 ( p3_u2957,n26108 );
   and U27555 ( n26110,n29867,n29868 );
   not U27556 ( p3_u2951,n26110 );
   and U27557 ( n26112,n29830,n29831 );
   not U27558 ( p3_u2955,n26112 );
   and U27559 ( n26114,n29785,n29786 );
   not U27560 ( p3_u2959,n26114 );
   and U27561 ( n26116,n29883,n29884 );
   not U27562 ( p3_u2949,n26116 );
   and U27563 ( n26118,n29928,n29929 );
   not U27564 ( p3_u2945,n26118 );
   and U27565 ( n26120,n30152,n30153 );
   not U27566 ( p3_u2922,n26120 );
   and U27567 ( n26122,n29642,n29643 );
   not U27568 ( p3_u2972,n26122 );
   and U27569 ( n26124,n30192,n30193 );
   not U27570 ( p3_u2917,n26124 );
   and U27571 ( n26126,n29715,n29716 );
   not U27572 ( p3_u2965,n26126 );
   and U27573 ( n26128,n29907,n29908 );
   not U27574 ( p3_u2947,n26128 );
   and U27575 ( n26130,n29602,n29603 );
   not U27576 ( p3_u2977,n26130 );
   and U27577 ( n26132,n29960,n29961 );
   not U27578 ( p3_u2941,n26132 );
   and U27579 ( n26134,n30168,n30169 );
   not U27580 ( p3_u2920,n26134 );
   and U27581 ( n26136,n30184,n30185 );
   not U27582 ( p3_u2918,n26136 );
   and U27583 ( n26138,n29527,n29528 );
   not U27584 ( p3_u2984,n26138 );
   and U27585 ( n26140,n29519,n29520 );
   not U27586 ( p3_u2985,n26140 );
   and U27587 ( n26142,n30200,n30201 );
   not U27588 ( p3_u2916,n26142 );
   and U27589 ( n26144,n29543,n29544 );
   not U27590 ( p3_u2982,n26144 );
   and U27591 ( n26146,n29748,n29749 );
   not U27592 ( p3_u2963,n26146 );
   and U27593 ( n26148,n29944,n29945 );
   not U27594 ( p3_u2943,n26148 );
   and U27595 ( n26150,n30139,n30140 );
   not U27596 ( p3_u2923,n26150 );
   and U27597 ( n26152,n29691,n29692 );
   not U27598 ( p3_u2968,n26152 );
   and U27599 ( n26154,n29952,n29953 );
   not U27600 ( p3_u2942,n26154 );
   and U27601 ( n26156,n29675,n29676 );
   not U27602 ( p3_u2970,n26156 );
   and U27603 ( n26158,n29891,n29892 );
   not U27604 ( p3_u2948,n26158 );
   and U27605 ( n26160,n29769,n29770 );
   not U27606 ( p3_u2961,n26160 );
   and U27607 ( n26162,n29723,n29724 );
   not U27608 ( p3_u2964,n26162 );
   and U27609 ( n26164,n29581,n29582 );
   not U27610 ( p3_u2979,n26164 );
   and U27611 ( n26166,n29683,n29684 );
   not U27612 ( p3_u2969,n26166 );
   and U27613 ( n26168,n29777,n29778 );
   not U27614 ( p3_u2960,n26168 );
   and U27615 ( n26170,n29498,n29499 );
   not U27616 ( p3_u2987,n26170 );
   and U27617 ( n26172,n29511,n29512 );
   not U27618 ( p3_u2986,n26172 );
   and U27619 ( n26174,n29843,n29844 );
   not U27620 ( p3_u2954,n26174 );
   and U27621 ( n26176,n29626,n29627 );
   not U27622 ( p3_u2974,n26176 );
   and U27623 ( n26178,n29551,n29552 );
   not U27624 ( p3_u2981,n26178 );
   and U27625 ( n26180,n29859,n29860 );
   not U27626 ( p3_u2952,n26180 );
   and U27627 ( n26182,n29618,n29619 );
   not U27628 ( p3_u2975,n26182 );
   and U27629 ( n26184,n29634,n29635 );
   not U27630 ( p3_u2973,n26184 );
   and U27631 ( n26186,n29707,n29708 );
   not U27632 ( p3_u2966,n26186 );
   and U27633 ( n26188,n30176,n30177 );
   not U27634 ( p3_u2919,n26188 );
   and U27635 ( n26190,n29662,n29663 );
   not U27636 ( p3_u2971,n26190 );
   and U27637 ( n26192,n29809,n29810 );
   not U27638 ( p3_u2956,n26192 );
   and U27639 ( n26194,n29968,n29969 );
   not U27640 ( p3_u2940,n26194 );
   and U27641 ( n26196,n29936,n29937 );
   not U27642 ( p3_u2944,n26196 );
   and U27643 ( n26198,n29793,n29794 );
   not U27644 ( p3_u2958,n26198 );
   and U27645 ( n26200,n29761,n29762 );
   not U27646 ( p3_u2962,n26200 );
   and U27647 ( n26202,n29699,n29700 );
   not U27648 ( p3_u2967,n26202 );
   and U27649 ( n26204,n29559,n29560 );
   not U27650 ( p3_u2980,n26204 );
   and U27651 ( n26206,n29875,n29876 );
   not U27652 ( p3_u2950,n26206 );
   and U27653 ( n26208,n29594,n29595 );
   not U27654 ( p3_u2978,n26208 );
   and U27655 ( n26210,n29610,n29611 );
   not U27656 ( p3_u2976,n26210 );
   and U27657 ( n26212,n28715,n28716 );
   not U27658 ( u219,n26212 );
   and U27659 ( n26214,n28727,n28728 );
   not U27660 ( u217,n26214 );
   and U27661 ( n26216,n28565,n28566 );
   not U27662 ( u244,n26216 );
   and U27663 ( n26218,n28709,n28710 );
   not U27664 ( u220,n26218 );
   and U27665 ( n26220,n30790,n30791 );
   not U27666 ( p3_u2863,n26220 );
   and U27667 ( n26222,n29535,n29536 );
   not U27668 ( p3_u2983,n26222 );
   and U27669 ( n26224,n28545,n28546 );
   not U27670 ( u247,n26224 );
   and U27671 ( n26226,n28697,n28698 );
   not U27672 ( u222,n26226 );
   and U27673 ( n26228,n28691,n28692 );
   not U27674 ( u223,n26228 );
   and U27675 ( n26230,n28673,n28674 );
   not U27676 ( u226,n26230 );
   and U27677 ( n26232,n28703,n28704 );
   not U27678 ( u221,n26232 );
   and U27679 ( n26234,n28721,n28722 );
   not U27680 ( u218,n26234 );
   and U27681 ( n26236,n31657,n31658 );
   not U27682 ( p3_u2833,n26236 );
   and U27683 ( n26238,n31545,n31546 );
   not U27684 ( p3_u2836,n26238 );
   and U27685 ( n26240,n31522,n31523 );
   not U27686 ( p3_u2837,n26240 );
   and U27687 ( n26242,n28553,n28554 );
   not U27688 ( u246,n26242 );
   and U27689 ( n26244,n28685,n28686 );
   not U27690 ( u224,n26244 );
   and U27691 ( n26246,n28679,n28680 );
   not U27692 ( u225,n26246 );
   and U27693 ( n26248,n44636,n44637 );
   not U27694 ( p2_u2821,n26248 );
   and U27695 ( n26250,n45368,n45369 );
   not U27696 ( p1_u3482,n26250 );
   and U27697 ( n26252,n28818,n28819 );
   not U27698 ( p3_u3293,n26252 );
   and U27699 ( n26254,n31143,n31144 );
   not U27700 ( p3_u2849,n26254 );
   and U27701 ( n26256,n31114,n31115 );
   not U27702 ( p3_u2850,n26256 );
   and U27703 ( n26258,n31260,n31261 );
   not U27704 ( p3_u2845,n26258 );
   and U27705 ( n26260,n30663,n30664 );
   not U27706 ( p3_u2873,n26260 );
   and U27707 ( n26262,n30706,n30707 );
   not U27708 ( p3_u2869,n26262 );
   and U27709 ( n26264,n30806,n30807 );
   not U27710 ( p3_u2862,n26264 );
   and U27711 ( n26266,n30695,n30696 );
   not U27712 ( p3_u2870,n26266 );
   and U27713 ( n26268,n44622,n44623 );
   not U27714 ( p2_u2823,n26268 );
   and U27715 ( n26270,n44628,n44629 );
   not U27716 ( p2_u2822,n26270 );
   and U27717 ( n26272,n41243,n41244 );
   not U27718 ( p2_u2916,n26272 );
   and U27719 ( n26274,n41222,n41223 );
   not U27720 ( p2_u2918,n26274 );
   and U27721 ( n26276,n30652,n30653 );
   not U27722 ( p3_u2874,n26276 );
   and U27723 ( n26278,n30634,n30635 );
   not U27724 ( p3_u2875,n26278 );
   and U27725 ( n26280,n30684,n30685 );
   not U27726 ( p3_u2871,n26280 );
   and U27727 ( n26282,n30674,n30675 );
   not U27728 ( p3_u2872,n26282 );
   and U27729 ( n26284,n39216,n39217 );
   not U27730 ( p2_u3025,n26284 );
   and U27731 ( n26286,n39189,n39190 );
   not U27732 ( p2_u3026,n26286 );
   and U27733 ( n26288,n39265,n39266 );
   not U27734 ( p2_u3023,n26288 );
   and U27735 ( n26290,n39026,n39027 );
   not U27736 ( p2_u3033,n26290 );
   and U27737 ( n26292,n41252,n41253 );
   not U27738 ( p2_u2915,n26292 );
   and U27739 ( n26294,n41233,n41234 );
   not U27740 ( p2_u2917,n26294 );
   and U27741 ( n26296,n33229,n33230 );
   not U27742 ( p3_u2770,n26296 );
   and U27743 ( n26298,n39284,n39285 );
   not U27744 ( p2_u3022,n26298 );
   and U27745 ( n26300,n39361,n39362 );
   not U27746 ( p2_u3019,n26300 );
   and U27747 ( n26302,n39399,n39400 );
   not U27748 ( p2_u3017,n26302 );
   and U27749 ( n26304,n39045,n39046 );
   not U27750 ( p2_u3032,n26304 );
   and U27751 ( n26306,n39332,n39333 );
   not U27752 ( p2_u3020,n26306 );
   and U27753 ( n26308,n40890,n40891 );
   not U27754 ( p2_u2981,n26308 );
   and U27755 ( n26310,n41012,n41013 );
   not U27756 ( p2_u2956,n26310 );
   and U27757 ( n26312,n33209,n33210 );
   not U27758 ( p3_u2775,n26312 );
   and U27759 ( n26314,n41004,n41005 );
   not U27760 ( p2_u2958,n26314 );
   and U27761 ( n26316,n40990,n40991 );
   not U27762 ( p2_u2961,n26316 );
   and U27763 ( n26318,n33099,n33100 );
   not U27764 ( p3_u2797,n26318 );
   and U27765 ( n26320,n33217,n33218 );
   not U27766 ( p3_u2773,n26320 );
   and U27767 ( n26322,n40995,n40996 );
   not U27768 ( p2_u2960,n26322 );
   and U27769 ( n26324,n33221,n33222 );
   not U27770 ( p3_u2772,n26324 );
   and U27771 ( n26326,n33204,n33205 );
   not U27772 ( p3_u2776,n26326 );
   and U27773 ( n26328,n33225,n33226 );
   not U27774 ( p3_u2771,n26328 );
   and U27775 ( n26330,n41024,n41025 );
   not U27776 ( p2_u2953,n26330 );
   and U27777 ( n26332,n41028,n41029 );
   not U27778 ( p2_u2952,n26332 );
   and U27779 ( n26334,n33213,n33214 );
   not U27780 ( p3_u2774,n26334 );
   and U27781 ( n26336,n40882,n40883 );
   not U27782 ( p2_u2982,n26336 );
   and U27783 ( n26338,n41000,n41001 );
   not U27784 ( p2_u2959,n26338 );
   and U27785 ( n26340,n41008,n41009 );
   not U27786 ( p2_u2957,n26340 );
   and U27787 ( n26342,n33237,n33238 );
   not U27788 ( p3_u2768,n26342 );
   and U27789 ( n26344,n31320,n31321 );
   not U27790 ( p3_u2843,n26344 );
   and U27791 ( n26346,n41020,n41021 );
   not U27792 ( p2_u2954,n26346 );
   and U27793 ( n26348,n33091,n33092 );
   not U27794 ( p3_u2798,n26348 );
   and U27795 ( n26350,n33233,n33234 );
   not U27796 ( p3_u2769,n26350 );
   and U27797 ( n26352,n33199,n33200 );
   not U27798 ( p3_u2777,n26352 );
   and U27799 ( n26354,n41016,n41017 );
   not U27800 ( p2_u2955,n26354 );
   and U27801 ( n26356,n39380,n39381 );
   not U27802 ( p2_u3018,n26356 );
   and U27803 ( n26358,n41263,n41264 );
   not U27804 ( p2_u2914,n26358 );
   and U27805 ( n26360,n38997,n38998 );
   not U27806 ( p2_u3034,n26360 );
   and U27807 ( n26362,n38852,n38853 );
   not U27808 ( p2_u3040,n26362 );
   and U27809 ( n26364,n38833,n38834 );
   not U27810 ( p2_u3041,n26364 );
   and U27811 ( n26366,n45489,n45490 );
   not U27812 ( p1_u3468,n26366 );
   and U27813 ( n26368,n41207,n41208 );
   not U27814 ( p2_u2919,n26368 );
   and U27815 ( n26370,n39313,n39314 );
   not U27816 ( p2_u3021,n26370 );
   and U27817 ( n26372,n39235,n39236 );
   not U27818 ( p2_u3024,n26372 );
   and U27819 ( n26374,n38806,n38807 );
   not U27820 ( p2_u3042,n26374 );
   and U27821 ( n26376,n39074,n39075 );
   not U27822 ( p2_u3031,n26376 );
   and U27823 ( n26378,n38881,n38882 );
   not U27824 ( p2_u3039,n26378 );
   and U27825 ( n26380,n35985,n35986 );
   not U27826 ( p3_u2646,n26380 );
   and U27827 ( n26382,n35893,n35894 );
   not U27828 ( p3_u2650,n26382 );
   and U27829 ( n26384,n29066,n29067 );
   not U27830 ( p3_u3031,n26384 );
   and U27831 ( n26386,n36773,n36774 );
   not U27832 ( p2_u3595,n26386 );
   and U27833 ( n26388,n41274,n41275 );
   not U27834 ( p2_u2913,n26388 );
   and U27835 ( n26390,n38738,n38739 );
   not U27836 ( p2_u3045,n26390 );
   and U27837 ( n26392,n45676,n45677 );
   not U27838 ( p1_u3196,n26392 );
   and U27839 ( n26394,n36124,n36125 );
   not U27840 ( p3_u2640,n26394 );
   and U27841 ( n26396,n35939,n35940 );
   not U27842 ( p3_u2648,n26396 );
   and U27843 ( n26398,n28875,n28876 );
   not U27844 ( p3_u3284,n26398 );
   and U27845 ( n26400,n36103,n36104 );
   not U27846 ( p3_u2641,n26400 );
   and U27847 ( n26402,n36032,n36033 );
   not U27848 ( p3_u2644,n26402 );
   and U27849 ( n26404,n29431,n29432 );
   not U27850 ( p3_u2991,n26404 );
   and U27851 ( n26406,n29378,n29379 );
   not U27852 ( p3_u2995,n26406 );
   and U27853 ( n26408,n29455,n29456 );
   not U27854 ( p3_u2989,n26408 );
   and U27855 ( n26410,n29419,n29420 );
   not U27856 ( p3_u2992,n26410 );
   and U27857 ( n26412,n29467,n29468 );
   not U27858 ( p3_u2988,n26412 );
   and U27859 ( n26414,n36963,n36964 );
   not U27860 ( p2_u3211,n26414 );
   and U27861 ( n26416,n47987,n47988 );
   not U27862 ( p1_u3008,n26416 );
   and U27863 ( n26418,n47868,n47869 );
   not U27864 ( p1_u3013,n26418 );
   and U27865 ( n26420,n31056,n31057 );
   not U27866 ( p3_u2852,n26420 );
   and U27867 ( n26422,n29407,n29408 );
   not U27868 ( p3_u2993,n26422 );
   and U27869 ( n26424,n29443,n29444 );
   not U27870 ( p3_u2990,n26424 );
   and U27871 ( n26426,n29395,n29396 );
   not U27872 ( p3_u2994,n26426 );
   and U27873 ( n26428,n47522,n47523 );
   not U27874 ( p1_u3028,n26428 );
   and U27875 ( n26430,n47587,n47588 );
   not U27876 ( p1_u3025,n26430 );
   and U27877 ( n26432,n47615,n47616 );
   not U27878 ( p1_u3024,n26432 );
   and U27879 ( n26434,n49606,n49607 );
   not U27880 ( p1_u2873,n26434 );
   and U27881 ( n26436,n48082,n48083 );
   not U27882 ( p1_u3004,n26436 );
   and U27883 ( n26438,n49830,n49831 );
   not U27884 ( p1_u2840,n26438 );
   and U27885 ( n26440,n37558,n37559 );
   not U27886 ( p2_u3147,n26440 );
   and U27887 ( n26442,n37542,n37543 );
   not U27888 ( p2_u3149,n26442 );
   and U27889 ( n26444,n37550,n37551 );
   not U27890 ( p2_u3148,n26444 );
   and U27891 ( n26446,n48125,n48126 );
   not U27892 ( p1_u3002,n26446 );
   and U27893 ( n26448,n47849,n47850 );
   not U27894 ( p1_u3014,n26448 );
   and U27895 ( n26450,n47774,n47775 );
   not U27896 ( p1_u3017,n26450 );
   and U27897 ( n26452,n32768,n32769 );
   not U27898 ( p3_u2803,n26452 );
   and U27899 ( n26454,n37534,n37535 );
   not U27900 ( p2_u3150,n26454 );
   and U27901 ( n26456,n37521,n37522 );
   not U27902 ( p2_u3151,n26456 );
   and U27903 ( n26458,n37582,n37583 );
   not U27904 ( p2_u3144,n26458 );
   and U27905 ( n26460,n37574,n37575 );
   not U27906 ( p2_u3145,n26460 );
   and U27907 ( n26462,n37566,n37567 );
   not U27908 ( p2_u3146,n26462 );
   and U27909 ( n26464,n37220,n37221 );
   not U27910 ( p2_u3175,n26464 );
   and U27911 ( n26466,n37237,n37238 );
   not U27912 ( p2_u3174,n26466 );
   and U27913 ( n26468,n37261,n37262 );
   not U27914 ( p2_u3172,n26468 );
   and U27915 ( n26470,n37273,n37274 );
   not U27916 ( p2_u3171,n26470 );
   and U27917 ( n26472,n37297,n37298 );
   not U27918 ( p2_u3169,n26472 );
   and U27919 ( n26474,n37309,n37310 );
   not U27920 ( p2_u3168,n26474 );
   and U27921 ( n26476,n39439,n39440 );
   not U27922 ( p2_u3015,n26476 );
   and U27923 ( n26478,n48527,n48528 );
   not U27924 ( p1_u2984,n26478 );
   and U27925 ( n26480,n48552,n48553 );
   not U27926 ( p1_u2983,n26480 );
   and U27927 ( n26482,n39642,n39643 );
   not U27928 ( p2_u3011,n26482 );
   and U27929 ( n26484,n37285,n37286 );
   not U27930 ( p2_u3170,n26484 );
   and U27931 ( n26486,n37249,n37250 );
   not U27932 ( p2_u3173,n26486 );
   and U27933 ( n26488,n38788,n38789 );
   not U27934 ( p2_u3043,n26488 );
   and U27935 ( n26490,n38929,n38930 );
   not U27936 ( p2_u3037,n26490 );
   and U27937 ( n26492,n48676,n48677 );
   not U27938 ( p1_u2976,n26492 );
   and U27939 ( n26494,n38978,n38979 );
   not U27940 ( p2_u3035,n26494 );
   and U27941 ( n26496,n48318,n48319 );
   not U27942 ( p1_u2997,n26496 );
   and U27943 ( n26498,n48588,n48589 );
   not U27944 ( p1_u2981,n26498 );
   and U27945 ( n26500,n30452,n30453 );
   not U27946 ( p3_u2892,n26500 );
   and U27947 ( n26502,n30537,n30538 );
   not U27948 ( p3_u2884,n26502 );
   and U27949 ( n26504,n30616,n30617 );
   not U27950 ( p3_u2876,n26504 );
   and U27951 ( n26506,n48412,n48413 );
   not U27952 ( p1_u2991,n26506 );
   and U27953 ( n26508,n38949,n38950 );
   not U27954 ( p2_u3036,n26508 );
   and U27955 ( n26510,n48512,n48513 );
   not U27956 ( p1_u2985,n26510 );
   and U27957 ( n26512,n30352,n30353 );
   not U27958 ( p3_u2902,n26512 );
   and U27959 ( n26514,n30529,n30530 );
   not U27960 ( p3_u2885,n26514 );
   and U27961 ( n26516,n30584,n30585 );
   not U27962 ( p3_u2880,n26516 );
   and U27963 ( n26518,n30436,n30437 );
   not U27964 ( p3_u2894,n26518 );
   and U27965 ( n26520,n30718,n30719 );
   not U27966 ( p3_u2868,n26520 );
   and U27967 ( n26522,n30372,n30373 );
   not U27968 ( p3_u2900,n26522 );
   and U27969 ( n26524,n30444,n30445 );
   not U27970 ( p3_u2893,n26524 );
   and U27971 ( n26526,n30362,n30363 );
   not U27972 ( p3_u2901,n26526 );
   and U27973 ( n26528,n30404,n30405 );
   not U27974 ( p3_u2898,n26528 );
   and U27975 ( n26530,n30568,n30569 );
   not U27976 ( p3_u2882,n26530 );
   and U27977 ( n26532,n30342,n30343 );
   not U27978 ( p3_u2903,n26532 );
   and U27979 ( n26534,n30592,n30593 );
   not U27980 ( p3_u2879,n26534 );
   and U27981 ( n26536,n30412,n30413 );
   not U27982 ( p3_u2897,n26536 );
   and U27983 ( n26538,n30600,n30601 );
   not U27984 ( p3_u2878,n26538 );
   and U27985 ( n26540,n30322,n30323 );
   not U27986 ( p3_u2905,n26540 );
   and U27987 ( n26542,n30420,n30421 );
   not U27988 ( p3_u2896,n26542 );
   and U27989 ( n26544,n30332,n30333 );
   not U27990 ( p3_u2904,n26544 );
   and U27991 ( n26546,n30312,n30313 );
   not U27992 ( p3_u2906,n26546 );
   and U27993 ( n26548,n30505,n30506 );
   not U27994 ( p3_u2888,n26548 );
   and U27995 ( n26550,n30489,n30490 );
   not U27996 ( p3_u2890,n26550 );
   and U27997 ( n26552,n30513,n30514 );
   not U27998 ( p3_u2887,n26552 );
   and U27999 ( n26554,n30497,n30498 );
   not U28000 ( p3_u2889,n26554 );
   and U28001 ( n26556,n30521,n30522 );
   not U28002 ( p3_u2886,n26556 );
   and U28003 ( n26558,n30576,n30577 );
   not U28004 ( p3_u2881,n26558 );
   and U28005 ( n26560,n30476,n30477 );
   not U28006 ( p3_u2891,n26560 );
   and U28007 ( n26562,n30391,n30392 );
   not U28008 ( p3_u2899,n26562 );
   and U28009 ( n26564,n30297,n30298 );
   not U28010 ( p3_u2907,n26564 );
   and U28011 ( n26566,n30555,n30556 );
   not U28012 ( p3_u2883,n26566 );
   and U28013 ( n26568,n30608,n30609 );
   not U28014 ( p3_u2877,n26568 );
   and U28015 ( n26570,n30428,n30429 );
   not U28016 ( p3_u2895,n26570 );
   and U28017 ( n26572,n48656,n48657 );
   not U28018 ( p1_u2977,n26572 );
   and U28019 ( n26574,n48482,n48483 );
   not U28020 ( p1_u2987,n26574 );
   and U28021 ( n26576,n48350,n48351 );
   not U28022 ( p1_u2995,n26576 );
   and U28023 ( n26578,n48728,n48729 );
   not U28024 ( p1_u2973,n26578 );
   and U28025 ( n26580,n48788,n48789 );
   not U28026 ( p1_u2970,n26580 );
   and U28027 ( n26582,n48803,n48804 );
   not U28028 ( p1_u2969,n26582 );
   and U28029 ( n26584,n47476,n47477 );
   not U28030 ( p1_u3030,n26584 );
   and U28031 ( n26586,n47493,n47494 );
   not U28032 ( p1_u3029,n26586 );
   and U28033 ( n26588,n32452,n32453 );
   not U28034 ( p3_u2812,n26588 );
   and U28035 ( n26590,n50469,n50470 );
   not U28036 ( p1_u2814,n26590 );
   and U28037 ( n26592,n32865,n32866 );
   not U28038 ( p3_u2800,n26592 );
   and U28039 ( n26594,n48606,n48607 );
   not U28040 ( p1_u2980,n26594 );
   and U28041 ( n26596,n48378,n48379 );
   not U28042 ( p1_u2993,n26596 );
   and U28043 ( n26598,n32513,n32514 );
   not U28044 ( p3_u2810,n26598 );
   and U28045 ( n26600,n48621,n48622 );
   not U28046 ( p1_u2979,n26600 );
   and U28047 ( n26602,n48695,n48696 );
   not U28048 ( p1_u2975,n26602 );
   and U28049 ( n26604,n32662,n32663 );
   not U28050 ( p3_u2806,n26604 );
   and U28051 ( n26606,n32381,n32382 );
   not U28052 ( p3_u2814,n26606 );
   and U28053 ( n26608,n35962,n35963 );
   not U28054 ( p3_u2647,n26608 );
   and U28055 ( n26610,n35847,n35848 );
   not U28056 ( p3_u2652,n26610 );
   and U28057 ( n26612,n48765,n48766 );
   not U28058 ( p1_u2971,n26612 );
   and U28059 ( n26614,n32590,n32591 );
   not U28060 ( p3_u2808,n26614 );
   and U28061 ( n26616,n32322,n32323 );
   not U28062 ( p3_u2816,n26616 );
   and U28063 ( n26618,n48446,n48447 );
   not U28064 ( p1_u2989,n26618 );
   and U28065 ( n26620,n35916,n35917 );
   not U28066 ( p3_u2649,n26620 );
   and U28067 ( n26622,n35742,n35743 );
   not U28068 ( p3_u2656,n26622 );
   and U28069 ( n26624,n36079,n36080 );
   not U28070 ( p3_u2642,n26624 );
   and U28071 ( n26626,n35540,n35541 );
   not U28072 ( p3_u2664,n26626 );
   and U28073 ( n26628,n36055,n36056 );
   not U28074 ( p3_u2643,n26628 );
   and U28075 ( n26630,n35871,n35872 );
   not U28076 ( p3_u2651,n26630 );
   and U28077 ( n26632,n39623,n39624 );
   not U28078 ( p2_u3012,n26632 );
   and U28079 ( n26634,n40185,n40186 );
   not U28080 ( p2_u2984,n26634 );
   and U28081 ( n26636,n50575,n50576 );
   not U28082 ( p1_u2809,n26636 );
   and U28083 ( n26638,n36008,n36009 );
   not U28084 ( p3_u2645,n26638 );
   and U28085 ( n26640,n35489,n35490 );
   not U28086 ( p3_u2666,n26640 );
   and U28087 ( n26642,n35694,n35695 );
   not U28088 ( p3_u2658,n26642 );
   and U28089 ( n26644,n37743,n37744 );
   not U28090 ( p2_u3130,n26644 );
   and U28091 ( n26646,n39605,n39606 );
   not U28092 ( p2_u3013,n26646 );
   and U28093 ( n26648,n49857,n49858 );
   not U28094 ( p1_u2839,n26648 );
   and U28095 ( n26650,n30823,n30824 );
   not U28096 ( p3_u2861,n26650 );
   and U28097 ( n26652,n41285,n41286 );
   not U28098 ( p2_u2912,n26652 );
   and U28099 ( n26654,n32087,n32088 );
   not U28100 ( p3_u2824,n26654 );
   and U28101 ( n26656,n49526,n49527 );
   not U28102 ( p1_u2880,n26656 );
   and U28103 ( n26658,n49434,n49435 );
   not U28104 ( p1_u2888,n26658 );
   and U28105 ( n26660,n49548,n49549 );
   not U28106 ( p1_u2878,n26660 );
   and U28107 ( n26662,n37698,n37699 );
   not U28108 ( p2_u3135,n26662 );
   and U28109 ( n26664,n37751,n37752 );
   not U28110 ( p2_u3129,n26664 );
   and U28111 ( n26666,n49504,n49505 );
   not U28112 ( p1_u2882,n26666 );
   and U28113 ( n26668,n49537,n49538 );
   not U28114 ( p1_u2879,n26668 );
   and U28115 ( n26670,n31918,n31919 );
   not U28116 ( p3_u2830,n26670 );
   and U28117 ( n26672,n49570,n49571 );
   not U28118 ( p1_u2876,n26672 );
   and U28119 ( n26674,n49515,n49516 );
   not U28120 ( p1_u2881,n26674 );
   and U28121 ( n26676,n49559,n49560 );
   not U28122 ( p1_u2877,n26676 );
   and U28123 ( n26678,n37735,n37736 );
   not U28124 ( p2_u3131,n26678 );
   and U28125 ( n26680,n37727,n37728 );
   not U28126 ( p2_u3132,n26680 );
   and U28127 ( n26682,n49493,n49494 );
   not U28128 ( p1_u2883,n26682 );
   and U28129 ( n26684,n37719,n37720 );
   not U28130 ( p2_u3133,n26684 );
   and U28131 ( n26686,n37711,n37712 );
   not U28132 ( p2_u3134,n26686 );
   and U28133 ( n26688,n37759,n37760 );
   not U28134 ( p2_u3128,n26688 );
   and U28135 ( n26690,n49581,n49582 );
   not U28136 ( p1_u2875,n26690 );
   and U28137 ( n26692,n46487,n46488 );
   not U28138 ( p1_u3108,n26692 );
   and U28139 ( n26694,n46578,n46579 );
   not U28140 ( p1_u3099,n26694 );
   and U28141 ( n26696,n46533,n46534 );
   not U28142 ( p1_u3104,n26696 );
   and U28143 ( n26698,n32044,n32045 );
   not U28144 ( p3_u2825,n26698 );
   and U28145 ( n26700,n49482,n49483 );
   not U28146 ( p1_u2884,n26700 );
   and U28147 ( n26702,n32143,n32144 );
   not U28148 ( p3_u2822,n26702 );
   and U28149 ( n26704,n46495,n46496 );
   not U28150 ( p1_u3107,n26704 );
   and U28151 ( n26706,n46337,n46338 );
   not U28152 ( p1_u3121,n26706 );
   and U28153 ( n26708,n37671,n37672 );
   not U28154 ( p2_u3136,n26708 );
   and U28155 ( n26710,n46546,n46547 );
   not U28156 ( p1_u3103,n26710 );
   and U28157 ( n26712,n46570,n46571 );
   not U28158 ( p1_u3100,n26712 );
   and U28159 ( n26714,n46450,n46451 );
   not U28160 ( p1_u3112,n26714 );
   and U28161 ( n26716,n46329,n46330 );
   not U28162 ( p1_u3122,n26716 );
   and U28163 ( n26718,n37663,n37664 );
   not U28164 ( p2_u3137,n26718 );
   and U28165 ( n26720,n46393,n46394 );
   not U28166 ( p1_u3117,n26720 );
   and U28167 ( n26722,n46511,n46512 );
   not U28168 ( p1_u3105,n26722 );
   and U28169 ( n26724,n46594,n46595 );
   not U28170 ( p1_u3097,n26724 );
   and U28171 ( n26726,n37631,n37632 );
   not U28172 ( p2_u3141,n26726 );
   and U28173 ( n26728,n37655,n37656 );
   not U28174 ( p2_u3138,n26728 );
   and U28175 ( n26730,n46276,n46277 );
   not U28176 ( p1_u3128,n26730 );
   and U28177 ( n26732,n30021,n30022 );
   not U28178 ( p3_u2935,n26732 );
   and U28179 ( n26734,n37610,n37611 );
   not U28180 ( p2_u3143,n26734 );
   and U28181 ( n26736,n37647,n37648 );
   not U28182 ( p2_u3139,n26736 );
   and U28183 ( n26738,n46313,n46314 );
   not U28184 ( p1_u3124,n26738 );
   and U28185 ( n26740,n46425,n46426 );
   not U28186 ( p1_u3113,n26740 );
   and U28187 ( n26742,n37623,n37624 );
   not U28188 ( p2_u3142,n26742 );
   and U28189 ( n26744,n46289,n46290 );
   not U28190 ( p1_u3127,n26744 );
   and U28191 ( n26746,n46401,n46402 );
   not U28192 ( p1_u3116,n26746 );
   and U28193 ( n26748,n46364,n46365 );
   not U28194 ( p1_u3120,n26748 );
   and U28195 ( n26750,n37639,n37640 );
   not U28196 ( p2_u3140,n26750 );
   and U28197 ( n26752,n31036,n31037 );
   not U28198 ( p3_u2853,n26752 );
   and U28199 ( n26754,n46321,n46322 );
   not U28200 ( p1_u3123,n26754 );
   and U28201 ( n26756,n30005,n30006 );
   not U28202 ( p3_u2937,n26756 );
   and U28203 ( n26758,n29997,n29998 );
   not U28204 ( p3_u2938,n26758 );
   and U28205 ( n26760,n37781,n37782 );
   not U28206 ( p2_u3127,n26760 );
   and U28207 ( n26762,n46409,n46410 );
   not U28208 ( p1_u3115,n26762 );
   and U28209 ( n26764,n46463,n46464 );
   not U28210 ( p1_u3111,n26764 );
   and U28211 ( n26766,n30037,n30038 );
   not U28212 ( p3_u2933,n26766 );
   and U28213 ( n26768,n46385,n46386 );
   not U28214 ( p1_u3118,n26768 );
   and U28215 ( n26770,n46297,n46298 );
   not U28216 ( p1_u3126,n26770 );
   and U28217 ( n26772,n46586,n46587 );
   not U28218 ( p1_u3098,n26772 );
   and U28219 ( n26774,n30013,n30014 );
   not U28220 ( p3_u2936,n26774 );
   and U28221 ( n26776,n30029,n30030 );
   not U28222 ( p3_u2934,n26776 );
   and U28223 ( n26778,n46471,n46472 );
   not U28224 ( p1_u3110,n26778 );
   and U28225 ( n26780,n30045,n30046 );
   not U28226 ( p3_u2932,n26780 );
   and U28227 ( n26782,n37834,n37835 );
   not U28228 ( p2_u3121,n26782 );
   and U28229 ( n26784,n29984,n29985 );
   not U28230 ( p3_u2939,n26784 );
   and U28231 ( n26786,n46503,n46504 );
   not U28232 ( p1_u3106,n26786 );
   and U28233 ( n26788,n46417,n46418 );
   not U28234 ( p1_u3114,n26788 );
   and U28235 ( n26790,n37826,n37827 );
   not U28236 ( p2_u3122,n26790 );
   and U28237 ( n26792,n46305,n46306 );
   not U28238 ( p1_u3125,n26792 );
   and U28239 ( n26794,n46377,n46378 );
   not U28240 ( p1_u3119,n26794 );
   and U28241 ( n26796,n46479,n46480 );
   not U28242 ( p1_u3109,n26796 );
   and U28243 ( n26798,n37842,n37843 );
   not U28244 ( p2_u3120,n26798 );
   and U28245 ( n26800,n37794,n37795 );
   not U28246 ( p2_u3126,n26800 );
   and U28247 ( n26802,n46554,n46555 );
   not U28248 ( p1_u3102,n26802 );
   and U28249 ( n26804,n37802,n37803 );
   not U28250 ( p2_u3125,n26804 );
   and U28251 ( n26806,n37810,n37811 );
   not U28252 ( p2_u3124,n26806 );
   and U28253 ( n26808,n37818,n37819 );
   not U28254 ( p2_u3123,n26808 );
   and U28255 ( n26810,n46562,n46563 );
   not U28256 ( p1_u3101,n26810 );
   and U28257 ( n26812,n41544,n41545 );
   not U28258 ( p2_u2890,n26812 );
   and U28259 ( n26814,n39662,n39663 );
   not U28260 ( p2_u3010,n26814 );
   and U28261 ( n26816,n46070,n46071 );
   not U28262 ( p1_u3145,n26816 );
   and U28263 ( n26818,n41512,n41513 );
   not U28264 ( p2_u2892,n26818 );
   and U28265 ( n26820,n50355,n50356 );
   not U28266 ( p1_u2819,n26820 );
   and U28267 ( n26822,n48636,n48637 );
   not U28268 ( p1_u2978,n26822 );
   and U28269 ( n26824,n46734,n46735 );
   not U28270 ( p1_u3085,n26824 );
   and U28271 ( n26826,n46705,n46706 );
   not U28272 ( p1_u3088,n26826 );
   and U28273 ( n26828,n41496,n41497 );
   not U28274 ( p2_u2893,n26828 );
   and U28275 ( n26830,n41432,n41433 );
   not U28276 ( p2_u2897,n26830 );
   and U28277 ( n26832,n46758,n46759 );
   not U28278 ( p1_u3082,n26832 );
   and U28279 ( n26834,n39720,n39721 );
   not U28280 ( p2_u3007,n26834 );
   and U28281 ( n26836,n40146,n40147 );
   not U28282 ( p2_u2986,n26836 );
   and U28283 ( n26838,n41528,n41529 );
   not U28284 ( p2_u2891,n26838 );
   and U28285 ( n26840,n39777,n39778 );
   not U28286 ( p2_u3004,n26840 );
   and U28287 ( n26842,n46030,n46031 );
   not U28288 ( p1_u3150,n26842 );
   and U28289 ( n26844,n46718,n46719 );
   not U28290 ( p1_u3087,n26844 );
   and U28291 ( n26846,n41400,n41401 );
   not U28292 ( p2_u2899,n26846 );
   and U28293 ( n26848,n46062,n46063 );
   not U28294 ( p1_u3146,n26848 );
   and U28295 ( n26850,n46726,n46727 );
   not U28296 ( p1_u3086,n26850 );
   and U28297 ( n26852,n46022,n46023 );
   not U28298 ( p1_u3151,n26852 );
   and U28299 ( n26854,n41708,n41709 );
   not U28300 ( p2_u2888,n26854 );
   and U28301 ( n26856,n41480,n41481 );
   not U28302 ( p2_u2894,n26856 );
   and U28303 ( n26858,n46054,n46055 );
   not U28304 ( p1_u3147,n26858 );
   and U28305 ( n26860,n39838,n39839 );
   not U28306 ( p2_u3001,n26860 );
   and U28307 ( n26862,n46046,n46047 );
   not U28308 ( p1_u3148,n26862 );
   and U28309 ( n26864,n46009,n46010 );
   not U28310 ( p1_u3152,n26864 );
   and U28311 ( n26866,n46766,n46767 );
   not U28312 ( p1_u3081,n26866 );
   and U28313 ( n26868,n39901,n39902 );
   not U28314 ( p2_u2998,n26868 );
   and U28315 ( n26870,n41464,n41465 );
   not U28316 ( p2_u2895,n26870 );
   and U28317 ( n26872,n46038,n46039 );
   not U28318 ( p1_u3149,n26872 );
   and U28319 ( n26874,n46742,n46743 );
   not U28320 ( p1_u3084,n26874 );
   and U28321 ( n26876,n41416,n41417 );
   not U28322 ( p2_u2898,n26876 );
   and U28323 ( n26878,n48709,n48710 );
   not U28324 ( p1_u2974,n26878 );
   and U28325 ( n26880,n48573,n48574 );
   not U28326 ( p1_u2982,n26880 );
   and U28327 ( n26882,n40017,n40018 );
   not U28328 ( p2_u2992,n26882 );
   and U28329 ( n26884,n39961,n39962 );
   not U28330 ( p2_u2995,n26884 );
   and U28331 ( n26886,n40203,n40204 );
   not U28332 ( p2_u2983,n26886 );
   and U28333 ( n26888,n46750,n46751 );
   not U28334 ( p1_u3083,n26888 );
   and U28335 ( n26890,n50447,n50448 );
   not U28336 ( p1_u2815,n26890 );
   and U28337 ( n26892,n41335,n41336 );
   not U28338 ( p2_u2903,n26892 );
   and U28339 ( n26894,n41448,n41449 );
   not U28340 ( p2_u2896,n26894 );
   and U28341 ( n26896,n30281,n30282 );
   not U28342 ( p3_u2908,n26896 );
   and U28343 ( n26898,n30249,n30250 );
   not U28344 ( p3_u2912,n26898 );
   and U28345 ( n26900,n30265,n30266 );
   not U28346 ( p3_u2910,n26900 );
   and U28347 ( n26902,n30241,n30242 );
   not U28348 ( p3_u2913,n26902 );
   and U28349 ( n26904,n30220,n30221 );
   not U28350 ( p3_u2915,n26904 );
   and U28351 ( n26906,n40088,n40089 );
   not U28352 ( p2_u2989,n26906 );
   and U28353 ( n26908,n39418,n39419 );
   not U28354 ( p2_u3016,n26908 );
   and U28355 ( n26910,n30273,n30274 );
   not U28356 ( p3_u2909,n26910 );
   and U28357 ( n26912,n45752,n45753 );
   not U28358 ( p1_u3163,n26912 );
   and U28359 ( n26914,n48829,n48830 );
   not U28360 ( p1_u2968,n26914 );
   and U28361 ( n26916,n31478,n31479 );
   not U28362 ( p3_u2838,n26916 );
   and U28363 ( n26918,n31405,n31406 );
   not U28364 ( p3_u2840,n26918 );
   and U28365 ( n26920,n46828,n46829 );
   not U28366 ( p1_u3076,n26920 );
   and U28367 ( n26922,n46804,n46805 );
   not U28368 ( p1_u3079,n26922 );
   and U28369 ( n26924,n38717,n38718 );
   not U28370 ( p2_u3046,n26924 );
   and U28371 ( n26926,n30233,n30234 );
   not U28372 ( p3_u2914,n26926 );
   and U28373 ( n26928,n31590,n31591 );
   not U28374 ( p3_u2835,n26928 );
   and U28375 ( n26930,n30257,n30258 );
   not U28376 ( p3_u2911,n26930 );
   and U28377 ( n26932,n46844,n46845 );
   not U28378 ( p1_u3074,n26932 );
   and U28379 ( n26934,n46112,n46113 );
   not U28380 ( p1_u3143,n26934 );
   and U28381 ( n26936,n48306,n48307 );
   not U28382 ( p1_u2998,n26936 );
   and U28383 ( n26938,n46128,n46129 );
   not U28384 ( p1_u3141,n26938 );
   and U28385 ( n26940,n38900,n38901 );
   not U28386 ( p2_u3038,n26940 );
   and U28387 ( n26942,n46160,n46161 );
   not U28388 ( p1_u3137,n26942 );
   and U28389 ( n26944,n40063,n40064 );
   not U28390 ( p2_u2990,n26944 );
   and U28391 ( n26946,n46136,n46137 );
   not U28392 ( p1_u3140,n26946 );
   and U28393 ( n26948,n40130,n40131 );
   not U28394 ( p2_u2987,n26948 );
   and U28395 ( n26950,n46099,n46100 );
   not U28396 ( p1_u3144,n26950 );
   and U28397 ( n26952,n46812,n46813 );
   not U28398 ( p1_u3078,n26952 );
   and U28399 ( n26954,n40166,n40167 );
   not U28400 ( p2_u2985,n26954 );
   and U28401 ( n26956,n39759,n39760 );
   not U28402 ( p2_u3005,n26956 );
   and U28403 ( n26958,n40001,n40002 );
   not U28404 ( p2_u2993,n26958 );
   and U28405 ( n26960,n39881,n39882 );
   not U28406 ( p2_u2999,n26960 );
   and U28407 ( n26962,n46852,n46853 );
   not U28408 ( p1_u3073,n26962 );
   and U28409 ( n26964,n39982,n39983 );
   not U28410 ( p2_u2994,n26964 );
   and U28411 ( n26966,n46144,n46145 );
   not U28412 ( p1_u3139,n26966 );
   and U28413 ( n26968,n46152,n46153 );
   not U28414 ( p1_u3138,n26968 );
   and U28415 ( n26970,n39093,n39094 );
   not U28416 ( p2_u3030,n26970 );
   and U28417 ( n26972,n31934,n31935 );
   not U28418 ( p3_u2829,n26972 );
   and U28419 ( n26974,n46836,n46837 );
   not U28420 ( p1_u3075,n26974 );
   and U28421 ( n26976,n46791,n46792 );
   not U28422 ( p1_u3080,n26976 );
   and U28423 ( n26978,n39122,n39123 );
   not U28424 ( p2_u3029,n26978 );
   and U28425 ( n26980,n39141,n39142 );
   not U28426 ( p2_u3028,n26980 );
   and U28427 ( n26982,n46820,n46821 );
   not U28428 ( p1_u3077,n26982 );
   and U28429 ( n26984,n39170,n39171 );
   not U28430 ( p2_u3027,n26984 );
   and U28431 ( n26986,n46120,n46121 );
   not U28432 ( p1_u3142,n26986 );
   and U28433 ( n26988,n39861,n39862 );
   not U28434 ( p2_u3000,n26988 );
   and U28435 ( n26990,n32247,n32248 );
   not U28436 ( p3_u2818,n26990 );
   and U28437 ( n26992,n35591,n35592 );
   not U28438 ( p3_u2662,n26992 );
   and U28439 ( n26994,n35643,n35644 );
   not U28440 ( p3_u2660,n26994 );
   and U28441 ( n26996,n38343,n38344 );
   not U28442 ( p2_u3073,n26996 );
   and U28443 ( n26998,n35426,n35427 );
   not U28444 ( p3_u2668,n26998 );
   and U28445 ( n27000,n38351,n38352 );
   not U28446 ( p2_u3072,n27000 );
   and U28447 ( n27002,n39701,n39702 );
   not U28448 ( p2_u3008,n27002 );
   and U28449 ( n27004,n38319,n38320 );
   not U28450 ( p2_u3076,n27004 );
   and U28451 ( n27006,n38327,n38328 );
   not U28452 ( p2_u3075,n27006 );
   and U28453 ( n27008,n38303,n38304 );
   not U28454 ( p2_u3078,n27008 );
   and U28455 ( n27010,n38311,n38312 );
   not U28456 ( p2_u3077,n27010 );
   and U28457 ( n27012,n38290,n38291 );
   not U28458 ( p2_u3079,n27012 );
   and U28459 ( n27014,n38335,n38336 );
   not U28460 ( p2_u3074,n27014 );
   and U28461 ( n27016,n45922,n45923 );
   not U28462 ( p1_u3157,n27016 );
   and U28463 ( n27018,n45910,n45911 );
   not U28464 ( p1_u3158,n27018 );
   and U28465 ( n27020,n46972,n46973 );
   not U28466 ( p1_u3063,n27020 );
   and U28467 ( n27022,n46996,n46997 );
   not U28468 ( p1_u3060,n27022 );
   and U28469 ( n27024,n45934,n45935 );
   not U28470 ( p1_u3156,n27024 );
   and U28471 ( n27026,n45958,n45959 );
   not U28472 ( p1_u3154,n27026 );
   and U28473 ( n27028,n46988,n46989 );
   not U28474 ( p1_u3061,n27028 );
   and U28475 ( n27030,n47020,n47021 );
   not U28476 ( p1_u3057,n27030 );
   and U28477 ( n27032,n45881,n45882 );
   not U28478 ( p1_u3160,n27032 );
   and U28479 ( n27034,n45946,n45947 );
   not U28480 ( p1_u3155,n27034 );
   and U28481 ( n27036,n46959,n46960 );
   not U28482 ( p1_u3064,n27036 );
   and U28483 ( n27038,n45898,n45899 );
   not U28484 ( p1_u3159,n27038 );
   and U28485 ( n27040,n38398,n38399 );
   not U28486 ( p2_u3069,n27040 );
   and U28487 ( n27042,n47004,n47005 );
   not U28488 ( p1_u3059,n27042 );
   and U28489 ( n27044,n47012,n47013 );
   not U28490 ( p1_u3058,n27044 );
   and U28491 ( n27046,n31616,n31617 );
   not U28492 ( p3_u2834,n27046 );
   and U28493 ( n27048,n46980,n46981 );
   not U28494 ( p1_u3062,n27048 );
   and U28495 ( n27050,n45970,n45971 );
   not U28496 ( p1_u3153,n27050 );
   and U28497 ( n27052,n38422,n38423 );
   not U28498 ( p2_u3066,n27052 );
   and U28499 ( n27054,n38406,n38407 );
   not U28500 ( p2_u3068,n27054 );
   and U28501 ( n27056,n38438,n38439 );
   not U28502 ( p2_u3064,n27056 );
   and U28503 ( n27058,n38430,n38431 );
   not U28504 ( p2_u3065,n27058 );
   and U28505 ( n27060,n38414,n38415 );
   not U28506 ( p2_u3067,n27060 );
   and U28507 ( n27062,n38390,n38391 );
   not U28508 ( p2_u3070,n27062 );
   and U28509 ( n27064,n38377,n38378 );
   not U28510 ( p2_u3071,n27064 );
   and U28511 ( n27066,n47263,n47264 );
   not U28512 ( p1_u3038,n27066 );
   and U28513 ( n27068,n47247,n47248 );
   not U28514 ( p1_u3039,n27068 );
   and U28515 ( n27070,n47047,n47048 );
   not U28516 ( p1_u3056,n27070 );
   and U28517 ( n27072,n47295,n47296 );
   not U28518 ( p1_u3036,n27072 );
   and U28519 ( n27074,n47223,n47224 );
   not U28520 ( p1_u3040,n27074 );
   and U28521 ( n27076,n47145,n47146 );
   not U28522 ( p1_u3047,n27076 );
   and U28523 ( n27078,n47131,n47132 );
   not U28524 ( p1_u3048,n27078 );
   and U28525 ( n27080,n47060,n47061 );
   not U28526 ( p1_u3055,n27080 );
   and U28527 ( n27082,n47076,n47077 );
   not U28528 ( p1_u3053,n27082 );
   and U28529 ( n27084,n47108,n47109 );
   not U28530 ( p1_u3049,n27084 );
   and U28531 ( n27086,n39943,n39944 );
   not U28532 ( p2_u2996,n27086 );
   and U28533 ( n27088,n40105,n40106 );
   not U28534 ( p2_u2988,n27088 );
   and U28535 ( n27090,n40045,n40046 );
   not U28536 ( p2_u2991,n27090 );
   and U28537 ( n27092,n47181,n47182 );
   not U28538 ( p1_u3043,n27092 );
   and U28539 ( n27094,n47311,n47312 );
   not U28540 ( p1_u3035,n27094 );
   and U28541 ( n27096,n39740,n39741 );
   not U28542 ( p2_u3006,n27096 );
   and U28543 ( n27098,n47092,n47093 );
   not U28544 ( p1_u3051,n27098 );
   and U28545 ( n27100,n47342,n47343 );
   not U28546 ( p1_u3033,n27100 );
   and U28547 ( n27102,n47154,n47155 );
   not U28548 ( p1_u3046,n27102 );
   and U28549 ( n27104,n47326,n47327 );
   not U28550 ( p1_u3034,n27104 );
   and U28551 ( n27106,n47279,n47280 );
   not U28552 ( p1_u3037,n27106 );
   and U28553 ( n27108,n47190,n47191 );
   not U28554 ( p1_u3042,n27108 );
   and U28555 ( n27110,n47068,n47069 );
   not U28556 ( p1_u3054,n27110 );
   and U28557 ( n27112,n47084,n47085 );
   not U28558 ( p1_u3052,n27112 );
   and U28559 ( n27114,n39797,n39798 );
   not U28560 ( p2_u3003,n27114 );
   and U28561 ( n27116,n37865,n37866 );
   not U28562 ( p2_u3119,n27116 );
   and U28563 ( n27118,n32117,n32118 );
   not U28564 ( p3_u2823,n27118 );
   and U28565 ( n27120,n39926,n39927 );
   not U28566 ( p2_u2997,n27120 );
   and U28567 ( n27122,n47100,n47101 );
   not U28568 ( p1_u3050,n27122 );
   and U28569 ( n27124,n47199,n47200 );
   not U28570 ( p1_u3041,n27124 );
   and U28571 ( n27126,n39681,n39682 );
   not U28572 ( p2_u3009,n27126 );
   and U28573 ( n27128,n48743,n48744 );
   not U28574 ( p1_u2972,n27128 );
   and U28575 ( n27130,n47172,n47173 );
   not U28576 ( p1_u3044,n27130 );
   and U28577 ( n27132,n47163,n47164 );
   not U28578 ( p1_u3045,n27132 );
   and U28579 ( n27134,n37878,n37879 );
   not U28580 ( p2_u3118,n27134 );
   and U28581 ( n27136,n37926,n37927 );
   not U28582 ( p2_u3112,n27136 );
   and U28583 ( n27138,n37918,n37919 );
   not U28584 ( p2_u3113,n27138 );
   and U28585 ( n27140,n37894,n37895 );
   not U28586 ( p2_u3116,n27140 );
   and U28587 ( n27142,n37910,n37911 );
   not U28588 ( p2_u3114,n27142 );
   and U28589 ( n27144,n37902,n37903 );
   not U28590 ( p2_u3115,n27144 );
   and U28591 ( n27146,n39816,n39817 );
   not U28592 ( p2_u3002,n27146 );
   and U28593 ( n27148,n38609,n38610 );
   not U28594 ( p2_u3052,n27148 );
   and U28595 ( n27150,n38577,n38578 );
   not U28596 ( p2_u3054,n27150 );
   and U28597 ( n27152,n38641,n38642 );
   not U28598 ( p2_u3050,n27152 );
   and U28599 ( n27154,n38593,n38594 );
   not U28600 ( p2_u3053,n27154 );
   and U28601 ( n27156,n38528,n38529 );
   not U28602 ( p2_u3056,n27156 );
   and U28603 ( n27158,n37886,n37887 );
   not U28604 ( p2_u3117,n27158 );
   and U28605 ( n27160,n38519,n38520 );
   not U28606 ( p2_u3057,n27160 );
   and U28607 ( n27162,n38657,n38658 );
   not U28608 ( p2_u3049,n27162 );
   and U28609 ( n27164,n38501,n38502 );
   not U28610 ( p2_u3059,n27164 );
   and U28611 ( n27166,n38483,n38484 );
   not U28612 ( p2_u3061,n27166 );
   and U28613 ( n27168,n38510,n38511 );
   not U28614 ( p2_u3058,n27168 );
   and U28615 ( n27170,n38552,n38553 );
   not U28616 ( p2_u3055,n27170 );
   and U28617 ( n27172,n38672,n38673 );
   not U28618 ( p2_u3048,n27172 );
   and U28619 ( n27174,n38492,n38493 );
   not U28620 ( p2_u3060,n27174 );
   and U28621 ( n27176,n49592,n49593 );
   not U28622 ( p1_u2874,n27176 );
   and U28623 ( n27178,n49460,n49461 );
   not U28624 ( p1_u2886,n27178 );
   and U28625 ( n27180,n49449,n49450 );
   not U28626 ( p1_u2887,n27180 );
   and U28627 ( n27182,n38625,n38626 );
   not U28628 ( p2_u3051,n27182 );
   and U28629 ( n27184,n32226,n32227 );
   not U28630 ( p3_u2819,n27184 );
   and U28631 ( n27186,n49471,n49472 );
   not U28632 ( p1_u2885,n27186 );
   and U28633 ( n27188,n31088,n31089 );
   not U28634 ( p3_u2851,n27188 );
   and U28635 ( n27190,n35362,n35363 );
   not U28636 ( p3_u2671,n27190 );
   and U28637 ( n27192,n38474,n38475 );
   not U28638 ( p2_u3062,n27192 );
   and U28639 ( n27194,n38460,n38461 );
   not U28640 ( p2_u3063,n27194 );
   and U28641 ( n27196,n38064,n38065 );
   not U28642 ( p2_u3100,n27196 );
   and U28643 ( n27198,n38048,n38049 );
   not U28644 ( p2_u3102,n27198 );
   and U28645 ( n27200,n38080,n38081 );
   not U28646 ( p2_u3098,n27200 );
   and U28647 ( n27202,n38072,n38073 );
   not U28648 ( p2_u3099,n27202 );
   and U28649 ( n27204,n38056,n38057 );
   not U28650 ( p2_u3101,n27204 );
   and U28651 ( n27206,n38035,n38036 );
   not U28652 ( p2_u3103,n27206 );
   and U28653 ( n27208,n46223,n46224 );
   not U28654 ( p1_u3132,n27208 );
   and U28655 ( n27210,n38088,n38089 );
   not U28656 ( p2_u3097,n27210 );
   and U28657 ( n27212,n32488,n32489 );
   not U28658 ( p3_u2811,n27212 );
   and U28659 ( n27214,n46215,n46216 );
   not U28660 ( p1_u3133,n27214 );
   and U28661 ( n27216,n46247,n46248 );
   not U28662 ( p1_u3129,n27216 );
   and U28663 ( n27218,n46912,n46913 );
   not U28664 ( p1_u3068,n27218 );
   and U28665 ( n27220,n46207,n46208 );
   not U28666 ( p1_u3134,n27220 );
   and U28667 ( n27222,n38096,n38097 );
   not U28668 ( p2_u3096,n27222 );
   and U28669 ( n27224,n46199,n46200 );
   not U28670 ( p1_u3135,n27224 );
   and U28671 ( n27226,n46920,n46921 );
   not U28672 ( p1_u3067,n27226 );
   and U28673 ( n27228,n46875,n46876 );
   not U28674 ( p1_u3072,n27228 );
   and U28675 ( n27230,n37368,n37369 );
   not U28676 ( p2_u3165,n27230 );
   and U28677 ( n27232,n37360,n37361 );
   not U28678 ( p2_u3166,n27232 );
   and U28679 ( n27234,n46186,n46187 );
   not U28680 ( p1_u3136,n27234 );
   and U28681 ( n27236,n33409,n33410 );
   not U28682 ( p3_u2735,n27236 );
   and U28683 ( n27238,n31948,n31949 );
   not U28684 ( p3_u2828,n27238 );
   and U28685 ( n27240,n32698,n32699 );
   not U28686 ( p3_u2805,n27240 );
   and U28687 ( n27242,n37347,n37348 );
   not U28688 ( p2_u3167,n27242 );
   and U28689 ( n27244,n46888,n46889 );
   not U28690 ( p1_u3071,n27244 );
   and U28691 ( n27246,n46231,n46232 );
   not U28692 ( p1_u3131,n27246 );
   and U28693 ( n27248,n46239,n46240 );
   not U28694 ( p1_u3130,n27248 );
   and U28695 ( n27250,n46896,n46897 );
   not U28696 ( p1_u3070,n27250 );
   and U28697 ( n27252,n46936,n46937 );
   not U28698 ( p1_u3065,n27252 );
   and U28699 ( n27254,n32357,n32358 );
   not U28700 ( p3_u2815,n27254 );
   and U28701 ( n27256,n37400,n37401 );
   not U28702 ( p2_u3161,n27256 );
   and U28703 ( n27258,n46904,n46905 );
   not U28704 ( p1_u3069,n27258 );
   and U28705 ( n27260,n37384,n37385 );
   not U28706 ( p2_u3163,n27260 );
   and U28707 ( n27262,n37392,n37393 );
   not U28708 ( p2_u3162,n27262 );
   and U28709 ( n27264,n37408,n37409 );
   not U28710 ( p2_u3160,n27264 );
   and U28711 ( n27266,n35380,n35381 );
   not U28712 ( p3_u2670,n27266 );
   and U28713 ( n27268,n38002,n38003 );
   not U28714 ( p2_u3105,n27268 );
   and U28715 ( n27270,n37994,n37995 );
   not U28716 ( p2_u3106,n27270 );
   and U28717 ( n27272,n38124,n38125 );
   not U28718 ( p2_u3095,n27272 );
   and U28719 ( n27274,n38010,n38011 );
   not U28720 ( p2_u3104,n27274 );
   and U28721 ( n27276,n46928,n46929 );
   not U28722 ( p1_u3066,n27276 );
   and U28723 ( n27278,n37376,n37377 );
   not U28724 ( p2_u3164,n27278 );
   and U28725 ( n27280,n37970,n37971 );
   not U28726 ( p2_u3109,n27280 );
   and U28727 ( n27282,n38137,n38138 );
   not U28728 ( p2_u3094,n27282 );
   and U28729 ( n27284,n37949,n37950 );
   not U28730 ( p2_u3111,n27284 );
   and U28731 ( n27286,n37962,n37963 );
   not U28732 ( p2_u3110,n27286 );
   and U28733 ( n27288,n37978,n37979 );
   not U28734 ( p2_u3108,n27288 );
   and U28735 ( n27290,n37986,n37987 );
   not U28736 ( p2_u3107,n27290 );
   and U28737 ( n27292,n38161,n38162 );
   not U28738 ( p2_u3091,n27292 );
   and U28739 ( n27294,n38145,n38146 );
   not U28740 ( p2_u3093,n27294 );
   and U28741 ( n27296,n38177,n38178 );
   not U28742 ( p2_u3089,n27296 );
   and U28743 ( n27298,n38169,n38170 );
   not U28744 ( p2_u3090,n27298 );
   and U28745 ( n27300,n38153,n38154 );
   not U28746 ( p2_u3092,n27300 );
   and U28747 ( n27302,n46678,n46679 );
   not U28748 ( p1_u3089,n27302 );
   and U28749 ( n27304,n46662,n46663 );
   not U28750 ( p1_u3091,n27304 );
   and U28751 ( n27306,n38185,n38186 );
   not U28752 ( p2_u3088,n27306 );
   and U28753 ( n27308,n46670,n46671 );
   not U28754 ( p1_u3090,n27308 );
   and U28755 ( n27310,n46617,n46618 );
   not U28756 ( p1_u3096,n27310 );
   and U28757 ( n27312,n46654,n46655 );
   not U28758 ( p1_u3092,n27312 );
   and U28759 ( n27314,n46646,n46647 );
   not U28760 ( p1_u3093,n27314 );
   and U28761 ( n27316,n38228,n38229 );
   not U28762 ( p2_u3085,n27316 );
   and U28763 ( n27318,n38207,n38208 );
   not U28764 ( p2_u3087,n27318 );
   and U28765 ( n27320,n38244,n38245 );
   not U28766 ( p2_u3083,n27320 );
   and U28767 ( n27322,n38236,n38237 );
   not U28768 ( p2_u3084,n27322 );
   and U28769 ( n27324,n38220,n38221 );
   not U28770 ( p2_u3086,n27324 );
   and U28771 ( n27326,n46630,n46631 );
   not U28772 ( p1_u3095,n27326 );
   and U28773 ( n27328,n45693,n45694 );
   not U28774 ( p1_u3195,n27328 );
   and U28775 ( n27330,n29084,n29085 );
   not U28776 ( p3_u3030,n27330 );
   and U28777 ( n27332,n38252,n38253 );
   not U28778 ( p2_u3082,n27332 );
   and U28779 ( n27334,n38268,n38269 );
   not U28780 ( p2_u3080,n27334 );
   and U28781 ( n27336,n38260,n38261 );
   not U28782 ( p2_u3081,n27336 );
   and U28783 ( n27338,n46638,n46639 );
   not U28784 ( p1_u3094,n27338 );
   and U28785 ( n27340,n41384,n41385 );
   not U28786 ( p2_u2900,n27340 );
   and U28787 ( n27342,n34039,n34040 );
   not U28788 ( p3_u2715,n27342 );
   and U28789 ( n27344,n37435,n37436 );
   not U28790 ( p2_u3159,n27344 );
   and U28791 ( n27346,n41352,n41353 );
   not U28792 ( p2_u2902,n27346 );
   and U28793 ( n27348,n41560,n41561 );
   not U28794 ( p2_u2889,n27348 );
   and U28795 ( n27350,n34069,n34070 );
   not U28796 ( p3_u2713,n27350 );
   and U28797 ( n27352,n34026,n34027 );
   not U28798 ( p3_u2716,n27352 );
   and U28799 ( n27354,n37448,n37449 );
   not U28800 ( p2_u3158,n27354 );
   and U28801 ( n27356,n34010,n34011 );
   not U28802 ( p3_u2717,n27356 );
   and U28803 ( n27358,n33979,n33980 );
   not U28804 ( p3_u2719,n27358 );
   and U28805 ( n27360,n41368,n41369 );
   not U28806 ( p2_u2901,n27360 );
   and U28807 ( n27362,n37456,n37457 );
   not U28808 ( p2_u3157,n27362 );
   and U28809 ( n27364,n37472,n37473 );
   not U28810 ( p2_u3155,n27364 );
   and U28811 ( n27366,n34056,n34057 );
   not U28812 ( p3_u2714,n27366 );
   and U28813 ( n27368,n37488,n37489 );
   not U28814 ( p2_u3153,n27368 );
   and U28815 ( n27370,n37480,n37481 );
   not U28816 ( p2_u3154,n27370 );
   and U28817 ( n27372,n37464,n37465 );
   not U28818 ( p2_u3156,n27372 );
   and U28819 ( n27374,n33997,n33998 );
   not U28820 ( p3_u2718,n27374 );
   and U28821 ( n27376,n33968,n33969 );
   not U28822 ( p3_u2720,n27376 );
   and U28823 ( n27378,n32797,n32798 );
   not U28824 ( p3_u2802,n27378 );
   and U28825 ( n27380,n33879,n33880 );
   not U28826 ( p3_u2727,n27380 );
   and U28827 ( n27382,n31280,n31281 );
   not U28828 ( p3_u2844,n27382 );
   and U28829 ( n27384,n34098,n34099 );
   not U28830 ( p3_u2711,n27384 );
   and U28831 ( n27386,n37496,n37497 );
   not U28832 ( p2_u3152,n27386 );
   and U28833 ( n27388,n50404,n50405 );
   not U28834 ( p1_u2817,n27388 );
   and U28835 ( n27390,n33904,n33905 );
   not U28836 ( p3_u2725,n27390 );
   and U28837 ( n27392,n50425,n50426 );
   not U28838 ( p1_u2816,n27392 );
   and U28839 ( n27394,n47801,n47802 );
   not U28840 ( p1_u3016,n27394 );
   and U28841 ( n27396,n36990,n36991 );
   not U28842 ( p2_u3209,n27396 );
   and U28843 ( n27398,n33929,n33930 );
   not U28844 ( p3_u2723,n27398 );
   and U28845 ( n27400,n32167,n32168 );
   not U28846 ( p3_u2821,n27400 );
   and U28847 ( n27402,n50377,n50378 );
   not U28848 ( p1_u2818,n27402 );
   and U28849 ( n27404,n33756,n33757 );
   not U28850 ( p3_u2729,n27404 );
   and U28851 ( n27406,n32014,n32015 );
   not U28852 ( p3_u2826,n27406 );
   and U28853 ( n27408,n29162,n29163 );
   not U28854 ( p3_u2996,n27408 );
   and U28855 ( n27410,n50516,n50517 );
   not U28856 ( p1_u2812,n27410 );
   and U28857 ( n27412,n50333,n50334 );
   not U28858 ( p1_u2820,n27412 );
   and U28859 ( n27414,n34186,n34187 );
   not U28860 ( p3_u2705,n27414 );
   and U28861 ( n27416,n47707,n47708 );
   not U28862 ( p1_u3020,n27416 );
   and U28863 ( n27418,n50538,n50539 );
   not U28864 ( p1_u2811,n27418 );
   and U28865 ( n27420,n50555,n50556 );
   not U28866 ( p1_u2810,n27420 );
   and U28867 ( n27422,n32888,n32889 );
   not U28868 ( p3_u2799,n27422 );
   and U28869 ( n27424,n33954,n33955 );
   not U28870 ( p3_u2721,n27424 );
   and U28871 ( n27426,n50494,n50495 );
   not U28872 ( p1_u2813,n27426 );
   and U28873 ( n27428,n33645,n33646 );
   not U28874 ( p3_u2731,n27428 );
   and U28875 ( n27430,n32192,n32193 );
   not U28876 ( p3_u2820,n27430 );
   and U28877 ( n27432,n33535,n33536 );
   not U28878 ( p3_u2733,n27432 );
   and U28879 ( n27434,n39583,n39584 );
   not U28880 ( p2_u3014,n27434 );
   and U28881 ( n27436,n47568,n47569 );
   not U28882 ( p1_u3026,n27436 );
   and U28883 ( n27438,n45773,n45774 );
   not U28884 ( p1_u3161,n27438 );
   and U28885 ( n27440,n31347,n31348 );
   not U28886 ( p3_u2842,n27440 );
   and U28887 ( n27442,n37047,n37048 );
   not U28888 ( p2_u3176,n27442 );
   and U28889 ( n27444,n31972,n31973 );
   not U28890 ( p3_u2827,n27444 );
   and U28891 ( n27446,n34143,n34144 );
   not U28892 ( p3_u2708,n27446 );
   and U28893 ( n27448,n34114,n34115 );
   not U28894 ( p3_u2710,n27448 );
   and U28895 ( n27450,n48290,n48291 );
   not U28896 ( p1_u2999,n27450 );
   and U28897 ( n27452,n48151,n48152 );
   not U28898 ( p1_u3000,n27452 );
   and U28899 ( n27454,n31201,n31202 );
   not U28900 ( p3_u2847,n27454 );
   and U28901 ( n27456,n30986,n30987 );
   not U28902 ( p3_u2855,n27456 );
   and U28903 ( n27458,n47461,n47462 );
   not U28904 ( p1_u3031,n27458 );
   and U28905 ( n27460,n34128,n34129 );
   not U28906 ( p3_u2709,n27460 );
   and U28907 ( n27462,n34157,n34158 );
   not U28908 ( p3_u2707,n27462 );
   and U28909 ( n27464,n31008,n31009 );
   not U28910 ( p3_u2854,n27464 );
   and U28911 ( n27466,n31229,n31230 );
   not U28912 ( p3_u2846,n27466 );
   and U28913 ( n27468,n47542,n47543 );
   not U28914 ( p1_u3027,n27468 );
   and U28915 ( n27470,n31165,n31166 );
   not U28916 ( p3_u2848,n27470 );
   and U28917 ( n27472,n28483,n28484 );
   not U28918 ( u281,n27472 );
   and U28919 ( n27474,n28525,n28526 );
   not U28920 ( u260,n27474 );
   and U28921 ( n27476,n28521,n28522 );
   not U28922 ( u262,n27476 );
   and U28923 ( n27478,n34169,n34170 );
   not U28924 ( p3_u2706,n27478 );
   and U28925 ( n27480,n34085,n34086 );
   not U28926 ( p3_u2712,n27480 );
   and U28927 ( n27482,n30843,n30844 );
   not U28928 ( p3_u2860,n27482 );
   and U28929 ( n27484,n28537,n28538 );
   not U28930 ( u254,n27484 );
   and U28931 ( n27486,n28511,n28512 );
   not U28932 ( u267,n27486 );
   and U28933 ( n27488,n28513,n28514 );
   not U28934 ( u266,n27488 );
   and U28935 ( n27490,n28480,n28481 );
   not U28936 ( u282,n27490 );
   and U28937 ( n27492,n28505,n28506 );
   not U28938 ( u270,n27492 );
   and U28939 ( n27494,n28529,n28530 );
   not U28940 ( u258,n27494 );
   and U28941 ( n27496,n28535,n28536 );
   not U28942 ( u255,n27496 );
   and U28943 ( n27498,n28541,n28542 );
   not U28944 ( u252,n27498 );
   and U28945 ( n27500,n28539,n28540 );
   not U28946 ( u253,n27500 );
   and U28947 ( n27502,n28543,n28544 );
   not U28948 ( u251,n27502 );
   and U28949 ( n27504,n28501,n28502 );
   not U28950 ( u272,n27504 );
   and U28951 ( n27506,n28531,n28532 );
   not U28952 ( u257,n27506 );
   and U28953 ( n27508,n28509,n28510 );
   not U28954 ( u268,n27508 );
   and U28955 ( n27510,n28487,n28488 );
   not U28956 ( u279,n27510 );
   and U28957 ( n27512,n28507,n28508 );
   not U28958 ( u269,n27512 );
   and U28959 ( n27514,n28519,n28520 );
   not U28960 ( u263,n27514 );
   and U28961 ( n27516,n28523,n28524 );
   not U28962 ( u261,n27516 );
   and U28963 ( n27518,n28491,n28492 );
   not U28964 ( u277,n27518 );
   and U28965 ( n27520,n28485,n28486 );
   not U28966 ( u280,n27520 );
   and U28967 ( n27522,n28503,n28504 );
   not U28968 ( u271,n27522 );
   and U28969 ( n27524,n28497,n28498 );
   not U28970 ( u274,n27524 );
   and U28971 ( n27526,n28493,n28494 );
   not U28972 ( u276,n27526 );
   and U28973 ( n27528,n28489,n28490 );
   not U28974 ( u278,n27528 );
   and U28975 ( n27530,n28495,n28496 );
   not U28976 ( u275,n27530 );
   and U28977 ( n27532,n34239,n34240 );
   not U28978 ( p3_u2702,n27532 );
   and U28979 ( n27534,n28499,n28500 );
   not U28980 ( u273,n27534 );
   and U28981 ( n27536,n28533,n28534 );
   not U28982 ( u256,n27536 );
   and U28983 ( n27538,n28515,n28516 );
   not U28984 ( u265,n27538 );
   and U28985 ( n27540,n28527,n28528 );
   not U28986 ( u259,n27540 );
   and U28987 ( n27542,n28517,n28518 );
   not U28988 ( u264,n27542 );
   and U28989 ( n27544,n47914,n47915 );
   not U28990 ( p1_u3011,n27544 );
   and U28991 ( n27546,n47634,n47635 );
   not U28992 ( p1_u3023,n27546 );
   and U28993 ( n27548,n48052,n48053 );
   not U28994 ( p1_u3005,n27548 );
   and U28995 ( n27550,n48006,n48007 );
   not U28996 ( p1_u3007,n27550 );
   and U28997 ( n27552,n48138,n48139 );
   not U28998 ( p1_u3001,n27552 );
   and U28999 ( n27554,n47680,n47681 );
   not U29000 ( p1_u3021,n27554 );
   and U29001 ( n27556,n47960,n47961 );
   not U29002 ( p1_u3009,n27556 );
   and U29003 ( n27558,n47728,n47729 );
   not U29004 ( p1_u3019,n27558 );
   and U29005 ( n27560,n47755,n47756 );
   not U29006 ( p1_u3018,n27560 );
   and U29007 ( n27562,n47822,n47823 );
   not U29008 ( p1_u3015,n27562 );
   and U29009 ( n27564,n47895,n47896 );
   not U29010 ( p1_u3012,n27564 );
   and U29011 ( n27566,n47941,n47942 );
   not U29012 ( p1_u3010,n27566 );
   and U29013 ( n27568,n33813,n33814 );
   not U29014 ( p3_u2728,n27568 );
   and U29015 ( n27570,n33918,n33919 );
   not U29016 ( p3_u2724,n27570 );
   and U29017 ( n27572,n33702,n33703 );
   not U29018 ( p3_u2730,n27572 );
   and U29019 ( n27574,n47661,n47662 );
   not U29020 ( p1_u3022,n27574 );
   and U29021 ( n27576,n48101,n48102 );
   not U29022 ( p1_u3003,n27576 );
   and U29023 ( n27578,n48033,n48034 );
   not U29024 ( p1_u3006,n27578 );
   and U29025 ( n27580,n29151,n29152 );
   not U29026 ( p3_u2997,n27580 );
   and U29027 ( n27582,n31688,n31689 );
   not U29028 ( p3_u2832,n27582 );
   and U29029 ( n27584,n33943,n33944 );
   not U29030 ( p3_u2722,n27584 );
   and U29031 ( n27586,n33893,n33894 );
   not U29032 ( p3_u2726,n27586 );
   and U29033 ( n27588,n33591,n33592 );
   not U29034 ( p3_u2732,n27588 );
   and U29035 ( n27590,n33481,n33482 );
   not U29036 ( p3_u2734,n27590 );
   and U29037 ( n27592,n36675,n36676 );
   not U29038 ( p2_u3604,n27592 );
   and U29039 ( n27594,n36663,n36664 );
   not U29040 ( p2_u3605,n27594 );
   and U29041 ( n27596,n28868,n28869 );
   not U29042 ( p3_u3285,n27596 );
   and U29043 ( n27598,n28857,n28858 );
   not U29044 ( p3_u3288,n27598 );
   and U29045 ( n27600,n28832,n28833 );
   not U29046 ( p3_u3290,n27600 );
   and U29047 ( n27602,n28844,n28845 );
   not U29048 ( p3_u3289,n27602 );
   and U29049 ( n27604,n45395,n45396 );
   not U29050 ( p1_u3477,n27604 );
   and U29051 ( n27606,n45409,n45410 );
   not U29052 ( p1_u3476,n27606 );
   and U29053 ( n27608,n45382,n45383 );
   not U29054 ( p1_u3478,n27608 );
   and U29055 ( n27610,n45423,n45424 );
   not U29056 ( p1_u3475,n27610 );
   and U29057 ( n27612,n36689,n36690 );
   not U29058 ( p2_u3603,n27612 );
   and U29059 ( n27614,n36703,n36704 );
   not U29060 ( p2_u3602,n27614 );
   and U29061 ( n27616,n28463,n28464 );
   not U29062 ( u351,n27616 );
   and U29063 ( n27618,n28469,n28470 );
   not U29064 ( u348,n27618 );
   and U29065 ( n27620,n28415,n28416 );
   not U29066 ( u375,n27620 );
   and U29067 ( n27622,n28467,n28468 );
   not U29068 ( u349,n27622 );
   and U29069 ( n27624,n28411,n28412 );
   not U29070 ( u376,n27624 );
   and U29071 ( n27626,n28471,n28472 );
   not U29072 ( u347,n27626 );
   and U29073 ( n27628,n45454,n45455 );
   not U29074 ( p1_u3473,n27628 );
   and U29075 ( n27630,n36766,n36767 );
   not U29076 ( p2_u3596,n27630 );
   and U29077 ( n27632,n36747,n36748 );
   not U29078 ( p2_u3599,n27632 );
   and U29079 ( n27634,n28459,n28460 );
   not U29080 ( u353,n27634 );
   and U29081 ( n27636,n28465,n28466 );
   not U29082 ( u350,n27636 );
   and U29083 ( n27638,n28461,n28462 );
   not U29084 ( u352,n27638 );
   and U29085 ( n27640,n33394,n33395 );
   not U29086 ( p3_u2738,n27640 );
   and U29087 ( n27642,n33384,n33385 );
   not U29088 ( p3_u2740,n27642 );
   and U29089 ( n27644,n33389,n33390 );
   not U29090 ( p3_u2739,n27644 );
   and U29091 ( n27646,n45482,n45483 );
   not U29092 ( p1_u3469,n27646 );
   and U29093 ( n27648,n36734,n36735 );
   not U29094 ( p2_u3600,n27648 );
   and U29095 ( n27650,n45467,n45468 );
   not U29096 ( p1_u3472,n27650 );
   and U29097 ( n27652,n28816,n28817 );
   not U29098 ( p3_u3294,n27652 );
   and U29099 ( n27654,n33379,n33380 );
   not U29100 ( p3_u2741,n27654 );
   and U29101 ( n27656,n33374,n33375 );
   not U29102 ( p3_u2742,n27656 );
   and U29103 ( n27658,n33254,n33255 );
   not U29104 ( p3_u2766,n27658 );
   and U29105 ( n27660,n33369,n33370 );
   not U29106 ( p3_u2743,n27660 );
   and U29107 ( n27662,n33246,n33247 );
   not U29108 ( p3_u2767,n27662 );
   and U29109 ( n27664,n36610,n36611 );
   not U29110 ( p2_u3612,n27664 );
   and U29111 ( n27666,n45499,n45500 );
   not U29112 ( p1_u3466,n27666 );
   and U29113 ( n27668,n45334,n45335 );
   not U29114 ( p1_u3485,n27668 );
   and U29115 ( n27670,n28782,n28783 );
   not U29116 ( p3_u3296,n27670 );
   and U29117 ( n27672,n45366,n45367 );
   not U29118 ( p1_u3483,n27672 );
   and U29119 ( n27674,n36661,n36662 );
   not U29120 ( p2_u3608,n27674 );
   and U29121 ( n27676,n50093,n50094 );
   not U29122 ( p1_u2830,n27676 );
   and U29123 ( n27678,n50311,n50312 );
   not U29124 ( p1_u2821,n27678 );
   and U29125 ( n27680,n50070,n50071 );
   not U29126 ( p1_u2831,n27680 );
   and U29127 ( n27682,n45361,n45362 );
   not U29128 ( p1_u3484,n27682 );
   and U29129 ( n27684,n49020,n52729 );
   not U29130 ( p1_u2806,n27684 );
   and U29131 ( n27686,n36792,n36793 );
   not U29132 ( p2_u3592,n27686 );
   and U29133 ( n27688,n50192,n50193 );
   not U29134 ( p1_u2826,n27688 );
   and U29135 ( n27690,n50119,n50120 );
   not U29136 ( p1_u2829,n27690 );
   and U29137 ( n27692,n50219,n50220 );
   not U29138 ( p1_u2825,n27692 );
   and U29139 ( n27694,n49940,n49941 );
   not U29140 ( p1_u2836,n27694 );
   and U29141 ( n27696,n49971,n49972 );
   not U29142 ( p1_u2835,n27696 );
   and U29143 ( n27698,n49997,n49998 );
   not U29144 ( p1_u2834,n27698 );
   and U29145 ( n27700,n50265,n50266 );
   not U29146 ( p1_u2823,n27700 );
   and U29147 ( n27702,n50145,n50146 );
   not U29148 ( p1_u2828,n27702 );
   and U29149 ( n27704,n50169,n50170 );
   not U29150 ( p1_u2827,n27704 );
   and U29151 ( n27706,n50240,n50241 );
   not U29152 ( p1_u2824,n27706 );
   and U29153 ( n27708,n50288,n50289 );
   not U29154 ( p1_u2822,n27708 );
   and U29155 ( n27710,n50046,n50047 );
   not U29156 ( p1_u2832,n27710 );
   and U29157 ( n27712,n35771,n35772 );
   not U29158 ( p3_u2655,n27712 );
   and U29159 ( n27714,n35566,n35567 );
   not U29160 ( p3_u2663,n27714 );
   and U29161 ( n27716,n35822,n35823 );
   not U29162 ( p3_u2653,n27716 );
   and U29163 ( n27718,n48497,n48498 );
   not U29164 ( p1_u2986,n27718 );
   and U29165 ( n27720,n48428,n48429 );
   not U29166 ( p1_u2990,n27720 );
   and U29167 ( n27722,n50025,n50026 );
   not U29168 ( p1_u2833,n27722 );
   and U29169 ( n27724,n43030,n43031 );
   not U29170 ( p2_u2844,n27724 );
   and U29171 ( n27726,n35717,n35718 );
   not U29172 ( p3_u2657,n27726 );
   and U29173 ( n27728,n35618,n35619 );
   not U29174 ( p3_u2661,n27728 );
   and U29175 ( n27730,n35457,n35458 );
   not U29176 ( p3_u2667,n27730 );
   and U29177 ( n27732,n35669,n35670 );
   not U29178 ( p3_u2659,n27732 );
   and U29179 ( n27734,n35515,n35516 );
   not U29180 ( p3_u2665,n27734 );
   and U29181 ( n27736,n43205,n43206 );
   not U29182 ( p2_u2838,n27736 );
   and U29183 ( n27738,n43056,n43057 );
   not U29184 ( p2_u2843,n27738 );
   and U29185 ( n27740,n42794,n42795 );
   not U29186 ( p2_u2850,n27740 );
   and U29187 ( n27742,n43115,n43116 );
   not U29188 ( p2_u2841,n27742 );
   and U29189 ( n27744,n43087,n43088 );
   not U29190 ( p2_u2842,n27744 );
   and U29191 ( n27746,n43233,n43234 );
   not U29192 ( p2_u2837,n27746 );
   and U29193 ( n27748,n42999,n43000 );
   not U29194 ( p2_u2845,n27748 );
   and U29195 ( n27750,n42882,n42883 );
   not U29196 ( p2_u2849,n27750 );
   and U29197 ( n27752,n35796,n35797 );
   not U29198 ( p3_u2654,n27752 );
   and U29199 ( n27754,n38760,n38761 );
   not U29200 ( p2_u3044,n27754 );
   and U29201 ( n27756,n43147,n43148 );
   not U29202 ( p2_u2840,n27756 );
   and U29203 ( n27758,n43173,n43174 );
   not U29204 ( p2_u2839,n27758 );
   and U29205 ( n27760,n32560,n32561 );
   not U29206 ( p3_u2809,n27760 );
   and U29207 ( n27762,n42685,n42686 );
   not U29208 ( p2_u2853,n27762 );
   and U29209 ( n27764,n49911,n49912 );
   not U29210 ( p1_u2837,n27764 );
   and U29211 ( n27766,n35318,n35319 );
   not U29212 ( p3_u2672,n27766 );
   and U29213 ( n27768,n42971,n42972 );
   not U29214 ( p2_u2846,n27768 );
   and U29215 ( n27770,n42723,n42724 );
   not U29216 ( p2_u2852,n27770 );
   and U29217 ( n27772,n32286,n32287 );
   not U29218 ( p3_u2817,n27772 );
   and U29219 ( n27774,n33089,n36286 );
   not U29220 ( p3_u2637,n27774 );
   and U29221 ( n27776,n28811,n28812 );
   not U29222 ( p3_u3295,n27776 );
   and U29223 ( n27778,n42658,n42659 );
   not U29224 ( p2_u2854,n27778 );
   and U29225 ( n27780,n32420,n32421 );
   not U29226 ( p3_u2813,n27780 );
   and U29227 ( n27782,n32628,n32629 );
   not U29228 ( p3_u2807,n27782 );
   and U29229 ( n27784,n43491,n43492 );
   not U29230 ( p2_u2828,n27784 );
   and U29231 ( n27786,n43265,n43266 );
   not U29232 ( p2_u2836,n27786 );
   and U29233 ( n27788,n43574,n43575 );
   not U29234 ( p2_u2825,n27788 );
   and U29235 ( n27790,n42941,n42942 );
   not U29236 ( p2_u2847,n27790 );
   and U29237 ( n27792,n32839,n32840 );
   not U29238 ( p3_u2801,n27792 );
   and U29239 ( n27794,n32726,n32727 );
   not U29240 ( p3_u2804,n27794 );
   and U29241 ( n27796,n43517,n43518 );
   not U29242 ( p2_u2827,n27796 );
   and U29243 ( n27798,n43347,n43348 );
   not U29244 ( p2_u2833,n27798 );
   and U29245 ( n27800,n43403,n43404 );
   not U29246 ( p2_u2831,n27800 );
   and U29247 ( n27802,n43547,n43548 );
   not U29248 ( p2_u2826,n27802 );
   and U29249 ( n27804,n28741,n28742 );
   not U29250 ( u213,n27804 );
   and U29251 ( n27806,n42912,n42913 );
   not U29252 ( p2_u2848,n27806 );
   and U29253 ( n27808,n43378,n43379 );
   not U29254 ( p2_u2832,n27808 );
   and U29255 ( n27810,n43322,n43323 );
   not U29256 ( p2_u2834,n27810 );
   and U29257 ( n27812,n49884,n49885 );
   not U29258 ( p1_u2838,n27812 );
   and U29259 ( n27814,n42757,n42758 );
   not U29260 ( p2_u2851,n27814 );
   and U29261 ( n27816,n43291,n43292 );
   not U29262 ( p2_u2835,n27816 );
   and U29263 ( n27818,n43460,n43461 );
   not U29264 ( p2_u2829,n27818 );
   and U29265 ( n27820,n30901,n30902 );
   not U29266 ( p3_u2858,n27820 );
   and U29267 ( n27822,n44728,n44729 );
   not U29268 ( p2_u2816,n27822 );
   and U29269 ( n27824,n42623,n42624 );
   not U29270 ( p2_u2855,n27824 );
   and U29271 ( n27826,n43435,n43436 );
   not U29272 ( p2_u2830,n27826 );
   and U29273 ( n27828,n35399,n35400 );
   not U29274 ( p3_u2669,n27828 );
   and U29275 ( n27830,n43610,n43611 );
   not U29276 ( p2_u2824,n27830 );
   and U29277 ( n27832,n48392,n48393 );
   not U29278 ( p1_u2992,n27832 );
   and U29279 ( n27834,n48336,n48337 );
   not U29280 ( p1_u2996,n27834 );
   and U29281 ( n27836,n48461,n48462 );
   not U29282 ( p1_u2988,n27836 );
   and U29283 ( n27838,n31452,n31453 );
   not U29284 ( p3_u2839,n27838 );
   and U29285 ( n27840,n31381,n31382 );
   not U29286 ( p3_u2841,n27840 );
   and U29287 ( n27842,n28889,n28890 );
   not U29288 ( p3_u3282,n27842 );
   and U29289 ( n27844,n37030,n37031 );
   not U29290 ( p2_u3178,n27844 );
   and U29291 ( n27846,n37036,n37037 );
   not U29292 ( p2_u3177,n27846 );
   and U29293 ( n27848,n45438,n45439 );
   not U29294 ( p1_u3474,n27848 );
   and U29295 ( n27850,n36719,n36720 );
   not U29296 ( p2_u3601,n27850 );
   and U29297 ( n27852,n52747,n52748 );
   not U29298 ( p1_u2803,n27852 );
   and U29299 ( n27854,n48364,n48365 );
   not U29300 ( p1_u2994,n27854 );
   and U29301 ( n27856,n36320,n36321 );
   not U29302 ( p3_u2634,n27856 );
   and U29303 ( n27858,n36788,n36789 );
   not U29304 ( p2_u3593,n27858 );
   and U29305 ( n27860,n45762,n45763 );
   not U29306 ( p1_u3162,n27860 );
   and U29307 ( n27862,n30745,n30746 );
   not U29308 ( p3_u2866,n27862 );
   and U29309 ( n27864,n30765,n30766 );
   not U29310 ( p3_u2865,n27864 );
   and U29311 ( n27866,n29143,n29144 );
   not U29312 ( p3_u2998,n27866 );
   and U29313 ( n27868,n28895,n36607 );
   not U29314 ( p3_u2633,n27868 );
   and U29315 ( n27870,n45506,n52755 );
   not U29316 ( p1_u2802,n27870 );
   and U29317 ( n27872,n28163,n44735 );
   not U29318 ( p2_u2815,n27872 );
   and U29319 ( n27874,n36621,n36622 );
   not U29320 ( p2_u3610,n27874 );
   and U29321 ( n27876,n52758,n52759 );
   not U29322 ( p1_u2801,n27876 );
   and U29323 ( n27878,n44738,n44739 );
   not U29324 ( p2_u2814,n27878 );
   buf U29325 ( n27880,n41126 );
   buf U29326 ( n27881,n49257 );
   not U29327 ( n27882,n30338 );
   not U29328 ( n27883,n30348 );
   not U29329 ( n27884,n30328 );
   not U29330 ( n27885,n30358 );
   not U29331 ( n27886,n30318 );
   not U29332 ( n27887,n30368 );
   not U29333 ( n27888,n30305 );
   not U29334 ( n27889,n30387 );
   not U29335 ( n27890,n28268 );
   not U29336 ( n27891,n28188 );
   not U29337 ( n27892,n45876 );
   buf U29338 ( n27893,n33414 );
   not U29339 ( n27894,n28329 );
   not U29340 ( n27895,p2_state2_reg_0_ );
   not U29341 ( n27896,n28280 );
   buf U29342 ( n27897,n42772 );
   not U29343 ( n27898,n42655 );
   or U29344 ( n27899,n28165,n37029 );
   not U29345 ( p2_u3179,n27899 );
   or U29346 ( n27901,n28164,n37028 );
   not U29347 ( p2_u3180,n27901 );
   or U29348 ( n27903,n28165,n37027 );
   not U29349 ( p2_u3181,n27903 );
   or U29350 ( n27905,n28166,n37026 );
   not U29351 ( p2_u3182,n27905 );
   or U29352 ( n27907,n28167,n37025 );
   not U29353 ( p2_u3183,n27907 );
   or U29354 ( n27909,n28165,n37024 );
   not U29355 ( p2_u3184,n27909 );
   or U29356 ( n27911,n28164,n37023 );
   not U29357 ( p2_u3185,n27911 );
   or U29358 ( n27913,n28167,n37022 );
   not U29359 ( p2_u3186,n27913 );
   or U29360 ( n27915,n28166,n37021 );
   not U29361 ( p2_u3187,n27915 );
   or U29362 ( n27917,n28166,n37020 );
   not U29363 ( p2_u3188,n27917 );
   or U29364 ( n27919,n28164,n37019 );
   not U29365 ( p2_u3189,n27919 );
   or U29366 ( n27921,n28164,n37018 );
   not U29367 ( p2_u3190,n27921 );
   or U29368 ( n27923,n28166,n37017 );
   not U29369 ( p2_u3191,n27923 );
   or U29370 ( n27925,n28167,n37016 );
   not U29371 ( p2_u3192,n27925 );
   or U29372 ( n27927,n28164,n37015 );
   not U29373 ( p2_u3193,n27927 );
   or U29374 ( n27929,n28166,n37014 );
   not U29375 ( p2_u3194,n27929 );
   or U29376 ( n27931,n28167,n37013 );
   not U29377 ( p2_u3195,n27931 );
   or U29378 ( n27933,n28166,n37012 );
   not U29379 ( p2_u3196,n27933 );
   or U29380 ( n27935,n28165,n37011 );
   not U29381 ( p2_u3197,n27935 );
   or U29382 ( n27937,n28165,n37010 );
   not U29383 ( p2_u3198,n27937 );
   or U29384 ( n27939,n28164,n37009 );
   not U29385 ( p2_u3199,n27939 );
   or U29386 ( n27941,n28166,n37008 );
   not U29387 ( p2_u3200,n27941 );
   or U29388 ( n27943,n28167,n37007 );
   not U29389 ( p2_u3201,n27943 );
   or U29390 ( n27945,n28164,n37006 );
   not U29391 ( p2_u3202,n27945 );
   or U29392 ( n27947,n28167,n37005 );
   not U29393 ( p2_u3203,n27947 );
   or U29394 ( n27949,n28165,n37004 );
   not U29395 ( p2_u3204,n27949 );
   or U29396 ( n27951,n28167,n37003 );
   not U29397 ( p2_u3205,n27951 );
   or U29398 ( n27953,n28166,n37002 );
   not U29399 ( p2_u3206,n27953 );
   or U29400 ( n27955,n28165,n37001 );
   not U29401 ( p2_u3207,n27955 );
   or U29402 ( n27957,n28165,n37000 );
   not U29403 ( p2_u3208,n27957 );
   or U29404 ( n27959,n28737,n41121 );
   not U29405 ( p2_u2920,n27959 );
   or U29406 ( n27961,n33401,n28475 );
   not U29407 ( p3_u2736,n27961 );
   not U29408 ( n27963,n53143 );
   not U29409 ( p1_u3193,n27963 );
   not U29410 ( n27965,n53144 );
   not U29411 ( p1_u3192,n27965 );
   not U29412 ( n27967,n53145 );
   not U29413 ( p1_u3191,n27967 );
   not U29414 ( n27969,n53146 );
   not U29415 ( p1_u3190,n27969 );
   not U29416 ( n27971,n53147 );
   not U29417 ( p1_u3189,n27971 );
   not U29418 ( n27973,n53148 );
   not U29419 ( p1_u3188,n27973 );
   not U29420 ( n27975,n53149 );
   not U29421 ( p1_u3187,n27975 );
   not U29422 ( n27977,n53150 );
   not U29423 ( p1_u3186,n27977 );
   not U29424 ( n27979,n53151 );
   not U29425 ( p1_u3185,n27979 );
   not U29426 ( n27981,n53152 );
   not U29427 ( p1_u3184,n27981 );
   not U29428 ( n27983,n53153 );
   not U29429 ( p1_u3183,n27983 );
   not U29430 ( n27985,n53154 );
   not U29431 ( p1_u3182,n27985 );
   not U29432 ( n27987,n53155 );
   not U29433 ( p1_u3181,n27987 );
   not U29434 ( n27989,n53156 );
   not U29435 ( p1_u3180,n27989 );
   not U29436 ( n27991,n53157 );
   not U29437 ( p1_u3179,n27991 );
   not U29438 ( n27993,n53158 );
   not U29439 ( p1_u3178,n27993 );
   not U29440 ( n27995,n53159 );
   not U29441 ( p1_u3177,n27995 );
   not U29442 ( n27997,n53160 );
   not U29443 ( p1_u3176,n27997 );
   not U29444 ( n27999,n53161 );
   not U29445 ( p1_u3175,n27999 );
   not U29446 ( n28001,n53162 );
   not U29447 ( p1_u3174,n28001 );
   not U29448 ( n28003,n53163 );
   not U29449 ( p1_u3173,n28003 );
   not U29450 ( n28005,n53164 );
   not U29451 ( p1_u3172,n28005 );
   not U29452 ( n28007,n53165 );
   not U29453 ( p1_u3171,n28007 );
   not U29454 ( n28009,n53166 );
   not U29455 ( p1_u3170,n28009 );
   not U29456 ( n28011,n53167 );
   not U29457 ( p1_u3169,n28011 );
   not U29458 ( n28013,n53168 );
   not U29459 ( p1_u3168,n28013 );
   not U29460 ( n28015,n53169 );
   not U29461 ( p1_u3167,n28015 );
   or U29462 ( n28017,n45508,n45749 );
   not U29463 ( p1_u3166,n28017 );
   not U29464 ( n28019,n53170 );
   not U29465 ( p1_u3165,n28019 );
   or U29466 ( n28021,n28156,n45751 );
   not U29467 ( p1_u3164,n28021 );
   or U29468 ( n28023,n31736,n31737 );
   not U29469 ( p3_u2831,n28023 );
   or U29470 ( n28025,n29232,n30744 );
   not U29471 ( p3_u2867,n28025 );
   not U29472 ( n28027,n53142 );
   not U29473 ( p3_u2999,n28027 );
   not U29474 ( n28029,n53141 );
   not U29475 ( p3_u3000,n28029 );
   not U29476 ( n28031,n53140 );
   not U29477 ( p3_u3001,n28031 );
   not U29478 ( n28033,n53139 );
   not U29479 ( p3_u3002,n28033 );
   not U29480 ( n28035,n53138 );
   not U29481 ( p3_u3003,n28035 );
   not U29482 ( n28037,n53137 );
   not U29483 ( p3_u3004,n28037 );
   not U29484 ( n28039,n53136 );
   not U29485 ( p3_u3005,n28039 );
   not U29486 ( n28041,n53135 );
   not U29487 ( p3_u3006,n28041 );
   not U29488 ( n28043,n53134 );
   not U29489 ( p3_u3007,n28043 );
   not U29490 ( n28045,n53133 );
   not U29491 ( p3_u3008,n28045 );
   not U29492 ( n28047,n53132 );
   not U29493 ( p3_u3009,n28047 );
   not U29494 ( n28049,n53131 );
   not U29495 ( p3_u3010,n28049 );
   not U29496 ( n28051,n53130 );
   not U29497 ( p3_u3011,n28051 );
   not U29498 ( n28053,n53129 );
   not U29499 ( p3_u3012,n28053 );
   not U29500 ( n28055,n53128 );
   not U29501 ( p3_u3013,n28055 );
   not U29502 ( n28057,n53127 );
   not U29503 ( p3_u3014,n28057 );
   not U29504 ( n28059,n53126 );
   not U29505 ( p3_u3015,n28059 );
   not U29506 ( n28061,n53125 );
   not U29507 ( p3_u3016,n28061 );
   not U29508 ( n28063,n53124 );
   not U29509 ( p3_u3017,n28063 );
   not U29510 ( n28065,n53123 );
   not U29511 ( p3_u3018,n28065 );
   not U29512 ( n28067,n53122 );
   not U29513 ( p3_u3019,n28067 );
   not U29514 ( n28069,n53121 );
   not U29515 ( p3_u3020,n28069 );
   not U29516 ( n28071,n53120 );
   not U29517 ( p3_u3021,n28071 );
   not U29518 ( n28073,n53119 );
   not U29519 ( p3_u3022,n28073 );
   not U29520 ( n28075,n53118 );
   not U29521 ( p3_u3023,n28075 );
   not U29522 ( n28077,n53117 );
   not U29523 ( p3_u3024,n28077 );
   not U29524 ( n28079,n53116 );
   not U29525 ( p3_u3025,n28079 );
   or U29526 ( n28081,n28158,n29115 );
   not U29527 ( p3_u3026,n28081 );
   or U29528 ( n28083,n28897,n29114 );
   not U29529 ( p3_u3027,n28083 );
   not U29530 ( n28085,n53115 );
   not U29531 ( p3_u3028,n28085 );
   or U29532 ( n28087,n28479,n49328 );
   not U29533 ( p1_u2905,n28087 );
   not U29534 ( n28089,n53114 );
   not U29535 ( n28090,n28260 );
   buf U29536 ( n28091,n41761 );
   not U29537 ( n28092,n42638 );
   buf U29538 ( n28093,n42634 );
   not U29539 ( n28095,p1_state2_reg_0_ );
   not U29540 ( n28094,p1_state2_reg_0_ );
   not U29541 ( n28096,n25182 );
   not U29542 ( n28098,n25182 );
   not U29543 ( n28097,n25182 );
   not U29544 ( n28099,n41044 );
   not U29545 ( n28101,n28099 );
   not U29546 ( n28100,n28099 );
   not U29547 ( n28103,n49818 );
   not U29548 ( n28102,n49818 );
   not U29549 ( n28104,n25183 );
   not U29550 ( n28106,n25183 );
   not U29551 ( n28105,n25183 );
   nor U29552 ( n28107,n49663,n47426 );
   not U29553 ( n28108,n28107 );
   not U29554 ( n28110,n28107 );
   not U29555 ( n28109,n28107 );
   nand U29556 ( n28112,n28790,n33401 );
   nand U29557 ( n28111,n28790,n33401 );
   nand U29558 ( n28114,n28374,n47473 );
   nand U29559 ( n28113,n28374,n47473 );
   nand U29560 ( n28116,n28132,n28160 );
   nand U29561 ( n28115,n28132,n28160 );
   and U29562 ( n28117,n45352,n28395 );
   not U29563 ( n28118,n28117 );
   not U29564 ( n28120,n28117 );
   not U29565 ( n28119,n28117 );
   not U29566 ( n28122,n44609 );
   not U29567 ( n28121,n44609 );
   nand U29568 ( n28124,n40865,p2_statebs16_reg );
   nand U29569 ( n28123,n40865,p2_statebs16_reg );
   nand U29570 ( n28126,n28808,n30836 );
   nand U29571 ( n28125,n28808,n30836 );
   not U29572 ( n28127,n33418 );
   not U29573 ( n28129,n28127 );
   not U29574 ( n28128,n28127 );
   and U29575 ( n28130,n28757,n28758 );
   not U29576 ( u214,n28130 );
   not U29577 ( n28132,n28130 );
   nand U29578 ( n28134,n33086,p3_statebs16_reg );
   nand U29579 ( n28133,n33086,p3_statebs16_reg );
   nand U29580 ( n28136,n28781,n29080 );
   nand U29581 ( n28135,n28781,n29080 );
   nand U29582 ( n28138,n45333,n45689 );
   nand U29583 ( n28137,n45333,n45689 );
   not U29584 ( n28139,n28250 );
   not U29585 ( n28141,n28250 );
   not U29586 ( n28140,n49841 );
   and U29587 ( n28142,n33241,n29304 );
   not U29588 ( n28143,n28142 );
   not U29589 ( n28146,n28142 );
   not U29590 ( n28144,n28142 );
   not U29591 ( n28145,n28142 );
   nand U29592 ( n28148,n37045,n42618 );
   nand U29593 ( n28147,n37045,n42618 );
   nand U29594 ( n28150,n44600,n44598 );
   nand U29595 ( n28149,n44600,n44598 );
   not U29596 ( n28151,n41765 );
   not U29597 ( n28152,n28151 );
   not U29598 ( n28153,n28151 );
   not U29599 ( n28154,n28151 );
   not U29600 ( n28156,n45506 );
   not U29601 ( n28155,n45506 );
   not U29602 ( n28158,n28895 );
   not U29603 ( n28157,n28895 );
   not U29604 ( n28159,n25181 );
   not U29605 ( n28162,n25181 );
   not U29606 ( n28160,n25181 );
   not U29607 ( n28161,n25181 );
   and U29608 ( n28163,n36987,n44736 );
   not U29609 ( n28164,n28163 );
   not U29610 ( n28167,n28163 );
   not U29611 ( n28165,n28163 );
   not U29612 ( n28166,n28163 );
   nand U29613 ( n28169,n32970,n32966 );
   nand U29614 ( n28168,n32970,n32966 );
   not U29615 ( n28170,n34238 );
   not U29616 ( n28171,n28170 );
   not U29617 ( n28173,n28170 );
   not U29618 ( n28172,n28170 );
   not U29619 ( n28174,n32131 );
   not U29620 ( n28175,n28174 );
   not U29621 ( n28176,n28174 );
   not U29622 ( n28177,n28174 );
   not U29623 ( n28178,p2_state2_reg_1_ );
   not U29624 ( n28181,p2_state2_reg_1_ );
   not U29625 ( n28179,p2_state2_reg_1_ );
   not U29626 ( n28180,p2_state2_reg_1_ );
   not U29627 ( n28182,n28407 );
   not U29628 ( n28185,n49843 );
   not U29629 ( n28183,n28408 );
   not U29630 ( n28184,n49843 );
   not U29631 ( n28186,n28089 );
   not U29632 ( u215,n28089 );
   buf U29633 ( n28188,n28739 );
   buf U29634 ( n28189,n45897 );
   buf U29635 ( n28190,n29388 );
   buf U29636 ( n28191,n29394 );
   buf U29637 ( n28192,n45890 );
   buf U29638 ( n28193,n37236 );
   buf U29639 ( n28194,n45909 );
   buf U29640 ( n28195,n29402 );
   buf U29641 ( n28196,n29406 );
   buf U29642 ( n28197,n37229 );
   buf U29643 ( n28198,n45905 );
   buf U29644 ( n28199,n37248 );
   buf U29645 ( n28200,n45921 );
   buf U29646 ( n28201,n29414 );
   buf U29647 ( n28202,n29418 );
   buf U29648 ( n28203,n37244 );
   buf U29649 ( n28204,n45917 );
   not U29650 ( n28205,n47512 );
   buf U29651 ( n28206,n37260 );
   buf U29652 ( n28207,n45933 );
   buf U29653 ( n28208,n29426 );
   buf U29654 ( n28209,n29430 );
   buf U29655 ( n28210,n37256 );
   buf U29656 ( n28211,n45929 );
   buf U29657 ( n28212,n49445 );
   not U29658 ( n28213,n47466 );
   buf U29659 ( n28214,n37272 );
   buf U29660 ( n28215,n45945 );
   buf U29661 ( n28216,n29438 );
   buf U29662 ( n28217,n29442 );
   buf U29663 ( n28218,n37268 );
   buf U29664 ( n28219,n45941 );
   not U29665 ( n28220,n50566 );
   not U29666 ( n28221,n30836 );
   not U29667 ( n28222,n31045 );
   buf U29668 ( n28223,n49448 );
   buf U29669 ( n28224,n49339 );
   buf U29670 ( n28225,n40889 );
   buf U29671 ( n28226,n37284 );
   buf U29672 ( n28227,n45957 );
   buf U29673 ( n28228,n29450 );
   buf U29674 ( n28229,n29454 );
   buf U29675 ( n28230,n37280 );
   buf U29676 ( n28231,n45953 );
   not U29677 ( n28232,n47473 );
   buf U29678 ( n28233,n33983 );
   not U29679 ( n28234,n39573 );
   buf U29680 ( n28235,n30811 );
   not U29681 ( n28236,n38769 );
   buf U29682 ( n28237,n41346 );
   not U29683 ( n28238,n47489 );
   buf U29684 ( n28239,n38601 );
   not U29685 ( n28240,n30851 );
   not U29686 ( n28241,n28262 );
   not U29687 ( n28242,n35376 );
   not U29688 ( n28243,n28261 );
   buf U29689 ( n28244,n37308 );
   buf U29690 ( n28245,n45969 );
   buf U29691 ( n28246,n29462 );
   buf U29692 ( n28247,n29466 );
   buf U29693 ( n28248,n37292 );
   buf U29694 ( n28249,n45965 );
   buf U29695 ( n28250,n49841 );
   not U29696 ( n28252,n49013 );
   not U29697 ( n28251,n49013 );
   nand U29698 ( n28253,n48159,n45444 );
   buf U29699 ( n28254,n33098 );
   buf U29700 ( n28255,n41045 );
   buf U29701 ( n28256,n41221 );
   buf U29702 ( n28257,n33251 );
   buf U29703 ( n28258,n49028 );
   not U29704 ( n28259,n41232 );
   buf U29705 ( n28260,n35448 );
   buf U29706 ( n28261,n49335 );
   buf U29707 ( n28262,n50737 );
   not U29708 ( n28263,n31956 );
   not U29709 ( n28264,n28379 );
   not U29710 ( n28265,n48647 );
   buf U29711 ( n28266,n30930 );
   buf U29712 ( n28267,n37296 );
   buf U29713 ( n28268,n48298 );
   not U29714 ( n28269,n38746 );
   buf U29715 ( n28270,n29488 );
   buf U29716 ( n28271,n29496 );
   buf U29717 ( n28272,n37304 );
   buf U29718 ( n28273,n45999 );
   buf U29719 ( n28274,n42987 );
   not U29720 ( n28275,n38744 );
   not U29721 ( n28276,n52625 );
   not U29722 ( n28277,n35379 );
   not U29723 ( n28278,n28352 );
   not U29724 ( n28279,n49882 );
   buf U29725 ( n28280,n36646 );
   not U29726 ( n28281,n45992 );
   not U29727 ( n28282,n40219 );
   buf U29728 ( n28283,n34233 );
   buf U29729 ( n28284,n49023 );
   not U29730 ( n28285,n40196 );
   buf U29731 ( n28286,n49851 );
   not U29732 ( n28288,n50593 );
   not U29733 ( n28287,n50593 );
   nand U29734 ( n28290,n49011,n49012 );
   nand U29735 ( n28289,n49011,n49012 );
   not U29736 ( n28291,n33413 );
   nand U29737 ( n28292,n48245,n48246 );
   not U29738 ( n28293,n28292 );
   not U29739 ( n28296,n28292 );
   not U29740 ( n28294,n28292 );
   not U29741 ( n28295,n28292 );
   nor U29742 ( n28297,n33251,n28771 );
   not U29743 ( n28298,n28297 );
   not U29744 ( n28299,n28297 );
   not U29745 ( n28300,n47613 );
   buf U29746 ( n28301,n38758 );
   buf U29747 ( n28302,n33417 );
   buf U29748 ( n28303,n37326 );
   not U29749 ( n28304,n38757 );
   buf U29750 ( n28305,n47466 );
   not U29751 ( n28306,n41862 );
   not U29752 ( n28307,n49443 );
   not U29753 ( n28308,n38472 );
   not U29754 ( n28309,n38482 );
   not U29755 ( n28310,n38491 );
   not U29756 ( n28311,n38500 );
   not U29757 ( n28312,n38509 );
   not U29758 ( n28313,n38518 );
   not U29759 ( n28314,n38527 );
   not U29760 ( n28315,n38551 );
   not U29761 ( n28316,n47143 );
   not U29762 ( n28317,n47153 );
   not U29763 ( n28318,n47162 );
   not U29764 ( n28319,n47171 );
   not U29765 ( n28320,n47180 );
   not U29766 ( n28321,n47189 );
   not U29767 ( n28322,n47198 );
   not U29768 ( n28323,n47222 );
   buf U29769 ( n28324,n37344 );
   buf U29770 ( n28325,n46006 );
   not U29771 ( n28326,n38937 );
   not U29772 ( n28327,n48996 );
   buf U29773 ( n28328,n37337 );
   buf U29774 ( n28329,n28765 );
   not U29775 ( n28330,n44156 );
   not U29776 ( n28331,n42664 );
   not U29777 ( n28332,n33401 );
   not U29778 ( n28333,n35378 );
   not U29779 ( n28334,n49979 );
   not U29780 ( n28335,n33241 );
   not U29781 ( n28336,n41032 );
   buf U29782 ( n28337,n30830 );
   buf U29783 ( n28338,n47519 );
   not U29784 ( n28339,n35386 );
   not U29785 ( n28340,n42639 );
   buf U29786 ( n28341,n48647 );
   not U29787 ( n28342,n52632 );
   not U29788 ( n28343,n38733 );
   not U29789 ( n28344,n48305 );
   not U29790 ( n28345,n39595 );
   not U29791 ( n28346,n39427 );
   not U29792 ( n28347,n39603 );
   buf U29793 ( n28348,n49663 );
   not U29794 ( n28349,n31929 );
   not U29795 ( n28350,n29487 );
   buf U29796 ( n28351,n30841 );
   buf U29797 ( n28352,n28414 );
   not U29798 ( n28353,n39596 );
   not U29799 ( n28354,n49856 );
   not U29800 ( n28355,n42744 );
   not U29801 ( n28356,n31923 );
   not U29802 ( n28357,n41121 );
   not U29803 ( n28358,n49837 );
   not U29804 ( n28359,n32178 );
   buf U29805 ( n28360,n42657 );
   not U29806 ( n28361,n42988 );
   not U29807 ( n28362,n28361 );
   not U29808 ( n28363,n28361 );
   not U29809 ( n28364,n49328 );
   not U29810 ( n28365,n33413 );
   not U29811 ( n28366,n28365 );
   not U29812 ( n28367,n28365 );
   not U29813 ( n28369,n44130 );
   not U29814 ( n28368,n44130 );
   not U29815 ( n28370,n28282 );
   not U29816 ( n28371,n28282 );
   not U29817 ( n28373,n41295 );
   not U29818 ( n28372,n41295 );
   not U29819 ( n28375,p1_state2_reg_2_ );
   not U29820 ( n28374,p1_state2_reg_2_ );
   not U29821 ( n28376,n28781 );
   not U29822 ( n28377,n36620 );
   not U29823 ( n28378,n45333 );
   nand U29824 ( n28380,n36215,n36216 );
   nand U29825 ( n28379,n36215,n36216 );
   nand U29826 ( n28382,n40878,n40879 );
   nand U29827 ( n28381,n40878,n40879 );
   not U29828 ( n28384,n43676 );
   not U29829 ( n28383,n43676 );
   not U29830 ( n28386,n36962 );
   not U29831 ( n28385,n36962 );
   not U29832 ( n28388,n36960 );
   not U29833 ( n28387,n36960 );
   not U29834 ( n28390,n43677 );
   not U29835 ( n28389,n43677 );
   not U29836 ( n28392,n29065 );
   not U29837 ( n28391,n29065 );
   not U29838 ( n28394,n45675 );
   not U29839 ( n28393,n45675 );
   nand U29840 ( n28396,n49017,n49018 );
   nand U29841 ( n28395,n49017,n49018 );
   nand U29842 ( n28397,n49171,n49172 );
   not U29843 ( n28398,n28397 );
   not U29844 ( n28401,n28397 );
   not U29845 ( n28399,n28397 );
   not U29846 ( n28400,n28397 );
   buf U29847 ( n28402,n45329 );
   not U29848 ( n28403,n28402 );
   not U29849 ( n28406,n28402 );
   not U29850 ( n28404,n28402 );
   not U29851 ( n28405,n28402 );
   nor U29852 ( n28408,p1_state2_reg_2_,p1_statebs16_reg );
   nor U29853 ( n28407,p1_state2_reg_2_,p1_statebs16_reg );
   nor U29854 ( n28410,n43894,n43658 );
   nor U29855 ( n28409,n43894,n43658 );
   nand U29856 ( n28412,p2_address_reg_0_,n28278 );
   nand U29857 ( n28411,n28414,p3_address_reg_0_ );
   nand U29858 ( n28416,p2_address_reg_10_,n28278 );
   nand U29859 ( n28415,n28352,p3_address_reg_10_ );
   nand U29860 ( n28418,p2_address_reg_11_,n28413 );
   nand U29861 ( n28417,n28352,p3_address_reg_11_ );
   nand U29862 ( n28420,p2_address_reg_12_,n28413 );
   nand U29863 ( n28419,n28414,p3_address_reg_12_ );
   nand U29864 ( n28422,p2_address_reg_13_,n28413 );
   nand U29865 ( n28421,n28414,p3_address_reg_13_ );
   nand U29866 ( n28424,p2_address_reg_14_,n28413 );
   nand U29867 ( n28423,n28414,p3_address_reg_14_ );
   nand U29868 ( n28426,p2_address_reg_15_,n28413 );
   nand U29869 ( n28425,n28414,p3_address_reg_15_ );
   nand U29870 ( n28428,p2_address_reg_16_,n28413 );
   nand U29871 ( n28427,n28414,p3_address_reg_16_ );
   nand U29872 ( n28430,p2_address_reg_17_,n28413 );
   nand U29873 ( n28429,n28414,p3_address_reg_17_ );
   nand U29874 ( n28432,p2_address_reg_18_,n28413 );
   nand U29875 ( n28431,n28414,p3_address_reg_18_ );
   nand U29876 ( n28434,p2_address_reg_19_,n28413 );
   nand U29877 ( n28433,n28414,p3_address_reg_19_ );
   nand U29878 ( n28436,p2_address_reg_1_,n28413 );
   nand U29879 ( n28435,n28414,p3_address_reg_1_ );
   nand U29880 ( n28438,p2_address_reg_20_,n28413 );
   nand U29881 ( n28437,n28414,p3_address_reg_20_ );
   nand U29882 ( n28440,p2_address_reg_21_,n28413 );
   nand U29883 ( n28439,n28414,p3_address_reg_21_ );
   nand U29884 ( n28442,p2_address_reg_22_,n28413 );
   nand U29885 ( n28441,n28414,p3_address_reg_22_ );
   nand U29886 ( n28444,p2_address_reg_23_,n28413 );
   nand U29887 ( n28443,n28414,p3_address_reg_23_ );
   nand U29888 ( n28446,p2_address_reg_24_,n28413 );
   nand U29889 ( n28445,n28352,p3_address_reg_24_ );
   nand U29890 ( n28448,p2_address_reg_25_,n28413 );
   nand U29891 ( n28447,n28352,p3_address_reg_25_ );
   nand U29892 ( n28450,p2_address_reg_26_,n28413 );
   nand U29893 ( n28449,n28352,p3_address_reg_26_ );
   nand U29894 ( n28452,p2_address_reg_27_,n28413 );
   nand U29895 ( n28451,n28352,p3_address_reg_27_ );
   nand U29896 ( n28454,p2_address_reg_28_,n28413 );
   nand U29897 ( n28453,n28352,p3_address_reg_28_ );
   nand U29898 ( n28456,p2_address_reg_29_,n28413 );
   nand U29899 ( n28455,n28352,p3_address_reg_29_ );
   nand U29900 ( n28458,p2_address_reg_2_,n28413 );
   nand U29901 ( n28457,n28352,p3_address_reg_2_ );
   nand U29902 ( n28460,p2_address_reg_3_,n28278 );
   nand U29903 ( n28459,n28352,p3_address_reg_3_ );
   nand U29904 ( n28462,p2_address_reg_4_,n28278 );
   nand U29905 ( n28461,n28352,p3_address_reg_4_ );
   nand U29906 ( n28464,p2_address_reg_5_,n28278 );
   nand U29907 ( n28463,n28352,p3_address_reg_5_ );
   nand U29908 ( n28466,p2_address_reg_6_,n28278 );
   nand U29909 ( n28465,n28352,p3_address_reg_6_ );
   nand U29910 ( n28468,p2_address_reg_7_,n28278 );
   nand U29911 ( n28467,n28352,p3_address_reg_7_ );
   nand U29912 ( n28470,p2_address_reg_8_,n28278 );
   nand U29913 ( n28469,n28352,p3_address_reg_8_ );
   nand U29914 ( n28472,p2_address_reg_9_,n28278 );
   nand U29915 ( n28471,n28414,p3_address_reg_9_ );
   not U29916 ( n28414,n28413 );
   nand U29917 ( n28413,n28473,n28474 );
   nand U29918 ( n28474,p3_datao_reg_30_,n28475 );
   nor U29919 ( n28473,n28476,n28477 );
   nor U29920 ( n28477,p2_datao_reg_31_,n28478 );
   and U29921 ( n28476,n28479,p1_datao_reg_30_ );
   nand U29922 ( n28481,buf2_reg_31_,n53114 );
   nand U29923 ( n28480,p2_datao_reg_31_,n28089 );
   nand U29924 ( n28484,buf2_reg_30_,n53114 );
   nand U29925 ( n28483,p2_datao_reg_30_,n28482 );
   nand U29926 ( n28486,buf2_reg_29_,n28186 );
   nand U29927 ( n28485,p2_datao_reg_29_,n28089 );
   nand U29928 ( n28488,buf2_reg_28_,n53114 );
   nand U29929 ( n28487,p2_datao_reg_28_,n28089 );
   nand U29930 ( n28490,buf2_reg_27_,n28186 );
   nand U29931 ( n28489,p2_datao_reg_27_,n28089 );
   nand U29932 ( n28492,buf2_reg_26_,n53114 );
   nand U29933 ( n28491,p2_datao_reg_26_,n28089 );
   nand U29934 ( n28494,buf2_reg_25_,n28186 );
   nand U29935 ( n28493,p2_datao_reg_25_,n28089 );
   nand U29936 ( n28496,buf2_reg_24_,n28186 );
   nand U29937 ( n28495,p2_datao_reg_24_,n28089 );
   nand U29938 ( n28498,buf2_reg_23_,n53114 );
   nand U29939 ( n28497,p2_datao_reg_23_,n28089 );
   nand U29940 ( n28500,buf2_reg_22_,n53114 );
   nand U29941 ( n28499,p2_datao_reg_22_,n28089 );
   nand U29942 ( n28502,buf2_reg_21_,n28186 );
   nand U29943 ( n28501,p2_datao_reg_21_,n28089 );
   nand U29944 ( n28504,buf2_reg_20_,n53114 );
   nand U29945 ( n28503,p2_datao_reg_20_,n28089 );
   nand U29946 ( n28506,buf2_reg_19_,n28186 );
   nand U29947 ( n28505,p2_datao_reg_19_,n28482 );
   nand U29948 ( n28508,buf2_reg_18_,n28186 );
   nand U29949 ( n28507,p2_datao_reg_18_,n28482 );
   nand U29950 ( n28510,buf2_reg_17_,n53114 );
   nand U29951 ( n28509,p2_datao_reg_17_,n28482 );
   nand U29952 ( n28512,buf2_reg_16_,n53114 );
   nand U29953 ( n28511,p2_datao_reg_16_,n28482 );
   nand U29954 ( n28514,buf2_reg_15_,n28186 );
   nand U29955 ( n28513,p2_datao_reg_15_,n28482 );
   nand U29956 ( n28516,buf2_reg_14_,n28186 );
   nand U29957 ( n28515,p2_datao_reg_14_,n28482 );
   nand U29958 ( n28518,buf2_reg_13_,n53114 );
   nand U29959 ( n28517,p2_datao_reg_13_,n28482 );
   nand U29960 ( n28520,buf2_reg_12_,n28186 );
   nand U29961 ( n28519,p2_datao_reg_12_,n28482 );
   nand U29962 ( n28522,buf2_reg_11_,n53114 );
   nand U29963 ( n28521,p2_datao_reg_11_,n28482 );
   nand U29964 ( n28524,buf2_reg_10_,n53114 );
   nand U29965 ( n28523,p2_datao_reg_10_,n28482 );
   nand U29966 ( n28526,buf2_reg_9_,n28186 );
   nand U29967 ( n28525,p2_datao_reg_9_,n28482 );
   nand U29968 ( n28528,buf2_reg_8_,n53114 );
   nand U29969 ( n28527,p2_datao_reg_8_,n28482 );
   nand U29970 ( n28530,buf2_reg_7_,n28186 );
   nand U29971 ( n28529,p2_datao_reg_7_,n28482 );
   nand U29972 ( n28532,buf2_reg_6_,n53114 );
   nand U29973 ( n28531,p2_datao_reg_6_,n28482 );
   nand U29974 ( n28534,buf2_reg_5_,n28186 );
   nand U29975 ( n28533,p2_datao_reg_5_,n28482 );
   nand U29976 ( n28536,buf2_reg_4_,n53114 );
   nand U29977 ( n28535,p2_datao_reg_4_,n28482 );
   nand U29978 ( n28538,buf2_reg_3_,n28186 );
   nand U29979 ( n28537,p2_datao_reg_3_,n28482 );
   nand U29980 ( n28540,buf2_reg_2_,n28186 );
   nand U29981 ( n28539,p2_datao_reg_2_,n28089 );
   nand U29982 ( n28542,buf2_reg_1_,n53114 );
   nand U29983 ( n28541,p2_datao_reg_1_,n28482 );
   nand U29984 ( n28544,buf2_reg_0_,n28186 );
   nand U29985 ( n28543,p2_datao_reg_0_,n28089 );
   nand U29986 ( n28546,p1_datao_reg_0_,n28130 );
   nor U29987 ( n28545,n28548,n28549 );
   nor U29988 ( n28549,n28162,n28550 );
   nor U29989 ( n28548,n28551,n28552 );
   not U29990 ( n28551,p2_datao_reg_0_ );
   nand U29991 ( n28554,p1_datao_reg_1_,n28130 );
   nor U29992 ( n28553,n28555,n28556 );
   nor U29993 ( n28556,n28159,n28557 );
   nor U29994 ( n28555,n28558,n28552 );
   not U29995 ( n28558,p2_datao_reg_1_ );
   nand U29996 ( n28560,p1_datao_reg_2_,n28547 );
   nor U29997 ( n28559,n28561,n28562 );
   nor U29998 ( n28562,n28161,n28563 );
   nor U29999 ( n28561,n28564,n28115 );
   not U30000 ( n28564,p2_datao_reg_2_ );
   nand U30001 ( n28566,p1_datao_reg_3_,n28130 );
   nor U30002 ( n28565,n28567,n28568 );
   nor U30003 ( n28568,n28160,n28569 );
   nor U30004 ( n28567,n28570,n28116 );
   not U30005 ( n28570,p2_datao_reg_3_ );
   nand U30006 ( n28572,p1_datao_reg_4_,n28547 );
   nor U30007 ( n28571,n28573,n28574 );
   nor U30008 ( n28574,n28162,n28575 );
   nor U30009 ( n28573,n28576,n28552 );
   not U30010 ( n28576,p2_datao_reg_4_ );
   nand U30011 ( n28578,p1_datao_reg_5_,n28547 );
   nor U30012 ( n28577,n28579,n28580 );
   nor U30013 ( n28580,n28159,n28581 );
   nor U30014 ( n28579,n28582,n28115 );
   not U30015 ( n28582,p2_datao_reg_5_ );
   nand U30016 ( n28584,p1_datao_reg_6_,n28547 );
   nor U30017 ( n28583,n28585,n28586 );
   nor U30018 ( n28586,n28161,n28587 );
   nor U30019 ( n28585,n28588,n28116 );
   not U30020 ( n28588,p2_datao_reg_6_ );
   nand U30021 ( n28590,p1_datao_reg_7_,n28547 );
   nor U30022 ( n28589,n28591,n28592 );
   nor U30023 ( n28592,n28160,n28593 );
   nor U30024 ( n28591,n28594,n28552 );
   not U30025 ( n28594,p2_datao_reg_7_ );
   nand U30026 ( n28596,p1_datao_reg_8_,n28547 );
   nor U30027 ( n28595,n28597,n28598 );
   nor U30028 ( n28598,n28162,n28599 );
   nor U30029 ( n28597,n28600,n28115 );
   not U30030 ( n28600,p2_datao_reg_8_ );
   nand U30031 ( n28602,p1_datao_reg_9_,n28547 );
   nor U30032 ( n28601,n28603,n28604 );
   nor U30033 ( n28604,n28159,n28605 );
   nor U30034 ( n28603,n28606,n28116 );
   not U30035 ( n28606,p2_datao_reg_9_ );
   nand U30036 ( n28608,p1_datao_reg_10_,n28547 );
   nor U30037 ( n28607,n28609,n28610 );
   nor U30038 ( n28610,n28161,n28611 );
   nor U30039 ( n28609,n28612,n28552 );
   not U30040 ( n28612,p2_datao_reg_10_ );
   nand U30041 ( n28614,p1_datao_reg_11_,n28547 );
   nor U30042 ( n28613,n28615,n28616 );
   nor U30043 ( n28616,n28160,n28617 );
   nor U30044 ( n28615,n28618,n28115 );
   not U30045 ( n28618,p2_datao_reg_11_ );
   nand U30046 ( n28620,p1_datao_reg_12_,n28547 );
   nor U30047 ( n28619,n28621,n28622 );
   nor U30048 ( n28622,n28162,n28623 );
   nor U30049 ( n28621,n28624,n28116 );
   not U30050 ( n28624,p2_datao_reg_12_ );
   nand U30051 ( n28626,p1_datao_reg_13_,n28547 );
   nor U30052 ( n28625,n28627,n28628 );
   nor U30053 ( n28628,n28159,n28629 );
   nor U30054 ( n28627,n28630,n28115 );
   not U30055 ( n28630,p2_datao_reg_13_ );
   nand U30056 ( n28632,p1_datao_reg_14_,n28547 );
   nor U30057 ( n28631,n28633,n28634 );
   nor U30058 ( n28634,n28161,n28635 );
   nor U30059 ( n28633,n28636,n28552 );
   not U30060 ( n28636,p2_datao_reg_14_ );
   nand U30061 ( n28638,p1_datao_reg_15_,n28547 );
   nor U30062 ( n28637,n28639,n28640 );
   nor U30063 ( n28640,n28160,n28641 );
   not U30064 ( n28641,buf1_reg_15_ );
   nor U30065 ( n28639,n28642,n28116 );
   not U30066 ( n28642,p2_datao_reg_15_ );
   nand U30067 ( n28644,p1_datao_reg_16_,n28547 );
   nor U30068 ( n28643,n28645,n28646 );
   nor U30069 ( n28646,n28162,n28647 );
   nor U30070 ( n28645,n28648,n28115 );
   not U30071 ( n28648,p2_datao_reg_16_ );
   nand U30072 ( n28650,p1_datao_reg_17_,n28547 );
   nor U30073 ( n28649,n28651,n28652 );
   nor U30074 ( n28652,n28159,n28653 );
   nor U30075 ( n28651,n28654,n28552 );
   not U30076 ( n28654,p2_datao_reg_17_ );
   nand U30077 ( n28656,p1_datao_reg_18_,n28547 );
   nor U30078 ( n28655,n28657,n28658 );
   nor U30079 ( n28658,n28161,n28659 );
   nor U30080 ( n28657,n28660,n28116 );
   not U30081 ( n28660,p2_datao_reg_18_ );
   nand U30082 ( n28662,p1_datao_reg_19_,n28547 );
   nor U30083 ( n28661,n28663,n28664 );
   nor U30084 ( n28664,n28160,n28665 );
   nor U30085 ( n28663,n28666,n28115 );
   not U30086 ( n28666,p2_datao_reg_19_ );
   nand U30087 ( n28668,p1_datao_reg_20_,n28547 );
   nor U30088 ( n28667,n28669,n28670 );
   nor U30089 ( n28670,n28162,n28671 );
   nor U30090 ( n28669,n28672,n28552 );
   not U30091 ( n28672,p2_datao_reg_20_ );
   nand U30092 ( n28674,p1_datao_reg_21_,n28130 );
   nor U30093 ( n28673,n28675,n28676 );
   nor U30094 ( n28676,n28159,n28677 );
   nor U30095 ( n28675,n28678,n28115 );
   not U30096 ( n28678,p2_datao_reg_21_ );
   nand U30097 ( n28680,p1_datao_reg_22_,n28130 );
   nor U30098 ( n28679,n28681,n28682 );
   nor U30099 ( n28682,n28161,n28683 );
   nor U30100 ( n28681,n28684,n28116 );
   not U30101 ( n28684,p2_datao_reg_22_ );
   nand U30102 ( n28686,p1_datao_reg_23_,n28130 );
   nor U30103 ( n28685,n28687,n28688 );
   nor U30104 ( n28688,n28160,n28689 );
   nor U30105 ( n28687,n28690,n28552 );
   not U30106 ( n28690,p2_datao_reg_23_ );
   nand U30107 ( n28692,p1_datao_reg_24_,n28130 );
   nor U30108 ( n28691,n28693,n28694 );
   nor U30109 ( n28694,n28162,n28695 );
   nor U30110 ( n28693,n28696,n28115 );
   not U30111 ( n28696,p2_datao_reg_24_ );
   nand U30112 ( n28698,p1_datao_reg_25_,n28130 );
   nor U30113 ( n28697,n28699,n28700 );
   nor U30114 ( n28700,n28159,n28701 );
   nor U30115 ( n28699,n28702,n28116 );
   not U30116 ( n28702,p2_datao_reg_25_ );
   nand U30117 ( n28704,p1_datao_reg_26_,n28130 );
   nor U30118 ( n28703,n28705,n28706 );
   nor U30119 ( n28706,n28161,n28707 );
   nor U30120 ( n28705,n28708,n28552 );
   not U30121 ( n28708,p2_datao_reg_26_ );
   nand U30122 ( n28710,p1_datao_reg_27_,n28130 );
   nor U30123 ( n28709,n28711,n28712 );
   nor U30124 ( n28712,n28160,n28713 );
   nor U30125 ( n28711,n28714,n28115 );
   not U30126 ( n28714,p2_datao_reg_27_ );
   nand U30127 ( n28716,p1_datao_reg_28_,n28130 );
   nor U30128 ( n28715,n28717,n28718 );
   nor U30129 ( n28718,n28162,n28719 );
   nor U30130 ( n28717,n28720,n28116 );
   not U30131 ( n28720,p2_datao_reg_28_ );
   nand U30132 ( n28722,p1_datao_reg_29_,n28130 );
   nor U30133 ( n28721,n28723,n28724 );
   nor U30134 ( n28724,n28159,n28725 );
   nor U30135 ( n28723,n28726,n28552 );
   not U30136 ( n28726,p2_datao_reg_29_ );
   nand U30137 ( n28728,p1_datao_reg_30_,n28130 );
   nor U30138 ( n28727,n28729,n28730 );
   nor U30139 ( n28730,n28161,n28731 );
   nor U30140 ( n28729,n28478,n28115 );
   not U30141 ( n28478,p2_datao_reg_30_ );
   nand U30142 ( n28733,p1_datao_reg_31_,n28547 );
   nor U30143 ( n28732,n28734,n28735 );
   nor U30144 ( n28735,n28160,n28736 );
   nor U30145 ( n28734,n28737,n28116 );
   nand U30146 ( n28552,n28132,n28160 );
   or U30147 ( n28738,n28739,n28740 );
   nor U30148 ( n28742,n28743,n28744 );
   or U30149 ( n28744,p3_be_n_reg_1_,p3_be_n_reg_2_ );
   nand U30150 ( n28743,n28745,n28746 );
   not U30151 ( n28746,p3_be_n_reg_3_ );
   nor U30152 ( n28745,p3_w_r_n_reg,p3_d_c_n_reg );
   nor U30153 ( n28741,n28747,n28748 );
   nand U30154 ( n28748,p3_m_io_n_reg,n28186 );
   not U30155 ( n53114,n28482 );
   nor U30156 ( n28482,n28740,p2_address_reg_29_ );
   or U30157 ( n28747,p3_ads_n_reg,p3_be_n_reg_0_ );
   nor U30158 ( n28749,n28547,n28740 );
   nand U30159 ( n28740,n28751,n28752 );
   nor U30160 ( n28752,n28753,n28754 );
   or U30161 ( n28754,p2_be_n_reg_1_,p2_be_n_reg_2_ );
   or U30162 ( n28753,p2_be_n_reg_3_,p2_d_c_n_reg );
   nor U30163 ( n28751,n28755,n28756 );
   nand U30164 ( n28756,p2_w_r_n_reg,p2_m_io_n_reg );
   or U30165 ( n28755,p2_ads_n_reg,p2_be_n_reg_0_ );
   not U30166 ( n28547,n28132 );
   nor U30167 ( n28758,n28759,n28760 );
   or U30168 ( n28760,p1_be_n_reg_0_,p1_be_n_reg_1_ );
   nand U30169 ( n28759,n28761,n28762 );
   not U30170 ( n28762,p1_be_n_reg_2_ );
   nor U30171 ( n28761,p1_d_c_n_reg,p1_be_n_reg_3_ );
   nor U30172 ( n28757,n28763,n28764 );
   nand U30173 ( n28764,p1_w_r_n_reg,p1_m_io_n_reg );
   or U30174 ( n28763,n28765,p1_ads_n_reg );
   nand U30175 ( n28767,p3_memoryfetch_reg,n28768 );
   nand U30176 ( n28766,n28769,n28770 );
   nand U30177 ( n28769,n28771,p3_state2_reg_2_ );
   nand U30178 ( n28773,n28768,p3_readrequest_reg );
   nand U30179 ( n28772,n28774,n28770 );
   not U30180 ( n28770,n28768 );
   nor U30181 ( n28768,n28775,n28776 );
   nand U30182 ( n28774,n28777,p3_state2_reg_2_ );
   nand U30183 ( n28779,p3_m_io_n_reg,n28376 );
   nand U30184 ( n28778,p3_memoryfetch_reg,n28781 );
   or U30185 ( n28783,n28784,n28785 );
   nand U30186 ( n28782,n28786,n28784 );
   nand U30187 ( n28784,n28787,n28788 );
   nand U30188 ( n28788,n28789,n28790 );
   nand U30189 ( n28789,n28791,n28792 );
   nand U30190 ( n28792,n28793,n28794 );
   nor U30191 ( n28787,n28795,n28776 );
   nand U30192 ( n28786,n28796,n28797 );
   nand U30193 ( n28797,p3_state2_reg_0_,n28798 );
   nand U30194 ( n28798,n28799,n28800 );
   nor U30195 ( n28800,n28801,n28802 );
   nor U30196 ( n28802,n28803,n28804 );
   nor U30197 ( n28803,n28805,n28806 );
   nor U30198 ( n28799,n28807,n28808 );
   nor U30199 ( n28807,n28809,n28810 );
   nand U30200 ( n28812,p3_more_reg,n28813 );
   or U30201 ( n28811,n28814,n28815 );
   or U30202 ( n28817,n28780,p3_readrequest_reg );
   nand U30203 ( n28816,p3_w_r_n_reg,n28376 );
   nor U30204 ( n28818,n28820,n28821 );
   nor U30205 ( n28821,n28822,n28823 );
   and U30206 ( n28820,n28822,p3_byteenable_reg_0_ );
   nand U30207 ( n28825,n28826,p3_reip_reg_0_ );
   nor U30208 ( n28824,n28827,n28828 );
   nor U30209 ( n28828,n28822,n28829 );
   nand U30210 ( n28829,n28830,n28831 );
   nand U30211 ( n28831,p3_reip_reg_0_,p3_datawidth_reg_0_ );
   nor U30212 ( n28830,p3_reip_reg_1_,p3_datawidth_reg_1_ );
   and U30213 ( n28827,n28822,p3_byteenable_reg_2_ );
   nand U30214 ( n28833,n28834,p3_instqueuerd_addr_reg_0_ );
   nand U30215 ( n28832,n28835,n28836 );
   nand U30216 ( n28835,n28837,n28838 );
   nand U30217 ( n28838,p3_state2_reg_1_,n28839 );
   nor U30218 ( n28837,n28840,n28841 );
   nor U30219 ( n28841,p3_instqueuerd_addr_reg_0_,n28842 );
   nor U30220 ( n28840,n28843,n28791 );
   nand U30221 ( n28845,n28834,p3_instqueuerd_addr_reg_1_ );
   nand U30222 ( n28844,n28846,n28836 );
   nand U30223 ( n28846,n28847,n28848 );
   nand U30224 ( n28848,n28849,n28850 );
   nor U30225 ( n28847,n28851,n28852 );
   nor U30226 ( n28852,n28853,n28791 );
   nor U30227 ( n28851,n28839,n28854 );
   or U30228 ( n28854,n28855,n28856 );
   nand U30229 ( n28858,n28834,p3_instqueuerd_addr_reg_2_ );
   nand U30230 ( n28857,n28859,n28836 );
   nand U30231 ( n28859,n28860,n28861 );
   nand U30232 ( n28861,n28850,n28862 );
   nor U30233 ( n28860,n28863,n28864 );
   and U30234 ( n28864,n28865,n28866 );
   nor U30235 ( n28863,n28839,n28867 );
   nand U30236 ( n28867,p3_state2_reg_1_,n28855 );
   xor U30237 ( n28855,p3_instaddrpointer_reg_31_,p3_instaddrpointer_reg_1_ );
   nand U30238 ( n28869,n28834,p3_instqueuerd_addr_reg_3_ );
   nand U30239 ( n28868,n28870,n28836 );
   nand U30240 ( n28870,n28871,n28872 );
   nand U30241 ( n28872,n28866,n28873 );
   nand U30242 ( n28871,n28850,n28874 );
   nand U30243 ( n28876,n28877,n28878 );
   nor U30244 ( n28877,n28879,n28791 );
   nor U30245 ( n28879,n28880,p3_instqueuerd_addr_reg_4_ );
   nor U30246 ( n28880,n28881,n28882 );
   nand U30247 ( n28882,p3_instqueuerd_addr_reg_1_,n28836 );
   not U30248 ( n28881,n28883 );
   nand U30249 ( n28875,n28834,p3_instqueuerd_addr_reg_4_ );
   not U30250 ( n28834,n28836 );
   nand U30251 ( n28836,n28884,n28885 );
   nand U30252 ( n28885,p3_state2_reg_3_,n28790 );
   nor U30253 ( n28884,n28886,n28887 );
   nor U30254 ( n28887,n28888,n28815 );
   nand U30255 ( n28890,p3_state2_reg_3_,n28891 );
   nand U30256 ( n28889,n28892,n28793 );
   nand U30257 ( n28894,n28895,p3_datawidth_reg_1_ );
   nand U30258 ( n28893,n28896,n28158 );
   nand U30259 ( n28896,n28898,n28899 );
   nand U30260 ( n28901,n28902,n28897 );
   nor U30261 ( n28902,bs16,n28903 );
   nand U30262 ( n28900,n28895,p3_datawidth_reg_0_ );
   nand U30263 ( n28905,p3_be_n_reg_0_,n28780 );
   nand U30264 ( n28904,p3_byteenable_reg_0_,n28781 );
   nand U30265 ( n28907,p3_be_n_reg_1_,n28780 );
   nand U30266 ( n28906,p3_byteenable_reg_1_,n28781 );
   nand U30267 ( n28909,p3_be_n_reg_2_,n28376 );
   nand U30268 ( n28908,p3_byteenable_reg_2_,n28781 );
   nand U30269 ( n28911,p3_be_n_reg_3_,n28376 );
   nand U30270 ( n28910,p3_byteenable_reg_3_,n28781 );
   nand U30271 ( n28913,p3_address_reg_29_,n28376 );
   nor U30272 ( n28912,n28914,n28915 );
   nor U30273 ( n28915,n28135,n28917 );
   nor U30274 ( n28914,n28918,n28919 );
   nand U30275 ( n28921,p3_address_reg_28_,n28376 );
   nor U30276 ( n28920,n28922,n28923 );
   nor U30277 ( n28923,n28919,n28136 );
   nor U30278 ( n28922,n28391,n28924 );
   nand U30279 ( n28926,p3_address_reg_27_,n28780 );
   nor U30280 ( n28925,n28927,n28928 );
   nor U30281 ( n28928,n28136,n28924 );
   nor U30282 ( n28927,n28918,n28929 );
   nand U30283 ( n28931,p3_address_reg_26_,n28376 );
   nor U30284 ( n28930,n28932,n28933 );
   nor U30285 ( n28933,n28916,n28929 );
   nor U30286 ( n28932,n28392,n28934 );
   nand U30287 ( n28936,p3_address_reg_25_,n28376 );
   nor U30288 ( n28935,n28937,n28938 );
   nor U30289 ( n28938,n28135,n28934 );
   nor U30290 ( n28937,n28391,n28939 );
   nand U30291 ( n28941,p3_address_reg_24_,n28376 );
   nor U30292 ( n28940,n28942,n28943 );
   nor U30293 ( n28943,n28136,n28939 );
   nor U30294 ( n28942,n28391,n28944 );
   nand U30295 ( n28946,p3_address_reg_23_,n28376 );
   nor U30296 ( n28945,n28947,n28948 );
   nor U30297 ( n28948,n28916,n28944 );
   nor U30298 ( n28947,n28918,n28949 );
   nand U30299 ( n28951,p3_address_reg_22_,n28376 );
   nor U30300 ( n28950,n28952,n28953 );
   nor U30301 ( n28953,n28916,n28949 );
   nor U30302 ( n28952,n28392,n28954 );
   nand U30303 ( n28956,p3_address_reg_21_,n28376 );
   nor U30304 ( n28955,n28957,n28958 );
   nor U30305 ( n28958,n28135,n28954 );
   nor U30306 ( n28957,n28391,n28959 );
   nand U30307 ( n28961,p3_address_reg_20_,n28780 );
   nor U30308 ( n28960,n28962,n28963 );
   nor U30309 ( n28963,n28136,n28959 );
   nor U30310 ( n28962,n28918,n28964 );
   nand U30311 ( n28966,p3_address_reg_19_,n28376 );
   nor U30312 ( n28965,n28967,n28968 );
   nor U30313 ( n28968,n28916,n28964 );
   nor U30314 ( n28967,n28392,n28969 );
   nand U30315 ( n28971,p3_address_reg_18_,n28780 );
   nor U30316 ( n28970,n28972,n28973 );
   nor U30317 ( n28973,n28135,n28969 );
   nor U30318 ( n28972,n28391,n28974 );
   nand U30319 ( n28976,p3_address_reg_17_,n28376 );
   nor U30320 ( n28975,n28977,n28978 );
   nor U30321 ( n28978,n28136,n28974 );
   nor U30322 ( n28977,n28918,n28979 );
   nand U30323 ( n28981,p3_address_reg_16_,n28376 );
   nor U30324 ( n28980,n28982,n28983 );
   nor U30325 ( n28983,n28916,n28979 );
   nor U30326 ( n28982,n28392,n28984 );
   nand U30327 ( n28986,p3_address_reg_15_,n28376 );
   nor U30328 ( n28985,n28987,n28988 );
   nor U30329 ( n28988,n28135,n28984 );
   nor U30330 ( n28987,n28392,n28989 );
   nand U30331 ( n28991,p3_address_reg_14_,n28376 );
   nor U30332 ( n28990,n28992,n28993 );
   nor U30333 ( n28993,n28136,n28989 );
   nor U30334 ( n28992,n28392,n28994 );
   nand U30335 ( n28996,p3_address_reg_13_,n28376 );
   nor U30336 ( n28995,n28997,n28998 );
   nor U30337 ( n28998,n28135,n28994 );
   nor U30338 ( n28997,n28918,n28999 );
   nand U30339 ( n29001,p3_address_reg_12_,n28780 );
   nor U30340 ( n29000,n29002,n29003 );
   nor U30341 ( n29003,n28916,n28999 );
   nor U30342 ( n29002,n28391,n29004 );
   nand U30343 ( n29006,p3_address_reg_11_,n28376 );
   nor U30344 ( n29005,n29007,n29008 );
   nor U30345 ( n29008,n28916,n29004 );
   nor U30346 ( n29007,n28391,n29009 );
   nand U30347 ( n29011,p3_address_reg_10_,n28376 );
   nor U30348 ( n29010,n29012,n29013 );
   nor U30349 ( n29013,n28135,n29009 );
   nor U30350 ( n29012,n28918,n29014 );
   nand U30351 ( n29016,p3_address_reg_9_,n28780 );
   nor U30352 ( n29015,n29017,n29018 );
   nor U30353 ( n29018,n28136,n29014 );
   nor U30354 ( n29017,n28392,n29019 );
   nand U30355 ( n29021,p3_address_reg_8_,n28780 );
   nor U30356 ( n29020,n29022,n29023 );
   nor U30357 ( n29023,n28916,n29019 );
   nor U30358 ( n29022,n28391,n29024 );
   nand U30359 ( n29026,p3_address_reg_7_,n28376 );
   nor U30360 ( n29025,n29027,n29028 );
   nor U30361 ( n29028,n28135,n29024 );
   nor U30362 ( n29027,n28918,n29029 );
   nand U30363 ( n29031,p3_address_reg_6_,n28780 );
   nor U30364 ( n29030,n29032,n29033 );
   nor U30365 ( n29033,n28136,n29029 );
   nor U30366 ( n29032,n28392,n29034 );
   nand U30367 ( n29036,p3_address_reg_5_,n28376 );
   nor U30368 ( n29035,n29037,n29038 );
   nor U30369 ( n29038,n28916,n29034 );
   nor U30370 ( n29037,n28391,n29039 );
   nand U30371 ( n29041,p3_address_reg_4_,n28780 );
   nor U30372 ( n29040,n29042,n29043 );
   nor U30373 ( n29043,n28135,n29039 );
   nor U30374 ( n29042,n28918,n29044 );
   nand U30375 ( n29046,p3_address_reg_3_,n28780 );
   nor U30376 ( n29045,n29047,n29048 );
   nor U30377 ( n29048,n28136,n29044 );
   nor U30378 ( n29047,n28392,n29049 );
   nand U30379 ( n29051,p3_address_reg_2_,n28780 );
   nor U30380 ( n29050,n29052,n29053 );
   nor U30381 ( n29053,n28916,n29049 );
   nor U30382 ( n29052,n28391,n29054 );
   nand U30383 ( n29056,p3_address_reg_1_,n28376 );
   nor U30384 ( n29055,n29057,n29058 );
   nor U30385 ( n29058,n28135,n29054 );
   nor U30386 ( n29057,n28918,n29059 );
   nand U30387 ( n29061,p3_address_reg_0_,n28780 );
   nor U30388 ( n29060,n29062,n29063 );
   nor U30389 ( n29063,n28136,n29059 );
   nor U30390 ( n29062,n29064,n28392 );
   not U30391 ( n28918,n29065 );
   nand U30392 ( n29067,n29068,n29069 );
   nor U30393 ( n29069,n29070,n29071 );
   nor U30394 ( n29071,n29072,n29073 );
   nor U30395 ( n29073,p3_requestpending_reg,n28899 );
   nor U30396 ( n29070,n29074,n29075 );
   nor U30397 ( n29068,n29076,n29077 );
   nor U30398 ( n29076,p3_requestpending_reg,hold );
   nor U30399 ( n29066,n29065,n29078 );
   nor U30400 ( n29078,n29079,n29080 );
   nor U30401 ( n29079,n29072,n29081 );
   nand U30402 ( n29081,n29082,n29083 );
   nand U30403 ( n29083,n29075,n29077 );
   nand U30404 ( n29082,hold,p3_state_reg_0_ );
   nor U30405 ( n29072,n29074,n28794 );
   nor U30406 ( n29065,n29080,n28780 );
   nor U30407 ( n29085,n29086,n29087 );
   nand U30408 ( n29087,n29088,n28135 );
   nand U30409 ( n28916,n28781,n29080 );
   nand U30410 ( n29088,n29089,p3_state_reg_1_ );
   nor U30411 ( n29089,n29090,n29091 );
   nor U30412 ( n29091,n28801,n29092 );
   nand U30413 ( n29092,n29093,n28785 );
   nor U30414 ( n29090,n29094,n29080 );
   nor U30415 ( n29094,n29095,n29077 );
   nor U30416 ( n29095,n28801,n29093 );
   nor U30417 ( n29086,n28899,n29096 );
   nand U30418 ( n29096,p3_state_reg_0_,p3_requestpending_reg );
   not U30419 ( n28899,n28903 );
   nor U30420 ( n29084,n29097,n29098 );
   nor U30421 ( n29098,n28780,n28794 );
   nor U30422 ( n29097,n29099,n29080 );
   nor U30423 ( n29099,n29100,n29101 );
   and U30424 ( n29100,n29074,n29102 );
   nand U30425 ( n29104,n29101,na );
   nor U30426 ( n29103,n29105,n29106 );
   nor U30427 ( n29106,p3_state_reg_2_,n29107 );
   nor U30428 ( n29107,n29077,n29108 );
   nand U30429 ( n29108,p3_requestpending_reg,n29109 );
   nand U30430 ( n29109,n28801,p3_state_reg_1_ );
   nor U30431 ( n29105,n29102,n29110 );
   nand U30432 ( n29110,n29111,n29112 );
   nand U30433 ( n29112,n29074,n29080 );
   not U30434 ( n29080,p3_state_reg_2_ );
   nand U30435 ( n29111,p3_state_reg_1_,n29077 );
   nor U30436 ( n29102,n28785,hold );
   not U30437 ( n28785,p3_requestpending_reg );
   nor U30438 ( n53115,n28157,n29113 );
   nor U30439 ( n53116,n28157,n29116 );
   nor U30440 ( n53117,n28897,n29117 );
   nor U30441 ( n53118,n28158,n29118 );
   nor U30442 ( n53119,n28158,n29119 );
   nor U30443 ( n53120,n28157,n29120 );
   nor U30444 ( n53121,n28897,n29121 );
   nor U30445 ( n53122,n28158,n29122 );
   nor U30446 ( n53123,n28157,n29123 );
   nor U30447 ( n53124,n28897,n29124 );
   nor U30448 ( n53125,n28157,n29125 );
   nor U30449 ( n53126,n28897,n29126 );
   nor U30450 ( n53127,n28897,n29127 );
   nor U30451 ( n53128,n28157,n29128 );
   nor U30452 ( n53129,n28158,n29129 );
   nor U30453 ( n53130,n28897,n29130 );
   nor U30454 ( n53131,n28157,n29131 );
   nor U30455 ( n53132,n28158,n29132 );
   nor U30456 ( n53133,n28157,n29133 );
   nor U30457 ( n53134,n28897,n29134 );
   nor U30458 ( n53135,n28158,n29135 );
   nor U30459 ( n53136,n28157,n29136 );
   nor U30460 ( n53137,n28897,n29137 );
   nor U30461 ( n53138,n28158,n29138 );
   nor U30462 ( n53139,n28157,n29139 );
   nor U30463 ( n53140,n28897,n29140 );
   nor U30464 ( n53141,n28158,n29141 );
   nor U30465 ( n53142,n28158,n29142 );
   nand U30466 ( n29144,p3_state2_reg_2_,n29145 );
   nand U30467 ( n29145,n28892,p3_state2_reg_1_ );
   nor U30468 ( n29143,n29146,n29147 );
   nor U30469 ( n29147,n28790,n29148 );
   nand U30470 ( n29148,n29149,n28794 );
   nor U30471 ( n29146,p3_state2_reg_0_,n29150 );
   nand U30472 ( n29150,p3_statebs16_reg,p3_state2_reg_1_ );
   nor U30473 ( n29152,n29153,n29154 );
   nor U30474 ( n29154,n28891,n29155 );
   nand U30475 ( n29155,n28866,n28794 );
   not U30476 ( n28891,n28892 );
   nor U30477 ( n28892,n28790,n29156 );
   nor U30478 ( n29151,n29157,n29158 );
   nor U30479 ( n29158,n29156,n28815 );
   nor U30480 ( n29157,n29159,n28856 );
   and U30481 ( n29159,n29160,n29161 );
   nor U30482 ( n29163,n29164,n29165 );
   nand U30483 ( n29165,n29160,n29166 );
   not U30484 ( n29166,n29167 );
   nand U30485 ( n29160,n29168,n28801 );
   nor U30486 ( n29168,p3_state2_reg_2_,n28790 );
   nor U30487 ( n29164,n29169,n29170 );
   not U30488 ( n29169,n29171 );
   nor U30489 ( n29162,n29172,n29173 );
   nand U30490 ( n29173,n29174,n29175 );
   nand U30491 ( n29175,n29176,n28790 );
   nor U30492 ( n29176,n29156,n29177 );
   nor U30493 ( n29177,n28842,n28796 );
   not U30494 ( n28842,n28850 );
   nand U30495 ( n29174,n29156,p3_state2_reg_0_ );
   not U30496 ( n29156,n29161 );
   nand U30497 ( n29161,n29178,n29179 );
   nand U30498 ( n29179,n29180,n29181 );
   nand U30499 ( n29180,n28801,n28793 );
   nand U30500 ( n29178,p3_state2_reg_0_,n29182 );
   nand U30501 ( n29182,n29183,n29184 );
   nor U30502 ( n29183,p3_state2_reg_1_,n29185 );
   nor U30503 ( n29185,n29186,n29187 );
   nor U30504 ( n29172,n29184,n28815 );
   and U30505 ( n29184,n29188,n29189 );
   nor U30506 ( n29189,n29190,n29191 );
   nand U30507 ( n29191,n29192,n29193 );
   nand U30508 ( n29193,n29194,n29195 );
   nand U30509 ( n29192,n28878,n29196 );
   nand U30510 ( n29196,n29197,n29198 );
   nand U30511 ( n29198,n28883,p3_instqueuerd_addr_reg_1_ );
   nand U30512 ( n29190,n29199,n28814 );
   nand U30513 ( n28814,n29200,n29201 );
   nand U30514 ( n29201,n29202,n29203 );
   nor U30515 ( n29203,n29204,n29205 );
   nand U30516 ( n29205,n29206,n29207 );
   nand U30517 ( n29207,n29208,n29209 );
   nand U30518 ( n29206,n29210,n29211 );
   nand U30519 ( n29204,n29212,n29213 );
   nand U30520 ( n29213,n29214,n29209 );
   nand U30521 ( n29212,n29215,n29216 );
   nor U30522 ( n29202,n29217,n29218 );
   nand U30523 ( n29218,n29219,n29220 );
   nand U30524 ( n29220,n29221,n29209 );
   nand U30525 ( n29219,n29222,n29211 );
   nor U30526 ( n29217,n29223,n29224 );
   nand U30527 ( n29199,n29225,n29226 );
   or U30528 ( n29226,p3_more_reg,p3_flush_reg );
   not U30529 ( n29225,n29200 );
   nor U30530 ( n29188,n29227,n29228 );
   nand U30531 ( n29228,n29229,n29230 );
   nand U30532 ( n29230,n29231,n29232 );
   nand U30533 ( n29231,n29233,n29234 );
   nand U30534 ( n29234,n29195,n29235 );
   nand U30535 ( n29233,n29236,n29237 );
   or U30536 ( n29237,n29195,n29235 );
   nand U30537 ( n29195,n29238,n29239 );
   nand U30538 ( n29239,n28888,p3_instqueuerd_addr_reg_3_ );
   nand U30539 ( n29238,n28873,n29240 );
   nand U30540 ( n28873,n29241,n29242 );
   nor U30541 ( n29242,n29243,n29244 );
   nor U30542 ( n29244,n29245,n29246 );
   nor U30543 ( n29243,n29247,n29248 );
   nand U30544 ( n29248,n29249,n29250 );
   not U30545 ( n29250,n28777 );
   nand U30546 ( n29249,n29251,n29245 );
   nor U30547 ( n29251,n29252,n29253 );
   nor U30548 ( n29253,n29254,n29255 );
   nand U30549 ( n29255,n29256,n29257 );
   nor U30550 ( n29252,p3_instqueuerd_addr_reg_3_,n29256 );
   nor U30551 ( n29241,n29258,n29259 );
   nor U30552 ( n29259,n29260,n29261 );
   nor U30553 ( n29258,n29262,n29254 );
   nor U30554 ( n29262,n29263,n29264 );
   nand U30555 ( n29264,n29265,n29266 );
   nand U30556 ( n29266,n29267,n29268 );
   nand U30557 ( n29268,n29269,n29270 );
   not U30558 ( n29270,n29271 );
   nor U30559 ( n29269,n29210,n29272 );
   nand U30560 ( n29265,n29273,n29274 );
   and U30561 ( n29263,n29275,n29272 );
   nor U30562 ( n29236,n29276,n29277 );
   nor U30563 ( n29277,n29278,n29194 );
   nor U30564 ( n29276,n29279,n29280 );
   nand U30565 ( n29280,n29281,n29282 );
   nand U30566 ( n29282,n29194,n29278 );
   nand U30567 ( n29194,n29283,n29284 );
   nand U30568 ( n29284,n28888,p3_instqueuerd_addr_reg_2_ );
   nand U30569 ( n29283,n28865,n29240 );
   nand U30570 ( n28865,n29285,n29286 );
   nor U30571 ( n29286,n29287,n29288 );
   nor U30572 ( n29288,p3_instqueuerd_addr_reg_2_,n29246 );
   nand U30573 ( n29246,p3_instqueuerd_addr_reg_1_,n29289 );
   nor U30574 ( n29287,n29290,n29257 );
   nor U30575 ( n29290,n29291,n29292 );
   nor U30576 ( n29292,p3_instqueuerd_addr_reg_1_,n29293 );
   nor U30577 ( n29291,n29294,n29295 );
   nor U30578 ( n29295,n29272,n29273 );
   nand U30579 ( n29273,n29296,n29297 );
   not U30580 ( n29297,n29298 );
   nor U30581 ( n29296,n29299,n29300 );
   nor U30582 ( n29300,n28777,n29301 );
   nor U30583 ( n29299,n29302,n29303 );
   nand U30584 ( n29303,n29304,n29305 );
   nand U30585 ( n29305,n29306,n29307 );
   nand U30586 ( n29307,n29308,n29309 );
   nor U30587 ( n29285,n29310,n29311 );
   nor U30588 ( n29311,n29312,n29260 );
   nor U30589 ( n29310,n28862,n29313 );
   or U30590 ( n29313,n29247,n28777 );
   nor U30591 ( n28777,n29314,n29315 );
   nand U30592 ( n29281,n29316,n29317 );
   nand U30593 ( n29317,n29318,p3_instqueuewr_addr_reg_0_ );
   nor U30594 ( n29318,n29319,n29320 );
   nor U30595 ( n29320,n29275,n29240 );
   nor U30596 ( n29319,n28888,n28843 );
   not U30597 ( n28843,n29321 );
   nand U30598 ( n29279,n29322,n29323 );
   nand U30599 ( n29323,n28888,n29324 );
   nand U30600 ( n29324,n29256,n29325 );
   nand U30601 ( n29325,p3_instqueuerd_addr_reg_1_,n29326 );
   nand U30602 ( n29322,n29327,n29240 );
   nor U30603 ( n29327,n28853,n29328 );
   nor U30604 ( n29328,n29321,n29326 );
   nand U30605 ( n29321,n29329,n29330 );
   nand U30606 ( n29330,n29331,n29275 );
   nand U30607 ( n29331,n29332,n29333 );
   nor U30608 ( n29333,n29208,n29334 );
   nor U30609 ( n29332,n29335,n29336 );
   nand U30610 ( n29329,p3_instqueuerd_addr_reg_0_,n29337 );
   nand U30611 ( n29337,n29293,n29260 );
   and U30612 ( n28853,n29338,n29339 );
   nand U30613 ( n29339,n29340,n29341 );
   or U30614 ( n29340,n29289,n28878 );
   nand U30615 ( n29289,n29293,n29342 );
   nand U30616 ( n29342,p3_instqueuerd_addr_reg_0_,n29343 );
   nand U30617 ( n29343,n29344,n29345 );
   nand U30618 ( n29345,n29346,n29315 );
   not U30619 ( n29344,n29336 );
   and U30620 ( n29293,n29347,n29348 );
   nand U30621 ( n29348,n29349,n29350 );
   and U30622 ( n29347,n29351,n29352 );
   nor U30623 ( n29338,n29353,n29354 );
   nor U30624 ( n29354,n29355,n29356 );
   nor U30625 ( n29355,n29334,n29336 );
   nand U30626 ( n29336,n29357,n29358 );
   nor U30627 ( n29358,n29359,n29360 );
   nor U30628 ( n29360,n29361,n29302 );
   and U30629 ( n29361,n29362,n29306 );
   nor U30630 ( n29357,n29298,n29272 );
   nand U30631 ( n29298,n29363,n29364 );
   nand U30632 ( n29364,n29365,n29366 );
   nor U30633 ( n29353,n29367,n29368 );
   nor U30634 ( n29367,n29335,n29208 );
   nand U30635 ( n29229,n28888,p3_instqueuerd_addr_reg_4_ );
   not U30636 ( n28888,n29240 );
   nand U30637 ( n29240,n29369,n29370 );
   nor U30638 ( n29370,n29371,n29372 );
   nor U30639 ( n29372,n29373,n29209 );
   nor U30640 ( n29371,n29374,n29375 );
   nand U30641 ( n29375,n28809,n28794 );
   nor U30642 ( n29369,n29376,n29377 );
   nor U30643 ( n29379,n29380,n29381 );
   nand U30644 ( n29381,n29382,n29383 );
   nand U30645 ( n29383,n29384,n29385 );
   nand U30646 ( n29382,p3_instqueue_reg_15__7_,n29386 );
   nor U30647 ( n29380,n29387,n28190 );
   nor U30648 ( n29378,n29389,n29390 );
   nor U30649 ( n29390,n29391,n29392 );
   nor U30650 ( n29389,n29393,n28191 );
   nor U30651 ( n29396,n29397,n29398 );
   nand U30652 ( n29398,n29399,n29400 );
   nand U30653 ( n29400,n29401,n29384 );
   nand U30654 ( n29399,p3_instqueue_reg_15__6_,n29386 );
   nor U30655 ( n29397,n29387,n28195 );
   nor U30656 ( n29395,n29403,n29404 );
   nor U30657 ( n29404,n29391,n29405 );
   nor U30658 ( n29403,n29393,n28196 );
   nor U30659 ( n29408,n29409,n29410 );
   nand U30660 ( n29410,n29411,n29412 );
   nand U30661 ( n29412,n29413,n29384 );
   nand U30662 ( n29411,p3_instqueue_reg_15__5_,n29386 );
   nor U30663 ( n29409,n29387,n28201 );
   nor U30664 ( n29407,n29415,n29416 );
   nor U30665 ( n29416,n29391,n29417 );
   nor U30666 ( n29415,n29393,n28202 );
   nor U30667 ( n29420,n29421,n29422 );
   nand U30668 ( n29422,n29423,n29424 );
   nand U30669 ( n29424,n29425,n29384 );
   nand U30670 ( n29423,p3_instqueue_reg_15__4_,n29386 );
   nor U30671 ( n29421,n29387,n28208 );
   nor U30672 ( n29419,n29427,n29428 );
   nor U30673 ( n29428,n29391,n29429 );
   nor U30674 ( n29427,n29393,n28209 );
   nor U30675 ( n29432,n29433,n29434 );
   nand U30676 ( n29434,n29435,n29436 );
   nand U30677 ( n29436,n29437,n29384 );
   nand U30678 ( n29435,p3_instqueue_reg_15__3_,n29386 );
   nor U30679 ( n29433,n29387,n28216 );
   nor U30680 ( n29431,n29439,n29440 );
   nor U30681 ( n29440,n29391,n29441 );
   nor U30682 ( n29439,n29393,n28217 );
   nor U30683 ( n29444,n29445,n29446 );
   nand U30684 ( n29446,n29447,n29448 );
   nand U30685 ( n29448,n29449,n29384 );
   nand U30686 ( n29447,p3_instqueue_reg_15__2_,n29386 );
   nor U30687 ( n29445,n29387,n28228 );
   nor U30688 ( n29443,n29451,n29452 );
   nor U30689 ( n29452,n29391,n29453 );
   nor U30690 ( n29451,n29393,n28229 );
   nor U30691 ( n29456,n29457,n29458 );
   nand U30692 ( n29458,n29459,n29460 );
   nand U30693 ( n29460,n29461,n29384 );
   nand U30694 ( n29459,p3_instqueue_reg_15__1_,n29386 );
   nor U30695 ( n29457,n29387,n28246 );
   nor U30696 ( n29455,n29463,n29464 );
   nor U30697 ( n29464,n29391,n29465 );
   nor U30698 ( n29463,n29393,n28247 );
   nor U30699 ( n29468,n29469,n29470 );
   nand U30700 ( n29470,n29471,n29472 );
   nand U30701 ( n29472,n29473,n29384 );
   nor U30702 ( n29384,n29474,n29475 );
   nand U30703 ( n29471,p3_instqueue_reg_15__0_,n29386 );
   nand U30704 ( n29386,n29476,n29477 );
   nand U30705 ( n29477,n29475,n29478 );
   nand U30706 ( n29478,n29479,n29480 );
   nand U30707 ( n29480,n29387,n29391 );
   and U30708 ( n29475,n29393,n29481 );
   nand U30709 ( n29481,n29482,n29483 );
   nand U30710 ( n29476,n29484,n29485 );
   nand U30711 ( n29485,n29486,n29487 );
   nor U30712 ( n29469,n29387,n28270 );
   nand U30713 ( n29387,n29489,n29490 );
   nor U30714 ( n29467,n29491,n29492 );
   nor U30715 ( n29492,n29391,n29493 );
   nand U30716 ( n29391,n29494,n29495 );
   nor U30717 ( n29491,n29393,n28271 );
   not U30718 ( n29393,n29486 );
   nor U30719 ( n29486,n29497,n29235 );
   nor U30720 ( n29499,n29500,n29501 );
   nand U30721 ( n29501,n29502,n29503 );
   nand U30722 ( n29503,n29504,n29385 );
   nand U30723 ( n29502,p3_instqueue_reg_14__7_,n29505 );
   nor U30724 ( n29500,n29388,n29506 );
   nor U30725 ( n29498,n29507,n29508 );
   nor U30726 ( n29508,n29392,n29509 );
   nor U30727 ( n29507,n29394,n29510 );
   nor U30728 ( n29512,n29513,n29514 );
   nand U30729 ( n29514,n29515,n29516 );
   nand U30730 ( n29516,n29504,n29401 );
   nand U30731 ( n29515,p3_instqueue_reg_14__6_,n29505 );
   nor U30732 ( n29513,n29402,n29506 );
   nor U30733 ( n29511,n29517,n29518 );
   nor U30734 ( n29518,n29405,n29509 );
   nor U30735 ( n29517,n29406,n29510 );
   nor U30736 ( n29520,n29521,n29522 );
   nand U30737 ( n29522,n29523,n29524 );
   nand U30738 ( n29524,n29504,n29413 );
   nand U30739 ( n29523,p3_instqueue_reg_14__5_,n29505 );
   nor U30740 ( n29521,n29414,n29506 );
   nor U30741 ( n29519,n29525,n29526 );
   nor U30742 ( n29526,n29417,n29509 );
   nor U30743 ( n29525,n29418,n29510 );
   nor U30744 ( n29528,n29529,n29530 );
   nand U30745 ( n29530,n29531,n29532 );
   nand U30746 ( n29532,n29504,n29425 );
   nand U30747 ( n29531,p3_instqueue_reg_14__4_,n29505 );
   nor U30748 ( n29529,n29426,n29506 );
   nor U30749 ( n29527,n29533,n29534 );
   nor U30750 ( n29534,n29429,n29509 );
   nor U30751 ( n29533,n29430,n29510 );
   nor U30752 ( n29536,n29537,n29538 );
   nand U30753 ( n29538,n29539,n29540 );
   nand U30754 ( n29540,n29504,n29437 );
   nand U30755 ( n29539,p3_instqueue_reg_14__3_,n29505 );
   nor U30756 ( n29537,n29438,n29506 );
   nor U30757 ( n29535,n29541,n29542 );
   nor U30758 ( n29542,n29441,n29509 );
   nor U30759 ( n29541,n29442,n29510 );
   nor U30760 ( n29544,n29545,n29546 );
   nand U30761 ( n29546,n29547,n29548 );
   nand U30762 ( n29548,n29504,n29449 );
   nand U30763 ( n29547,p3_instqueue_reg_14__2_,n29505 );
   nor U30764 ( n29545,n29450,n29506 );
   nor U30765 ( n29543,n29549,n29550 );
   nor U30766 ( n29550,n29453,n29509 );
   nor U30767 ( n29549,n29454,n29510 );
   nor U30768 ( n29552,n29553,n29554 );
   nand U30769 ( n29554,n29555,n29556 );
   nand U30770 ( n29556,n29504,n29461 );
   nand U30771 ( n29555,p3_instqueue_reg_14__1_,n29505 );
   nor U30772 ( n29553,n29462,n29506 );
   nor U30773 ( n29551,n29557,n29558 );
   nor U30774 ( n29558,n29465,n29509 );
   nor U30775 ( n29557,n29466,n29510 );
   nor U30776 ( n29560,n29561,n29562 );
   nand U30777 ( n29562,n29563,n29564 );
   nand U30778 ( n29564,n29504,n29473 );
   and U30779 ( n29504,n29565,n29566 );
   nor U30780 ( n29565,n29474,n29567 );
   nand U30781 ( n29563,p3_instqueue_reg_14__0_,n29505 );
   nand U30782 ( n29505,n29568,n29569 );
   nand U30783 ( n29569,n29567,n29566 );
   nand U30784 ( n29566,n29479,n29570 );
   nand U30785 ( n29570,n29506,n29509 );
   and U30786 ( n29567,n29510,n29571 );
   nand U30787 ( n29571,n29572,n29483 );
   nand U30788 ( n29568,n29484,n29573 );
   or U30789 ( n29573,n29510,n28350 );
   nor U30790 ( n29561,n29488,n29506 );
   nand U30791 ( n29506,n29575,n29489 );
   nor U30792 ( n29559,n29576,n29577 );
   nor U30793 ( n29577,n29493,n29509 );
   nand U30794 ( n29509,n29578,n29495 );
   nor U30795 ( n29576,n29496,n29510 );
   nand U30796 ( n29510,n29579,n29580 );
   nor U30797 ( n29582,n29583,n29584 );
   nand U30798 ( n29584,n29585,n29586 );
   nand U30799 ( n29586,n29587,n29385 );
   nand U30800 ( n29585,p3_instqueue_reg_13__7_,n29588 );
   nor U30801 ( n29583,n29388,n29589 );
   nor U30802 ( n29581,n29590,n29591 );
   nor U30803 ( n29591,n29392,n29592 );
   nor U30804 ( n29590,n29394,n29593 );
   nor U30805 ( n29595,n29596,n29597 );
   nand U30806 ( n29597,n29598,n29599 );
   nand U30807 ( n29599,n29587,n29401 );
   nand U30808 ( n29598,p3_instqueue_reg_13__6_,n29588 );
   nor U30809 ( n29596,n29402,n29589 );
   nor U30810 ( n29594,n29600,n29601 );
   nor U30811 ( n29601,n29405,n29592 );
   nor U30812 ( n29600,n29406,n29593 );
   nor U30813 ( n29603,n29604,n29605 );
   nand U30814 ( n29605,n29606,n29607 );
   nand U30815 ( n29607,n29587,n29413 );
   nand U30816 ( n29606,p3_instqueue_reg_13__5_,n29588 );
   nor U30817 ( n29604,n29414,n29589 );
   nor U30818 ( n29602,n29608,n29609 );
   nor U30819 ( n29609,n29417,n29592 );
   nor U30820 ( n29608,n29418,n29593 );
   nor U30821 ( n29611,n29612,n29613 );
   nand U30822 ( n29613,n29614,n29615 );
   nand U30823 ( n29615,n29587,n29425 );
   nand U30824 ( n29614,p3_instqueue_reg_13__4_,n29588 );
   nor U30825 ( n29612,n29426,n29589 );
   nor U30826 ( n29610,n29616,n29617 );
   nor U30827 ( n29617,n29429,n29592 );
   nor U30828 ( n29616,n29430,n29593 );
   nor U30829 ( n29619,n29620,n29621 );
   nand U30830 ( n29621,n29622,n29623 );
   nand U30831 ( n29623,n29587,n29437 );
   nand U30832 ( n29622,p3_instqueue_reg_13__3_,n29588 );
   nor U30833 ( n29620,n29438,n29589 );
   nor U30834 ( n29618,n29624,n29625 );
   nor U30835 ( n29625,n29441,n29592 );
   nor U30836 ( n29624,n29442,n29593 );
   nor U30837 ( n29627,n29628,n29629 );
   nand U30838 ( n29629,n29630,n29631 );
   nand U30839 ( n29631,n29587,n29449 );
   nand U30840 ( n29630,p3_instqueue_reg_13__2_,n29588 );
   nor U30841 ( n29628,n29450,n29589 );
   nor U30842 ( n29626,n29632,n29633 );
   nor U30843 ( n29633,n29453,n29592 );
   nor U30844 ( n29632,n29454,n29593 );
   nor U30845 ( n29635,n29636,n29637 );
   nand U30846 ( n29637,n29638,n29639 );
   nand U30847 ( n29639,n29587,n29461 );
   nand U30848 ( n29638,p3_instqueue_reg_13__1_,n29588 );
   nor U30849 ( n29636,n29462,n29589 );
   nor U30850 ( n29634,n29640,n29641 );
   nor U30851 ( n29641,n29465,n29592 );
   nor U30852 ( n29640,n29466,n29593 );
   nor U30853 ( n29643,n29644,n29645 );
   nand U30854 ( n29645,n29646,n29647 );
   nand U30855 ( n29647,n29587,n29473 );
   and U30856 ( n29587,n29648,n29649 );
   nor U30857 ( n29648,n29474,n29650 );
   nand U30858 ( n29646,p3_instqueue_reg_13__0_,n29588 );
   nand U30859 ( n29588,n29651,n29652 );
   nand U30860 ( n29652,n29650,n29649 );
   nand U30861 ( n29649,n29479,n29653 );
   nand U30862 ( n29653,n29589,n29592 );
   and U30863 ( n29650,n29593,n29654 );
   nand U30864 ( n29654,n29655,n29483 );
   nand U30865 ( n29651,n29484,n29656 );
   or U30866 ( n29656,n29593,n28350 );
   nor U30867 ( n29644,n29488,n29589 );
   nand U30868 ( n29589,n29657,n29489 );
   nor U30869 ( n29642,n29658,n29659 );
   nor U30870 ( n29659,n29493,n29592 );
   nand U30871 ( n29592,n29660,n29495 );
   nor U30872 ( n29658,n29496,n29593 );
   nand U30873 ( n29593,n29661,n29580 );
   nor U30874 ( n29663,n29664,n29665 );
   nand U30875 ( n29665,n29666,n29667 );
   nand U30876 ( n29667,n29668,n29385 );
   nand U30877 ( n29666,p3_instqueue_reg_12__7_,n29669 );
   nor U30878 ( n29664,n29388,n29670 );
   nor U30879 ( n29662,n29671,n29672 );
   nor U30880 ( n29672,n29392,n29673 );
   nor U30881 ( n29671,n29394,n29674 );
   nor U30882 ( n29676,n29677,n29678 );
   nand U30883 ( n29678,n29679,n29680 );
   nand U30884 ( n29680,n29668,n29401 );
   nand U30885 ( n29679,p3_instqueue_reg_12__6_,n29669 );
   nor U30886 ( n29677,n29402,n29670 );
   nor U30887 ( n29675,n29681,n29682 );
   nor U30888 ( n29682,n29405,n29673 );
   nor U30889 ( n29681,n29406,n29674 );
   nor U30890 ( n29684,n29685,n29686 );
   nand U30891 ( n29686,n29687,n29688 );
   nand U30892 ( n29688,n29668,n29413 );
   nand U30893 ( n29687,p3_instqueue_reg_12__5_,n29669 );
   nor U30894 ( n29685,n29414,n29670 );
   nor U30895 ( n29683,n29689,n29690 );
   nor U30896 ( n29690,n29417,n29673 );
   nor U30897 ( n29689,n29418,n29674 );
   nor U30898 ( n29692,n29693,n29694 );
   nand U30899 ( n29694,n29695,n29696 );
   nand U30900 ( n29696,n29668,n29425 );
   nand U30901 ( n29695,p3_instqueue_reg_12__4_,n29669 );
   nor U30902 ( n29693,n29426,n29670 );
   nor U30903 ( n29691,n29697,n29698 );
   nor U30904 ( n29698,n29429,n29673 );
   nor U30905 ( n29697,n29430,n29674 );
   nor U30906 ( n29700,n29701,n29702 );
   nand U30907 ( n29702,n29703,n29704 );
   nand U30908 ( n29704,n29668,n29437 );
   nand U30909 ( n29703,p3_instqueue_reg_12__3_,n29669 );
   nor U30910 ( n29701,n29438,n29670 );
   nor U30911 ( n29699,n29705,n29706 );
   nor U30912 ( n29706,n29441,n29673 );
   nor U30913 ( n29705,n29442,n29674 );
   nor U30914 ( n29708,n29709,n29710 );
   nand U30915 ( n29710,n29711,n29712 );
   nand U30916 ( n29712,n29668,n29449 );
   nand U30917 ( n29711,p3_instqueue_reg_12__2_,n29669 );
   nor U30918 ( n29709,n29450,n29670 );
   nor U30919 ( n29707,n29713,n29714 );
   nor U30920 ( n29714,n29453,n29673 );
   nor U30921 ( n29713,n29454,n29674 );
   nor U30922 ( n29716,n29717,n29718 );
   nand U30923 ( n29718,n29719,n29720 );
   nand U30924 ( n29720,n29668,n29461 );
   nand U30925 ( n29719,p3_instqueue_reg_12__1_,n29669 );
   nor U30926 ( n29717,n29462,n29670 );
   nor U30927 ( n29715,n29721,n29722 );
   nor U30928 ( n29722,n29465,n29673 );
   nor U30929 ( n29721,n29466,n29674 );
   nor U30930 ( n29724,n29725,n29726 );
   nand U30931 ( n29726,n29727,n29728 );
   nand U30932 ( n29728,n29668,n29473 );
   and U30933 ( n29668,n29729,n29483 );
   nand U30934 ( n29727,p3_instqueue_reg_12__0_,n29669 );
   nand U30935 ( n29669,n29730,n29731 );
   nand U30936 ( n29731,n29732,n29733 );
   nand U30937 ( n29733,n29479,n29734 );
   nand U30938 ( n29734,n29673,n29670 );
   nand U30939 ( n29732,n29735,n29483 );
   nor U30940 ( n29483,n29736,n29737 );
   nand U30941 ( n29730,n29484,n29738 );
   or U30942 ( n29738,n29674,n28350 );
   nor U30943 ( n29725,n29488,n29670 );
   nand U30944 ( n29670,n29739,n29489 );
   nor U30945 ( n29489,n29740,n29741 );
   nor U30946 ( n29723,n29742,n29743 );
   nor U30947 ( n29743,n29493,n29673 );
   nand U30948 ( n29673,n29744,n29495 );
   nor U30949 ( n29495,n29745,n29746 );
   nor U30950 ( n29742,n29496,n29674 );
   nand U30951 ( n29674,n29747,n29580 );
   nor U30952 ( n29580,n29278,n29235 );
   nor U30953 ( n29749,n29750,n29751 );
   nand U30954 ( n29751,n29752,n29753 );
   nand U30955 ( n29753,n29754,n29385 );
   nand U30956 ( n29752,p3_instqueue_reg_11__7_,n29755 );
   nor U30957 ( n29750,n29388,n29756 );
   nor U30958 ( n29748,n29757,n29758 );
   nor U30959 ( n29758,n29392,n29759 );
   nor U30960 ( n29757,n29394,n29760 );
   nor U30961 ( n29762,n29763,n29764 );
   nand U30962 ( n29764,n29765,n29766 );
   nand U30963 ( n29766,n29754,n29401 );
   nand U30964 ( n29765,p3_instqueue_reg_11__6_,n29755 );
   nor U30965 ( n29763,n29402,n29756 );
   nor U30966 ( n29761,n29767,n29768 );
   nor U30967 ( n29768,n29405,n29759 );
   nor U30968 ( n29767,n29406,n29760 );
   nor U30969 ( n29770,n29771,n29772 );
   nand U30970 ( n29772,n29773,n29774 );
   nand U30971 ( n29774,n29754,n29413 );
   nand U30972 ( n29773,p3_instqueue_reg_11__5_,n29755 );
   nor U30973 ( n29771,n29414,n29756 );
   nor U30974 ( n29769,n29775,n29776 );
   nor U30975 ( n29776,n29417,n29759 );
   nor U30976 ( n29775,n29418,n29760 );
   nor U30977 ( n29778,n29779,n29780 );
   nand U30978 ( n29780,n29781,n29782 );
   nand U30979 ( n29782,n29754,n29425 );
   nand U30980 ( n29781,p3_instqueue_reg_11__4_,n29755 );
   nor U30981 ( n29779,n29426,n29756 );
   nor U30982 ( n29777,n29783,n29784 );
   nor U30983 ( n29784,n29429,n29759 );
   nor U30984 ( n29783,n29430,n29760 );
   nor U30985 ( n29786,n29787,n29788 );
   nand U30986 ( n29788,n29789,n29790 );
   nand U30987 ( n29790,n29754,n29437 );
   nand U30988 ( n29789,p3_instqueue_reg_11__3_,n29755 );
   nor U30989 ( n29787,n29438,n29756 );
   nor U30990 ( n29785,n29791,n29792 );
   nor U30991 ( n29792,n29441,n29759 );
   nor U30992 ( n29791,n29442,n29760 );
   nor U30993 ( n29794,n29795,n29796 );
   nand U30994 ( n29796,n29797,n29798 );
   nand U30995 ( n29798,n29754,n29449 );
   nand U30996 ( n29797,p3_instqueue_reg_11__2_,n29755 );
   nor U30997 ( n29795,n29450,n29756 );
   nor U30998 ( n29793,n29799,n29800 );
   nor U30999 ( n29800,n29453,n29759 );
   nor U31000 ( n29799,n29454,n29760 );
   nor U31001 ( n29802,n29803,n29804 );
   nand U31002 ( n29804,n29805,n29806 );
   nand U31003 ( n29806,n29754,n29461 );
   nand U31004 ( n29805,p3_instqueue_reg_11__1_,n29755 );
   nor U31005 ( n29803,n29462,n29756 );
   nor U31006 ( n29801,n29807,n29808 );
   nor U31007 ( n29808,n29465,n29759 );
   nor U31008 ( n29807,n29466,n29760 );
   nor U31009 ( n29810,n29811,n29812 );
   nand U31010 ( n29812,n29813,n29814 );
   nand U31011 ( n29814,n29754,n29473 );
   and U31012 ( n29754,n29815,n29816 );
   nor U31013 ( n29815,n29474,n29817 );
   nand U31014 ( n29813,p3_instqueue_reg_11__0_,n29755 );
   nand U31015 ( n29755,n29818,n29819 );
   nand U31016 ( n29819,n29817,n29816 );
   nand U31017 ( n29816,n29479,n29820 );
   nand U31018 ( n29820,n29756,n29759 );
   and U31019 ( n29817,n29760,n29821 );
   nand U31020 ( n29821,n29822,n29482 );
   nand U31021 ( n29818,n29484,n29823 );
   or U31022 ( n29823,n29760,n28350 );
   nor U31023 ( n29811,n29488,n29756 );
   nand U31024 ( n29756,n29824,n29490 );
   nor U31025 ( n29809,n29825,n29826 );
   nor U31026 ( n29826,n29493,n29759 );
   nand U31027 ( n29759,n29827,n29494 );
   nor U31028 ( n29825,n29496,n29760 );
   nand U31029 ( n29760,n29828,n29829 );
   nor U31030 ( n29831,n29832,n29833 );
   nand U31031 ( n29833,n29834,n29835 );
   nand U31032 ( n29835,n29836,n29385 );
   nand U31033 ( n29834,p3_instqueue_reg_10__7_,n29837 );
   nor U31034 ( n29832,n29388,n29838 );
   nor U31035 ( n29830,n29839,n29840 );
   nor U31036 ( n29840,n29392,n29841 );
   nor U31037 ( n29839,n29394,n29842 );
   nor U31038 ( n29844,n29845,n29846 );
   nand U31039 ( n29846,n29847,n29848 );
   nand U31040 ( n29848,n29836,n29401 );
   nand U31041 ( n29847,p3_instqueue_reg_10__6_,n29837 );
   nor U31042 ( n29845,n29402,n29838 );
   nor U31043 ( n29843,n29849,n29850 );
   nor U31044 ( n29850,n29405,n29841 );
   nor U31045 ( n29849,n29406,n29842 );
   nor U31046 ( n29852,n29853,n29854 );
   nand U31047 ( n29854,n29855,n29856 );
   nand U31048 ( n29856,n29836,n29413 );
   nand U31049 ( n29855,p3_instqueue_reg_10__5_,n29837 );
   nor U31050 ( n29853,n29414,n29838 );
   nor U31051 ( n29851,n29857,n29858 );
   nor U31052 ( n29858,n29417,n29841 );
   nor U31053 ( n29857,n29418,n29842 );
   nor U31054 ( n29860,n29861,n29862 );
   nand U31055 ( n29862,n29863,n29864 );
   nand U31056 ( n29864,n29836,n29425 );
   nand U31057 ( n29863,p3_instqueue_reg_10__4_,n29837 );
   nor U31058 ( n29861,n29426,n29838 );
   nor U31059 ( n29859,n29865,n29866 );
   nor U31060 ( n29866,n29429,n29841 );
   nor U31061 ( n29865,n29430,n29842 );
   nor U31062 ( n29868,n29869,n29870 );
   nand U31063 ( n29870,n29871,n29872 );
   nand U31064 ( n29872,n29836,n29437 );
   nand U31065 ( n29871,p3_instqueue_reg_10__3_,n29837 );
   nor U31066 ( n29869,n29438,n29838 );
   nor U31067 ( n29867,n29873,n29874 );
   nor U31068 ( n29874,n29441,n29841 );
   nor U31069 ( n29873,n29442,n29842 );
   nor U31070 ( n29876,n29877,n29878 );
   nand U31071 ( n29878,n29879,n29880 );
   nand U31072 ( n29880,n29836,n29449 );
   nand U31073 ( n29879,p3_instqueue_reg_10__2_,n29837 );
   nor U31074 ( n29877,n29450,n29838 );
   nor U31075 ( n29875,n29881,n29882 );
   nor U31076 ( n29882,n29453,n29841 );
   nor U31077 ( n29881,n29454,n29842 );
   nor U31078 ( n29884,n29885,n29886 );
   nand U31079 ( n29886,n29887,n29888 );
   nand U31080 ( n29888,n29836,n29461 );
   nand U31081 ( n29887,p3_instqueue_reg_10__1_,n29837 );
   nor U31082 ( n29885,n29462,n29838 );
   nor U31083 ( n29883,n29889,n29890 );
   nor U31084 ( n29890,n29465,n29841 );
   nor U31085 ( n29889,n29466,n29842 );
   nor U31086 ( n29892,n29893,n29894 );
   nand U31087 ( n29894,n29895,n29896 );
   nand U31088 ( n29896,n29836,n29473 );
   and U31089 ( n29836,n29897,n29898 );
   nor U31090 ( n29897,n29474,n29899 );
   nand U31091 ( n29895,p3_instqueue_reg_10__0_,n29837 );
   nand U31092 ( n29837,n29900,n29901 );
   nand U31093 ( n29901,n29899,n29898 );
   nand U31094 ( n29898,n29479,n29902 );
   nand U31095 ( n29902,n29838,n29841 );
   and U31096 ( n29899,n29842,n29903 );
   nand U31097 ( n29903,n29822,n29572 );
   nand U31098 ( n29900,n29484,n29904 );
   or U31099 ( n29904,n29842,n28350 );
   nor U31100 ( n29893,n29488,n29838 );
   nand U31101 ( n29838,n29824,n29575 );
   nor U31102 ( n29891,n29905,n29906 );
   nor U31103 ( n29906,n29493,n29841 );
   nand U31104 ( n29841,n29827,n29578 );
   nor U31105 ( n29905,n29496,n29842 );
   nand U31106 ( n29842,n29828,n29579 );
   nor U31107 ( n29908,n29909,n29910 );
   nand U31108 ( n29910,n29911,n29912 );
   nand U31109 ( n29912,n29913,n29385 );
   nand U31110 ( n29911,p3_instqueue_reg_9__7_,n29914 );
   nor U31111 ( n29909,n29388,n29915 );
   nor U31112 ( n29907,n29916,n29917 );
   nor U31113 ( n29917,n29392,n29918 );
   nor U31114 ( n29916,n29394,n29919 );
   nor U31115 ( n29921,n29922,n29923 );
   nand U31116 ( n29923,n29924,n29925 );
   nand U31117 ( n29925,n29913,n29401 );
   nand U31118 ( n29924,p3_instqueue_reg_9__6_,n29914 );
   nor U31119 ( n29922,n29402,n29915 );
   nor U31120 ( n29920,n29926,n29927 );
   nor U31121 ( n29927,n29405,n29918 );
   nor U31122 ( n29926,n29406,n29919 );
   nor U31123 ( n29929,n29930,n29931 );
   nand U31124 ( n29931,n29932,n29933 );
   nand U31125 ( n29933,n29913,n29413 );
   nand U31126 ( n29932,p3_instqueue_reg_9__5_,n29914 );
   nor U31127 ( n29930,n29414,n29915 );
   nor U31128 ( n29928,n29934,n29935 );
   nor U31129 ( n29935,n29417,n29918 );
   nor U31130 ( n29934,n29418,n29919 );
   nor U31131 ( n29937,n29938,n29939 );
   nand U31132 ( n29939,n29940,n29941 );
   nand U31133 ( n29941,n29913,n29425 );
   nand U31134 ( n29940,p3_instqueue_reg_9__4_,n29914 );
   nor U31135 ( n29938,n29426,n29915 );
   nor U31136 ( n29936,n29942,n29943 );
   nor U31137 ( n29943,n29429,n29918 );
   nor U31138 ( n29942,n29430,n29919 );
   nor U31139 ( n29945,n29946,n29947 );
   nand U31140 ( n29947,n29948,n29949 );
   nand U31141 ( n29949,n29913,n29437 );
   nand U31142 ( n29948,p3_instqueue_reg_9__3_,n29914 );
   nor U31143 ( n29946,n29438,n29915 );
   nor U31144 ( n29944,n29950,n29951 );
   nor U31145 ( n29951,n29441,n29918 );
   nor U31146 ( n29950,n29442,n29919 );
   nor U31147 ( n29953,n29954,n29955 );
   nand U31148 ( n29955,n29956,n29957 );
   nand U31149 ( n29957,n29913,n29449 );
   nand U31150 ( n29956,p3_instqueue_reg_9__2_,n29914 );
   nor U31151 ( n29954,n29450,n29915 );
   nor U31152 ( n29952,n29958,n29959 );
   nor U31153 ( n29959,n29453,n29918 );
   nor U31154 ( n29958,n29454,n29919 );
   nor U31155 ( n29961,n29962,n29963 );
   nand U31156 ( n29963,n29964,n29965 );
   nand U31157 ( n29965,n29913,n29461 );
   nand U31158 ( n29964,p3_instqueue_reg_9__1_,n29914 );
   nor U31159 ( n29962,n29462,n29915 );
   nor U31160 ( n29960,n29966,n29967 );
   nor U31161 ( n29967,n29465,n29918 );
   nor U31162 ( n29966,n29466,n29919 );
   nor U31163 ( n29969,n29970,n29971 );
   nand U31164 ( n29971,n29972,n29973 );
   nand U31165 ( n29973,n29913,n29473 );
   and U31166 ( n29913,n29974,n29975 );
   nor U31167 ( n29974,n29474,n29976 );
   nand U31168 ( n29972,p3_instqueue_reg_9__0_,n29914 );
   nand U31169 ( n29914,n29977,n29978 );
   nand U31170 ( n29978,n29976,n29975 );
   nand U31171 ( n29975,n29479,n29979 );
   nand U31172 ( n29979,n29915,n29918 );
   and U31173 ( n29976,n29919,n29980 );
   nand U31174 ( n29980,n29822,n29655 );
   nand U31175 ( n29977,n29484,n29981 );
   or U31176 ( n29981,n29919,n28350 );
   nor U31177 ( n29970,n29488,n29915 );
   nand U31178 ( n29915,n29824,n29657 );
   nor U31179 ( n29968,n29982,n29983 );
   nor U31180 ( n29983,n29493,n29918 );
   nand U31181 ( n29918,n29827,n29660 );
   nor U31182 ( n29982,n29496,n29919 );
   nand U31183 ( n29919,n29828,n29661 );
   nor U31184 ( n29985,n29986,n29987 );
   nand U31185 ( n29987,n29988,n29989 );
   nand U31186 ( n29989,n29990,n29385 );
   nand U31187 ( n29988,p3_instqueue_reg_8__7_,n29991 );
   nor U31188 ( n29986,n28190,n29992 );
   nor U31189 ( n29984,n29993,n29994 );
   nor U31190 ( n29994,n29392,n29995 );
   nor U31191 ( n29993,n28191,n29996 );
   nor U31192 ( n29998,n29999,n30000 );
   nand U31193 ( n30000,n30001,n30002 );
   nand U31194 ( n30002,n29990,n29401 );
   nand U31195 ( n30001,p3_instqueue_reg_8__6_,n29991 );
   nor U31196 ( n29999,n28195,n29992 );
   nor U31197 ( n29997,n30003,n30004 );
   nor U31198 ( n30004,n29405,n29995 );
   nor U31199 ( n30003,n28196,n29996 );
   nor U31200 ( n30006,n30007,n30008 );
   nand U31201 ( n30008,n30009,n30010 );
   nand U31202 ( n30010,n29990,n29413 );
   nand U31203 ( n30009,p3_instqueue_reg_8__5_,n29991 );
   nor U31204 ( n30007,n28201,n29992 );
   nor U31205 ( n30005,n30011,n30012 );
   nor U31206 ( n30012,n29417,n29995 );
   nor U31207 ( n30011,n28202,n29996 );
   nor U31208 ( n30014,n30015,n30016 );
   nand U31209 ( n30016,n30017,n30018 );
   nand U31210 ( n30018,n29990,n29425 );
   nand U31211 ( n30017,p3_instqueue_reg_8__4_,n29991 );
   nor U31212 ( n30015,n28208,n29992 );
   nor U31213 ( n30013,n30019,n30020 );
   nor U31214 ( n30020,n29429,n29995 );
   nor U31215 ( n30019,n28209,n29996 );
   nor U31216 ( n30022,n30023,n30024 );
   nand U31217 ( n30024,n30025,n30026 );
   nand U31218 ( n30026,n29990,n29437 );
   nand U31219 ( n30025,p3_instqueue_reg_8__3_,n29991 );
   nor U31220 ( n30023,n28216,n29992 );
   nor U31221 ( n30021,n30027,n30028 );
   nor U31222 ( n30028,n29441,n29995 );
   nor U31223 ( n30027,n28217,n29996 );
   nor U31224 ( n30030,n30031,n30032 );
   nand U31225 ( n30032,n30033,n30034 );
   nand U31226 ( n30034,n29990,n29449 );
   nand U31227 ( n30033,p3_instqueue_reg_8__2_,n29991 );
   nor U31228 ( n30031,n28228,n29992 );
   nor U31229 ( n30029,n30035,n30036 );
   nor U31230 ( n30036,n29453,n29995 );
   nor U31231 ( n30035,n28229,n29996 );
   nor U31232 ( n30038,n30039,n30040 );
   nand U31233 ( n30040,n30041,n30042 );
   nand U31234 ( n30042,n29990,n29461 );
   nand U31235 ( n30041,p3_instqueue_reg_8__1_,n29991 );
   nor U31236 ( n30039,n28246,n29992 );
   nor U31237 ( n30037,n30043,n30044 );
   nor U31238 ( n30044,n29465,n29995 );
   nor U31239 ( n30043,n28247,n29996 );
   nor U31240 ( n30046,n30047,n30048 );
   nand U31241 ( n30048,n30049,n30050 );
   nand U31242 ( n30050,n29990,n29473 );
   and U31243 ( n29990,n29822,n29729 );
   nand U31244 ( n30049,p3_instqueue_reg_8__0_,n29991 );
   nand U31245 ( n29991,n30051,n30052 );
   nand U31246 ( n30052,n30053,n30054 );
   nand U31247 ( n30054,n29479,n30055 );
   nand U31248 ( n30055,n29995,n29992 );
   nand U31249 ( n30053,n29822,n29735 );
   nand U31250 ( n30051,n29484,n30056 );
   or U31251 ( n30056,n29996,n28350 );
   nor U31252 ( n30047,n28270,n29992 );
   nand U31253 ( n29992,n29824,n29739 );
   nor U31254 ( n30045,n30057,n30058 );
   nor U31255 ( n30058,n29493,n29995 );
   nand U31256 ( n29995,n29827,n29744 );
   not U31257 ( n29827,n30059 );
   nor U31258 ( n30057,n28271,n29996 );
   nand U31259 ( n29996,n29828,n29747 );
   nor U31260 ( n29828,n29235,p3_instqueuewr_addr_reg_2_ );
   nor U31261 ( n30061,n30062,n30063 );
   nand U31262 ( n30063,n30064,n30065 );
   nand U31263 ( n30065,n30066,n29385 );
   nand U31264 ( n30064,p3_instqueue_reg_7__7_,n30067 );
   nor U31265 ( n30062,n29392,n30068 );
   nor U31266 ( n30060,n30069,n30070 );
   nor U31267 ( n30070,n29388,n30071 );
   nor U31268 ( n30069,n29394,n30072 );
   nor U31269 ( n30074,n30075,n30076 );
   nand U31270 ( n30076,n30077,n30078 );
   nand U31271 ( n30078,n30066,n29401 );
   nand U31272 ( n30077,p3_instqueue_reg_7__6_,n30067 );
   nor U31273 ( n30075,n29405,n30068 );
   nor U31274 ( n30073,n30079,n30080 );
   nor U31275 ( n30080,n29402,n30071 );
   nor U31276 ( n30079,n29406,n30072 );
   nor U31277 ( n30082,n30083,n30084 );
   nand U31278 ( n30084,n30085,n30086 );
   nand U31279 ( n30086,n30066,n29413 );
   nand U31280 ( n30085,p3_instqueue_reg_7__5_,n30067 );
   nor U31281 ( n30083,n29417,n30068 );
   nor U31282 ( n30081,n30087,n30088 );
   nor U31283 ( n30088,n29414,n30071 );
   nor U31284 ( n30087,n29418,n30072 );
   nor U31285 ( n30090,n30091,n30092 );
   nand U31286 ( n30092,n30093,n30094 );
   nand U31287 ( n30094,n30066,n29425 );
   nand U31288 ( n30093,p3_instqueue_reg_7__4_,n30067 );
   nor U31289 ( n30091,n29429,n30068 );
   nor U31290 ( n30089,n30095,n30096 );
   nor U31291 ( n30096,n29426,n30071 );
   nor U31292 ( n30095,n29430,n30072 );
   nor U31293 ( n30098,n30099,n30100 );
   nand U31294 ( n30100,n30101,n30102 );
   nand U31295 ( n30102,n30066,n29437 );
   nand U31296 ( n30101,p3_instqueue_reg_7__3_,n30067 );
   nor U31297 ( n30099,n29441,n30068 );
   nor U31298 ( n30097,n30103,n30104 );
   nor U31299 ( n30104,n29438,n30071 );
   nor U31300 ( n30103,n29442,n30072 );
   nor U31301 ( n30106,n30107,n30108 );
   nand U31302 ( n30108,n30109,n30110 );
   nand U31303 ( n30110,n30066,n29449 );
   nand U31304 ( n30109,p3_instqueue_reg_7__2_,n30067 );
   nor U31305 ( n30107,n29453,n30068 );
   nor U31306 ( n30105,n30111,n30112 );
   nor U31307 ( n30112,n29450,n30071 );
   nor U31308 ( n30111,n29454,n30072 );
   nor U31309 ( n30114,n30115,n30116 );
   nand U31310 ( n30116,n30117,n30118 );
   nand U31311 ( n30118,n30066,n29461 );
   nand U31312 ( n30117,p3_instqueue_reg_7__1_,n30067 );
   nor U31313 ( n30115,n29465,n30068 );
   nor U31314 ( n30113,n30119,n30120 );
   nor U31315 ( n30120,n29462,n30071 );
   nor U31316 ( n30119,n29466,n30072 );
   nor U31317 ( n30122,n30123,n30124 );
   nand U31318 ( n30124,n30125,n30126 );
   nand U31319 ( n30126,n30066,n29473 );
   and U31320 ( n30066,n30127,n30128 );
   nand U31321 ( n30125,p3_instqueue_reg_7__0_,n30067 );
   nand U31322 ( n30067,n30129,n30130 );
   nand U31323 ( n30130,n29484,n30072 );
   nor U31324 ( n30129,n29574,n30131 );
   nor U31325 ( n30131,n30132,n30127 );
   or U31326 ( n30127,n30133,n30134 );
   nor U31327 ( n30132,n30135,n30136 );
   and U31328 ( n30135,n30071,n30068 );
   nor U31329 ( n30123,n29493,n30068 );
   nor U31330 ( n30121,n30137,n30138 );
   nor U31331 ( n30138,n29496,n30072 );
   nor U31332 ( n30137,n29488,n30071 );
   nor U31333 ( n30140,n30141,n30142 );
   nand U31334 ( n30142,n30143,n30144 );
   nand U31335 ( n30144,n30145,n29385 );
   nand U31336 ( n30143,p3_instqueue_reg_6__7_,n30146 );
   nor U31337 ( n30141,n29388,n30147 );
   nor U31338 ( n30139,n30148,n30149 );
   nor U31339 ( n30149,n29392,n30150 );
   nor U31340 ( n30148,n29394,n30151 );
   nor U31341 ( n30153,n30154,n30155 );
   nand U31342 ( n30155,n30156,n30157 );
   nand U31343 ( n30157,n30145,n29401 );
   nand U31344 ( n30156,p3_instqueue_reg_6__6_,n30146 );
   nor U31345 ( n30154,n29402,n30147 );
   nor U31346 ( n30152,n30158,n30159 );
   nor U31347 ( n30159,n29405,n30150 );
   nor U31348 ( n30158,n29406,n30151 );
   nor U31349 ( n30161,n30162,n30163 );
   nand U31350 ( n30163,n30164,n30165 );
   nand U31351 ( n30165,n30145,n29413 );
   nand U31352 ( n30164,p3_instqueue_reg_6__5_,n30146 );
   nor U31353 ( n30162,n29414,n30147 );
   nor U31354 ( n30160,n30166,n30167 );
   nor U31355 ( n30167,n29417,n30150 );
   nor U31356 ( n30166,n29418,n30151 );
   nor U31357 ( n30169,n30170,n30171 );
   nand U31358 ( n30171,n30172,n30173 );
   nand U31359 ( n30173,n30145,n29425 );
   nand U31360 ( n30172,p3_instqueue_reg_6__4_,n30146 );
   nor U31361 ( n30170,n29426,n30147 );
   nor U31362 ( n30168,n30174,n30175 );
   nor U31363 ( n30175,n29429,n30150 );
   nor U31364 ( n30174,n29430,n30151 );
   nor U31365 ( n30177,n30178,n30179 );
   nand U31366 ( n30179,n30180,n30181 );
   nand U31367 ( n30181,n30145,n29437 );
   nand U31368 ( n30180,p3_instqueue_reg_6__3_,n30146 );
   nor U31369 ( n30178,n29438,n30147 );
   nor U31370 ( n30176,n30182,n30183 );
   nor U31371 ( n30183,n29441,n30150 );
   nor U31372 ( n30182,n29442,n30151 );
   nor U31373 ( n30185,n30186,n30187 );
   nand U31374 ( n30187,n30188,n30189 );
   nand U31375 ( n30189,n30145,n29449 );
   nand U31376 ( n30188,p3_instqueue_reg_6__2_,n30146 );
   nor U31377 ( n30186,n29450,n30147 );
   nor U31378 ( n30184,n30190,n30191 );
   nor U31379 ( n30191,n29453,n30150 );
   nor U31380 ( n30190,n29454,n30151 );
   nor U31381 ( n30193,n30194,n30195 );
   nand U31382 ( n30195,n30196,n30197 );
   nand U31383 ( n30197,n30145,n29461 );
   nand U31384 ( n30196,p3_instqueue_reg_6__1_,n30146 );
   nor U31385 ( n30194,n29462,n30147 );
   nor U31386 ( n30192,n30198,n30199 );
   nor U31387 ( n30199,n29465,n30150 );
   nor U31388 ( n30198,n29466,n30151 );
   nor U31389 ( n30201,n30202,n30203 );
   nand U31390 ( n30203,n30204,n30205 );
   nand U31391 ( n30205,n30145,n29473 );
   and U31392 ( n30145,n30206,n30207 );
   nor U31393 ( n30206,n29474,n30208 );
   nand U31394 ( n30204,p3_instqueue_reg_6__0_,n30146 );
   nand U31395 ( n30146,n30209,n30210 );
   nand U31396 ( n30210,n30208,n30207 );
   nand U31397 ( n30207,n29479,n30211 );
   nand U31398 ( n30211,n30147,n30150 );
   and U31399 ( n30208,n30151,n30212 );
   nand U31400 ( n30212,n29572,n30213 );
   nand U31401 ( n30209,n29484,n30214 );
   or U31402 ( n30214,n30151,n28350 );
   nor U31403 ( n30202,n29488,n30147 );
   nand U31404 ( n30147,n29575,n30215 );
   nor U31405 ( n30200,n30216,n30217 );
   nor U31406 ( n30217,n29493,n30150 );
   nand U31407 ( n30150,n30218,n29578 );
   nor U31408 ( n30216,n29496,n30151 );
   nand U31409 ( n30151,n30219,n29579 );
   nor U31410 ( n30221,n30222,n30223 );
   nand U31411 ( n30223,n30224,n30225 );
   nand U31412 ( n30225,n30226,n29385 );
   nand U31413 ( n30224,p3_instqueue_reg_5__7_,n30227 );
   nor U31414 ( n30222,n28190,n30228 );
   nor U31415 ( n30220,n30229,n30230 );
   nor U31416 ( n30230,n27888,n30231 );
   nor U31417 ( n30229,n28191,n30232 );
   nor U31418 ( n30234,n30235,n30236 );
   nand U31419 ( n30236,n30237,n30238 );
   nand U31420 ( n30238,n30226,n29401 );
   nand U31421 ( n30237,p3_instqueue_reg_5__6_,n30227 );
   nor U31422 ( n30235,n28195,n30228 );
   nor U31423 ( n30233,n30239,n30240 );
   nor U31424 ( n30240,n27886,n30231 );
   nor U31425 ( n30239,n28196,n30232 );
   nor U31426 ( n30242,n30243,n30244 );
   nand U31427 ( n30244,n30245,n30246 );
   nand U31428 ( n30246,n30226,n29413 );
   nand U31429 ( n30245,p3_instqueue_reg_5__5_,n30227 );
   nor U31430 ( n30243,n28201,n30228 );
   nor U31431 ( n30241,n30247,n30248 );
   nor U31432 ( n30248,n27884,n30231 );
   nor U31433 ( n30247,n28202,n30232 );
   nor U31434 ( n30250,n30251,n30252 );
   nand U31435 ( n30252,n30253,n30254 );
   nand U31436 ( n30254,n30226,n29425 );
   nand U31437 ( n30253,p3_instqueue_reg_5__4_,n30227 );
   nor U31438 ( n30251,n28208,n30228 );
   nor U31439 ( n30249,n30255,n30256 );
   nor U31440 ( n30256,n27882,n30231 );
   nor U31441 ( n30255,n28209,n30232 );
   nor U31442 ( n30258,n30259,n30260 );
   nand U31443 ( n30260,n30261,n30262 );
   nand U31444 ( n30262,n30226,n29437 );
   nand U31445 ( n30261,p3_instqueue_reg_5__3_,n30227 );
   nor U31446 ( n30259,n28216,n30228 );
   nor U31447 ( n30257,n30263,n30264 );
   nor U31448 ( n30264,n27883,n30231 );
   nor U31449 ( n30263,n28217,n30232 );
   nor U31450 ( n30266,n30267,n30268 );
   nand U31451 ( n30268,n30269,n30270 );
   nand U31452 ( n30270,n30226,n29449 );
   nand U31453 ( n30269,p3_instqueue_reg_5__2_,n30227 );
   nor U31454 ( n30267,n28228,n30228 );
   nor U31455 ( n30265,n30271,n30272 );
   nor U31456 ( n30272,n27885,n30231 );
   nor U31457 ( n30271,n28229,n30232 );
   nor U31458 ( n30274,n30275,n30276 );
   nand U31459 ( n30276,n30277,n30278 );
   nand U31460 ( n30278,n30226,n29461 );
   nand U31461 ( n30277,p3_instqueue_reg_5__1_,n30227 );
   nor U31462 ( n30275,n28246,n30228 );
   nor U31463 ( n30273,n30279,n30280 );
   nor U31464 ( n30280,n27887,n30231 );
   nor U31465 ( n30279,n28247,n30232 );
   nor U31466 ( n30282,n30283,n30284 );
   nand U31467 ( n30284,n30285,n30286 );
   nand U31468 ( n30286,n30226,n29473 );
   and U31469 ( n30226,n30287,n30288 );
   nor U31470 ( n30287,n29474,n30289 );
   nand U31471 ( n30285,p3_instqueue_reg_5__0_,n30227 );
   nand U31472 ( n30227,n30290,n30291 );
   nand U31473 ( n30291,n30289,n30288 );
   nand U31474 ( n30288,n29479,n30292 );
   nand U31475 ( n30292,n30228,n30231 );
   and U31476 ( n30289,n30232,n30293 );
   nand U31477 ( n30293,n29655,n30213 );
   nand U31478 ( n30290,n29484,n30294 );
   or U31479 ( n30294,n30232,n28350 );
   nor U31480 ( n30283,n28270,n30228 );
   nand U31481 ( n30228,n29657,n30215 );
   nor U31482 ( n30281,n30295,n30296 );
   nor U31483 ( n30296,n27889,n30231 );
   nand U31484 ( n30231,n30218,n29660 );
   nor U31485 ( n30295,n28271,n30232 );
   nand U31486 ( n30232,n30219,n29661 );
   nor U31487 ( n30298,n30299,n30300 );
   nand U31488 ( n30300,n30301,n30302 );
   nand U31489 ( n30302,p3_instqueue_reg_4__7_,n30303 );
   nand U31490 ( n30301,n30304,n30305 );
   nor U31491 ( n30299,n30306,n30307 );
   nor U31492 ( n30297,n30308,n30309 );
   nor U31493 ( n30309,n28191,n30310 );
   nor U31494 ( n30308,n28190,n30311 );
   nor U31495 ( n30313,n30314,n30315 );
   nand U31496 ( n30315,n30316,n30317 );
   nand U31497 ( n30317,p3_instqueue_reg_4__6_,n30303 );
   nand U31498 ( n30316,n30304,n30318 );
   nor U31499 ( n30314,n30319,n30307 );
   nor U31500 ( n30312,n30320,n30321 );
   nor U31501 ( n30321,n28196,n30310 );
   nor U31502 ( n30320,n28195,n30311 );
   nor U31503 ( n30323,n30324,n30325 );
   nand U31504 ( n30325,n30326,n30327 );
   nand U31505 ( n30327,p3_instqueue_reg_4__5_,n30303 );
   nand U31506 ( n30326,n30304,n30328 );
   nor U31507 ( n30324,n30329,n30307 );
   nor U31508 ( n30322,n30330,n30331 );
   nor U31509 ( n30331,n28202,n30310 );
   nor U31510 ( n30330,n28201,n30311 );
   nor U31511 ( n30333,n30334,n30335 );
   nand U31512 ( n30335,n30336,n30337 );
   nand U31513 ( n30337,p3_instqueue_reg_4__4_,n30303 );
   nand U31514 ( n30336,n30304,n30338 );
   nor U31515 ( n30334,n30339,n30307 );
   nor U31516 ( n30332,n30340,n30341 );
   nor U31517 ( n30341,n28209,n30310 );
   nor U31518 ( n30340,n28208,n30311 );
   nor U31519 ( n30343,n30344,n30345 );
   nand U31520 ( n30345,n30346,n30347 );
   nand U31521 ( n30347,p3_instqueue_reg_4__3_,n30303 );
   nand U31522 ( n30346,n30304,n30348 );
   nor U31523 ( n30344,n30349,n30307 );
   nor U31524 ( n30342,n30350,n30351 );
   nor U31525 ( n30351,n28217,n30310 );
   nor U31526 ( n30350,n28216,n30311 );
   nor U31527 ( n30353,n30354,n30355 );
   nand U31528 ( n30355,n30356,n30357 );
   nand U31529 ( n30357,p3_instqueue_reg_4__2_,n30303 );
   nand U31530 ( n30356,n30304,n30358 );
   nor U31531 ( n30354,n30359,n30307 );
   nor U31532 ( n30352,n30360,n30361 );
   nor U31533 ( n30361,n28229,n30310 );
   nor U31534 ( n30360,n28228,n30311 );
   nor U31535 ( n30363,n30364,n30365 );
   nand U31536 ( n30365,n30366,n30367 );
   nand U31537 ( n30367,p3_instqueue_reg_4__1_,n30303 );
   nand U31538 ( n30366,n30304,n30368 );
   nor U31539 ( n30364,n30369,n30307 );
   nor U31540 ( n30362,n30370,n30371 );
   nor U31541 ( n30371,n28247,n30310 );
   nor U31542 ( n30370,n28246,n30311 );
   nor U31543 ( n30373,n30374,n30375 );
   nand U31544 ( n30375,n30376,n30377 );
   nand U31545 ( n30377,p3_instqueue_reg_4__0_,n30303 );
   nand U31546 ( n30303,n30378,n30379 );
   nand U31547 ( n30379,n30310,n29484 );
   nor U31548 ( n30378,n29574,n30380 );
   nor U31549 ( n30380,n30381,n30382 );
   nor U31550 ( n30382,n30383,n30384 );
   nor U31551 ( n30381,n30385,n30136 );
   nor U31552 ( n30385,n30304,n30386 );
   not U31553 ( n30386,n30311 );
   nand U31554 ( n30376,n30304,n30387 );
   and U31555 ( n30304,n30218,n29744 );
   nor U31556 ( n30374,n30388,n30307 );
   nand U31557 ( n30307,n29729,n30213 );
   nor U31558 ( n30372,n30389,n30390 );
   nor U31559 ( n30390,n28271,n30310 );
   nand U31560 ( n30310,n30219,n29747 );
   nor U31561 ( n30219,n29278,p3_instqueuewr_addr_reg_3_ );
   nor U31562 ( n30389,n28270,n30311 );
   nand U31563 ( n30311,n29739,n30215 );
   nor U31564 ( n30392,n30393,n30394 );
   nand U31565 ( n30394,n30395,n30396 );
   nand U31566 ( n30396,p3_instqueue_reg_3__7_,n30397 );
   nand U31567 ( n30395,n30398,n30305 );
   nor U31568 ( n30393,n30306,n30399 );
   nor U31569 ( n30391,n30400,n30401 );
   nor U31570 ( n30401,n28191,n30402 );
   nor U31571 ( n30400,n28190,n30403 );
   nor U31572 ( n30405,n30406,n30407 );
   nand U31573 ( n30407,n30408,n30409 );
   nand U31574 ( n30409,p3_instqueue_reg_3__6_,n30397 );
   nand U31575 ( n30408,n30398,n30318 );
   nor U31576 ( n30406,n30319,n30399 );
   nor U31577 ( n30404,n30410,n30411 );
   nor U31578 ( n30411,n28196,n30402 );
   nor U31579 ( n30410,n28195,n30403 );
   nor U31580 ( n30413,n30414,n30415 );
   nand U31581 ( n30415,n30416,n30417 );
   nand U31582 ( n30417,p3_instqueue_reg_3__5_,n30397 );
   nand U31583 ( n30416,n30398,n30328 );
   nor U31584 ( n30414,n30329,n30399 );
   nor U31585 ( n30412,n30418,n30419 );
   nor U31586 ( n30419,n28202,n30402 );
   nor U31587 ( n30418,n28201,n30403 );
   nor U31588 ( n30421,n30422,n30423 );
   nand U31589 ( n30423,n30424,n30425 );
   nand U31590 ( n30425,p3_instqueue_reg_3__4_,n30397 );
   nand U31591 ( n30424,n30398,n30338 );
   nor U31592 ( n30422,n30339,n30399 );
   nor U31593 ( n30420,n30426,n30427 );
   nor U31594 ( n30427,n28209,n30402 );
   nor U31595 ( n30426,n28208,n30403 );
   nor U31596 ( n30429,n30430,n30431 );
   nand U31597 ( n30431,n30432,n30433 );
   nand U31598 ( n30433,p3_instqueue_reg_3__3_,n30397 );
   nand U31599 ( n30432,n30398,n30348 );
   nor U31600 ( n30430,n30349,n30399 );
   nor U31601 ( n30428,n30434,n30435 );
   nor U31602 ( n30435,n28217,n30402 );
   nor U31603 ( n30434,n28216,n30403 );
   nor U31604 ( n30437,n30438,n30439 );
   nand U31605 ( n30439,n30440,n30441 );
   nand U31606 ( n30441,p3_instqueue_reg_3__2_,n30397 );
   nand U31607 ( n30440,n30398,n30358 );
   nor U31608 ( n30438,n30359,n30399 );
   nor U31609 ( n30436,n30442,n30443 );
   nor U31610 ( n30443,n28229,n30402 );
   nor U31611 ( n30442,n28228,n30403 );
   nor U31612 ( n30445,n30446,n30447 );
   nand U31613 ( n30447,n30448,n30449 );
   nand U31614 ( n30449,p3_instqueue_reg_3__1_,n30397 );
   nand U31615 ( n30448,n30398,n30368 );
   nor U31616 ( n30446,n30369,n30399 );
   nor U31617 ( n30444,n30450,n30451 );
   nor U31618 ( n30451,n28247,n30402 );
   nor U31619 ( n30450,n28246,n30403 );
   nor U31620 ( n30453,n30454,n30455 );
   nand U31621 ( n30455,n30456,n30457 );
   nand U31622 ( n30457,p3_instqueue_reg_3__0_,n30397 );
   nand U31623 ( n30397,n30458,n30459 );
   nand U31624 ( n30459,n30402,n29484 );
   nor U31625 ( n30458,n29574,n30460 );
   nor U31626 ( n30460,n30461,n30462 );
   nand U31627 ( n30462,n30463,n30402 );
   nand U31628 ( n30463,n29479,n30464 );
   nand U31629 ( n30464,n30403,n30465 );
   nor U31630 ( n30461,n30466,n30467 );
   nand U31631 ( n30456,n30398,n30387 );
   not U31632 ( n30398,n30465 );
   nand U31633 ( n30465,n30468,n29494 );
   nor U31634 ( n30454,n30388,n30399 );
   nand U31635 ( n30399,n30128,n30469 );
   nand U31636 ( n30469,n30470,n30402 );
   nand U31637 ( n30470,n30471,n29482 );
   nor U31638 ( n30452,n30472,n30473 );
   nor U31639 ( n30473,n28271,n30402 );
   nand U31640 ( n30402,n30474,n29829 );
   nor U31641 ( n30472,n28270,n30403 );
   nand U31642 ( n30403,n30475,n29490 );
   nor U31643 ( n30477,n30478,n30479 );
   nand U31644 ( n30479,n30480,n30481 );
   nand U31645 ( n30481,p3_instqueue_reg_2__7_,n30482 );
   nand U31646 ( n30480,n30483,n30305 );
   nor U31647 ( n30478,n30306,n30484 );
   nor U31648 ( n30476,n30485,n30486 );
   nor U31649 ( n30486,n28191,n30487 );
   nor U31650 ( n30485,n28190,n30488 );
   nor U31651 ( n30490,n30491,n30492 );
   nand U31652 ( n30492,n30493,n30494 );
   nand U31653 ( n30494,p3_instqueue_reg_2__6_,n30482 );
   nand U31654 ( n30493,n30483,n30318 );
   nor U31655 ( n30491,n30319,n30484 );
   nor U31656 ( n30489,n30495,n30496 );
   nor U31657 ( n30496,n28196,n30487 );
   nor U31658 ( n30495,n28195,n30488 );
   nor U31659 ( n30498,n30499,n30500 );
   nand U31660 ( n30500,n30501,n30502 );
   nand U31661 ( n30502,p3_instqueue_reg_2__5_,n30482 );
   nand U31662 ( n30501,n30483,n30328 );
   nor U31663 ( n30499,n30329,n30484 );
   nor U31664 ( n30497,n30503,n30504 );
   nor U31665 ( n30504,n28202,n30487 );
   nor U31666 ( n30503,n28201,n30488 );
   nor U31667 ( n30506,n30507,n30508 );
   nand U31668 ( n30508,n30509,n30510 );
   nand U31669 ( n30510,p3_instqueue_reg_2__4_,n30482 );
   nand U31670 ( n30509,n30483,n30338 );
   nor U31671 ( n30507,n30339,n30484 );
   nor U31672 ( n30505,n30511,n30512 );
   nor U31673 ( n30512,n28209,n30487 );
   nor U31674 ( n30511,n28208,n30488 );
   nor U31675 ( n30514,n30515,n30516 );
   nand U31676 ( n30516,n30517,n30518 );
   nand U31677 ( n30518,p3_instqueue_reg_2__3_,n30482 );
   nand U31678 ( n30517,n30483,n30348 );
   nor U31679 ( n30515,n30349,n30484 );
   nor U31680 ( n30513,n30519,n30520 );
   nor U31681 ( n30520,n28217,n30487 );
   nor U31682 ( n30519,n28216,n30488 );
   nor U31683 ( n30522,n30523,n30524 );
   nand U31684 ( n30524,n30525,n30526 );
   nand U31685 ( n30526,p3_instqueue_reg_2__2_,n30482 );
   nand U31686 ( n30525,n30483,n30358 );
   nor U31687 ( n30523,n30359,n30484 );
   nor U31688 ( n30521,n30527,n30528 );
   nor U31689 ( n30528,n28229,n30487 );
   nor U31690 ( n30527,n28228,n30488 );
   nor U31691 ( n30530,n30531,n30532 );
   nand U31692 ( n30532,n30533,n30534 );
   nand U31693 ( n30534,p3_instqueue_reg_2__1_,n30482 );
   nand U31694 ( n30533,n30483,n30368 );
   nor U31695 ( n30531,n30369,n30484 );
   nor U31696 ( n30529,n30535,n30536 );
   nor U31697 ( n30536,n28247,n30487 );
   nor U31698 ( n30535,n28246,n30488 );
   nor U31699 ( n30538,n30539,n30540 );
   nand U31700 ( n30540,n30541,n30542 );
   nand U31701 ( n30542,p3_instqueue_reg_2__0_,n30482 );
   nand U31702 ( n30482,n30543,n30544 );
   nand U31703 ( n30544,n30487,n29484 );
   nor U31704 ( n30543,n29574,n30545 );
   nor U31705 ( n30545,n30546,n30547 );
   nand U31706 ( n30547,n30548,n30487 );
   nand U31707 ( n30548,n29479,n30549 );
   nand U31708 ( n30549,n30488,n30550 );
   and U31709 ( n30546,n29572,n30471 );
   nand U31710 ( n30541,n30483,n30387 );
   not U31711 ( n30483,n30550 );
   nand U31712 ( n30550,n30468,n29578 );
   nor U31713 ( n30539,n30388,n30484 );
   nand U31714 ( n30484,n30128,n30551 );
   nand U31715 ( n30551,n30552,n30487 );
   nand U31716 ( n30552,n30471,n29572 );
   nor U31717 ( n30537,n30553,n30554 );
   nor U31718 ( n30554,n28271,n30487 );
   nand U31719 ( n30487,n30474,n29579 );
   nor U31720 ( n30553,n28270,n30488 );
   nand U31721 ( n30488,n30475,n29575 );
   nor U31722 ( n30556,n30557,n30558 );
   nand U31723 ( n30558,n30559,n30560 );
   nand U31724 ( n30560,p3_instqueue_reg_1__7_,n30561 );
   nand U31725 ( n30559,n30562,n30305 );
   nor U31726 ( n30557,n30306,n30563 );
   not U31727 ( n30306,n29385 );
   nor U31728 ( n30555,n30564,n30565 );
   nor U31729 ( n30565,n28191,n30566 );
   nor U31730 ( n30564,n28190,n30567 );
   nor U31731 ( n30569,n30570,n30571 );
   nand U31732 ( n30571,n30572,n30573 );
   nand U31733 ( n30573,p3_instqueue_reg_1__6_,n30561 );
   nand U31734 ( n30572,n30562,n30318 );
   nor U31735 ( n30570,n30319,n30563 );
   not U31736 ( n30319,n29401 );
   nor U31737 ( n30568,n30574,n30575 );
   nor U31738 ( n30575,n28196,n30566 );
   nor U31739 ( n30574,n28195,n30567 );
   nor U31740 ( n30577,n30578,n30579 );
   nand U31741 ( n30579,n30580,n30581 );
   nand U31742 ( n30581,p3_instqueue_reg_1__5_,n30561 );
   nand U31743 ( n30580,n30562,n30328 );
   nor U31744 ( n30578,n30329,n30563 );
   not U31745 ( n30329,n29413 );
   nor U31746 ( n30576,n30582,n30583 );
   nor U31747 ( n30583,n28202,n30566 );
   nor U31748 ( n30582,n28201,n30567 );
   nor U31749 ( n30585,n30586,n30587 );
   nand U31750 ( n30587,n30588,n30589 );
   nand U31751 ( n30589,p3_instqueue_reg_1__4_,n30561 );
   nand U31752 ( n30588,n30562,n30338 );
   nor U31753 ( n30586,n30339,n30563 );
   not U31754 ( n30339,n29425 );
   nor U31755 ( n30584,n30590,n30591 );
   nor U31756 ( n30591,n28209,n30566 );
   nor U31757 ( n30590,n28208,n30567 );
   nor U31758 ( n30593,n30594,n30595 );
   nand U31759 ( n30595,n30596,n30597 );
   nand U31760 ( n30597,p3_instqueue_reg_1__3_,n30561 );
   nand U31761 ( n30596,n30562,n30348 );
   nor U31762 ( n30594,n30349,n30563 );
   not U31763 ( n30349,n29437 );
   nor U31764 ( n30592,n30598,n30599 );
   nor U31765 ( n30599,n28217,n30566 );
   nor U31766 ( n30598,n28216,n30567 );
   nor U31767 ( n30601,n30602,n30603 );
   nand U31768 ( n30603,n30604,n30605 );
   nand U31769 ( n30605,p3_instqueue_reg_1__2_,n30561 );
   nand U31770 ( n30604,n30562,n30358 );
   nor U31771 ( n30602,n30359,n30563 );
   not U31772 ( n30359,n29449 );
   nor U31773 ( n30600,n30606,n30607 );
   nor U31774 ( n30607,n28229,n30566 );
   nor U31775 ( n30606,n28228,n30567 );
   nor U31776 ( n30609,n30610,n30611 );
   nand U31777 ( n30611,n30612,n30613 );
   nand U31778 ( n30613,p3_instqueue_reg_1__1_,n30561 );
   nand U31779 ( n30612,n30562,n30368 );
   nor U31780 ( n30610,n30369,n30563 );
   not U31781 ( n30369,n29461 );
   nor U31782 ( n30608,n30614,n30615 );
   nor U31783 ( n30615,n28247,n30566 );
   nor U31784 ( n30614,n28246,n30567 );
   nor U31785 ( n30617,n30618,n30619 );
   nand U31786 ( n30619,n30620,n30621 );
   nand U31787 ( n30621,p3_instqueue_reg_1__0_,n30561 );
   nand U31788 ( n30561,n30622,n30623 );
   nand U31789 ( n30623,n30566,n29484 );
   nor U31790 ( n30622,n29574,n30624 );
   nor U31791 ( n30624,n30625,n30626 );
   nand U31792 ( n30626,n30627,n30566 );
   nand U31793 ( n30627,n29479,n30628 );
   nand U31794 ( n30628,n30567,n30629 );
   not U31795 ( n29479,n30136 );
   and U31796 ( n30625,n29655,n30471 );
   nand U31797 ( n30620,n30562,n30387 );
   not U31798 ( n30562,n30629 );
   nand U31799 ( n30629,n30468,n29660 );
   nor U31800 ( n30618,n30388,n30563 );
   nand U31801 ( n30563,n30128,n30630 );
   nand U31802 ( n30630,n30631,n30566 );
   nand U31803 ( n30631,n30471,n29655 );
   not U31804 ( n30128,n29474 );
   nor U31805 ( n30616,n30632,n30633 );
   nor U31806 ( n30633,n28271,n30566 );
   nand U31807 ( n30566,n30474,n29661 );
   nor U31808 ( n30632,n28270,n30567 );
   nand U31809 ( n30567,n30475,n29657 );
   nor U31810 ( n30635,n30636,n30637 );
   nand U31811 ( n30637,n30638,n30639 );
   nand U31812 ( n30639,n30640,n30305 );
   not U31813 ( n30305,n29392 );
   nand U31814 ( n29392,n30641,buf2_reg_31_ );
   nand U31815 ( n30638,n30642,n29385 );
   nor U31816 ( n29385,n30643,n28350 );
   nor U31817 ( n30636,n29394,n30644 );
   nand U31818 ( n29394,n30645,n30646 );
   nor U31819 ( n30634,n30647,n30648 );
   nor U31820 ( n30648,n30649,n30650 );
   nor U31821 ( n30647,n29388,n30651 );
   nand U31822 ( n29388,n30641,buf2_reg_23_ );
   nor U31823 ( n30653,n30654,n30655 );
   nand U31824 ( n30655,n30656,n30657 );
   nand U31825 ( n30657,n30640,n30318 );
   not U31826 ( n30318,n29405 );
   nand U31827 ( n29405,n30641,buf2_reg_30_ );
   nand U31828 ( n30656,n30642,n29401 );
   nor U31829 ( n29401,n30658,n28350 );
   nor U31830 ( n30654,n29406,n30644 );
   nand U31831 ( n29406,n30645,n30659 );
   nor U31832 ( n30652,n30660,n30661 );
   nor U31833 ( n30661,n30649,n30662 );
   nor U31834 ( n30660,n29402,n30651 );
   nand U31835 ( n29402,n30641,buf2_reg_22_ );
   nor U31836 ( n30664,n30665,n30666 );
   nand U31837 ( n30666,n30667,n30668 );
   nand U31838 ( n30668,n30640,n30328 );
   not U31839 ( n30328,n29417 );
   nand U31840 ( n29417,n30641,buf2_reg_29_ );
   nand U31841 ( n30667,n30642,n29413 );
   nor U31842 ( n29413,n30669,n28350 );
   nor U31843 ( n30665,n29418,n30644 );
   nand U31844 ( n29418,n30645,n30670 );
   nor U31845 ( n30663,n30671,n30672 );
   nor U31846 ( n30672,n30649,n30673 );
   nor U31847 ( n30671,n29414,n30651 );
   nand U31848 ( n29414,n30641,buf2_reg_21_ );
   nor U31849 ( n30675,n30676,n30677 );
   nand U31850 ( n30677,n30678,n30679 );
   nand U31851 ( n30679,n30640,n30338 );
   not U31852 ( n30338,n29429 );
   nand U31853 ( n29429,n30641,buf2_reg_28_ );
   nand U31854 ( n30678,n30642,n29425 );
   nor U31855 ( n29425,n30680,n29574 );
   nor U31856 ( n30676,n29430,n30644 );
   nand U31857 ( n29430,n30645,n29309 );
   nor U31858 ( n30674,n30681,n30682 );
   nor U31859 ( n30682,n30649,n30683 );
   nor U31860 ( n30681,n29426,n30651 );
   nand U31861 ( n29426,n30641,buf2_reg_20_ );
   nor U31862 ( n30685,n30686,n30687 );
   nand U31863 ( n30687,n30688,n30689 );
   nand U31864 ( n30689,n30640,n30348 );
   not U31865 ( n30348,n29441 );
   nand U31866 ( n29441,n30641,buf2_reg_27_ );
   nand U31867 ( n30688,n30642,n29437 );
   nor U31868 ( n29437,n30690,n28350 );
   nor U31869 ( n30686,n29442,n30644 );
   nand U31870 ( n29442,n30645,n30691 );
   nor U31871 ( n30684,n30692,n30693 );
   nor U31872 ( n30693,n30649,n30694 );
   nor U31873 ( n30692,n29438,n30651 );
   nand U31874 ( n29438,n30641,buf2_reg_19_ );
   nor U31875 ( n30696,n30697,n30698 );
   nand U31876 ( n30698,n30699,n30700 );
   nand U31877 ( n30700,n30640,n30358 );
   not U31878 ( n30358,n29453 );
   nand U31879 ( n29453,n30641,buf2_reg_26_ );
   nand U31880 ( n30699,n30642,n29449 );
   nor U31881 ( n29449,n30701,n29574 );
   nor U31882 ( n30697,n29454,n30644 );
   nand U31883 ( n29454,n30645,n30702 );
   nor U31884 ( n30695,n30703,n30704 );
   nor U31885 ( n30704,n30649,n30705 );
   nor U31886 ( n30703,n29450,n30651 );
   nand U31887 ( n29450,n30641,buf2_reg_18_ );
   nor U31888 ( n30707,n30708,n30709 );
   nand U31889 ( n30709,n30710,n30711 );
   nand U31890 ( n30711,n30640,n30368 );
   not U31891 ( n30368,n29465 );
   nand U31892 ( n29465,n30641,buf2_reg_25_ );
   nand U31893 ( n30710,n30642,n29461 );
   nor U31894 ( n29461,n30712,n29574 );
   not U31895 ( n30642,n30713 );
   nor U31896 ( n30708,n29466,n30644 );
   nand U31897 ( n29466,n30645,n29366 );
   nor U31898 ( n30706,n30714,n30715 );
   nor U31899 ( n30715,n30649,n30716 );
   not U31900 ( n30649,n30717 );
   nor U31901 ( n30714,n29462,n30651 );
   nand U31902 ( n29462,n30641,buf2_reg_17_ );
   nor U31903 ( n30719,n30720,n30721 );
   nand U31904 ( n30721,n30722,n30723 );
   nand U31905 ( n30723,p3_instqueue_reg_0__0_,n30717 );
   nand U31906 ( n30717,n30724,n30725 );
   nand U31907 ( n30725,n30644,n29484 );
   nand U31908 ( n29484,n29487,n30726 );
   nor U31909 ( n30724,n29574,n30727 );
   nor U31910 ( n30727,n30728,n30729 );
   nor U31911 ( n30729,n30383,n30467 );
   not U31912 ( n30467,n30471 );
   nor U31913 ( n30728,n30730,n30136 );
   nor U31914 ( n30730,n30640,n30731 );
   not U31915 ( n30731,n30651 );
   nand U31916 ( n30722,n30640,n30387 );
   not U31917 ( n30387,n29493 );
   nand U31918 ( n29493,n30641,buf2_reg_24_ );
   and U31919 ( n30640,n30468,n29744 );
   and U31920 ( n29744,n30732,p3_instqueuewr_addr_reg_0_ );
   and U31921 ( n30468,n29746,n29745 );
   nor U31922 ( n30720,n30388,n30713 );
   nand U31923 ( n30713,n30471,n29729 );
   nor U31924 ( n29729,n30383,n29474 );
   nor U31925 ( n29474,n30136,n30733 );
   nand U31926 ( n30136,n30734,n28808 );
   nor U31927 ( n30471,n30735,n30736 );
   not U31928 ( n30388,n29473 );
   nor U31929 ( n29473,n30737,n29574 );
   nor U31930 ( n30718,n30738,n30739 );
   nor U31931 ( n30739,n29496,n30644 );
   nand U31932 ( n30644,n30474,n29747 );
   nor U31933 ( n29747,p3_instqueuewr_addr_reg_1_,p3_instqueuewr_addr_reg_0_ );
   nor U31934 ( n30474,p3_instqueuewr_addr_reg_3_,p3_instqueuewr_addr_reg_2_ );
   nand U31935 ( n29496,n30645,n29350 );
   nor U31936 ( n30645,n30726,n28350 );
   nor U31937 ( n30738,n29488,n30651 );
   nand U31938 ( n30651,n30475,n29739 );
   nor U31939 ( n29739,n30740,p3_instqueuewr_addr_reg_0_ );
   nor U31940 ( n30475,n30741,n30742 );
   nand U31941 ( n29488,n30641,buf2_reg_16_ );
   nor U31942 ( n30641,n30743,n28350 );
   not U31943 ( n29232,p3_instqueuewr_addr_reg_4_ );
   nand U31944 ( n30746,p3_instqueuewr_addr_reg_3_,n30747 );
   nand U31945 ( n30747,n30744,n30748 );
   nand U31946 ( n30748,p3_state2_reg_3_,n29497 );
   nand U31947 ( n30745,n30749,n30744 );
   nand U31948 ( n30749,n30750,n30751 );
   nand U31949 ( n30751,n30133,p3_state2_reg_3_ );
   nor U31950 ( n30750,n30752,n30753 );
   and U31951 ( n30753,n30741,n30754 );
   nor U31952 ( n30752,n30755,n30743 );
   nor U31953 ( n30755,n30756,n30757 );
   nand U31954 ( n30757,n30068,n30059 );
   nand U31955 ( n30059,n29745,n30758 );
   nand U31956 ( n30068,n30218,n29494 );
   nor U31957 ( n30218,n30758,n29745 );
   nor U31958 ( n30756,n29494,n29746 );
   not U31959 ( n29746,n30758 );
   nand U31960 ( n30758,n30759,n30760 );
   or U31961 ( n30760,n29741,n29490 );
   nor U31962 ( n30759,n29824,n30761 );
   not U31963 ( n30761,n30071 );
   nand U31964 ( n30071,n29490,n30215 );
   nor U31965 ( n30215,n30741,n29740 );
   nor U31966 ( n29824,n30742,n29741 );
   not U31967 ( n29741,n30741 );
   nand U31968 ( n30741,n30762,n30763 );
   nand U31969 ( n30763,n30735,n30466 );
   nor U31970 ( n30762,n30134,n29822 );
   nor U31971 ( n29822,n29737,n30736 );
   not U31972 ( n29737,n30735 );
   nor U31973 ( n30134,n30384,n30466 );
   not U31974 ( n30466,n29482 );
   not U31975 ( n30384,n30213 );
   nor U31976 ( n30213,n30735,n29736 );
   nand U31977 ( n30735,n30072,n30764 );
   nand U31978 ( n30764,p3_instqueuewr_addr_reg_3_,n29497 );
   not U31979 ( n30072,n30133 );
   nor U31980 ( n30133,n29497,p3_instqueuewr_addr_reg_3_ );
   nand U31981 ( n30766,p3_instqueuewr_addr_reg_2_,n30767 );
   nand U31982 ( n30767,n30744,n30768 );
   nand U31983 ( n30768,p3_state2_reg_3_,n29326 );
   nand U31984 ( n30765,n30769,n30744 );
   nand U31985 ( n30769,n30770,n30771 );
   nand U31986 ( n30771,n30742,n30754 );
   nor U31987 ( n30770,n30772,n30773 );
   nor U31988 ( n30773,n30774,n30743 );
   xor U31989 ( n30774,n29494,n29745 );
   xor U31990 ( n29745,n29740,n29490 );
   nor U31991 ( n29490,n30775,n30776 );
   not U31992 ( n29740,n30742 );
   xor U31993 ( n30742,n30736,n29482 );
   nor U31994 ( n29482,n29735,p3_instqueuewr_addr_reg_0_ );
   not U31995 ( n30736,n29736 );
   nand U31996 ( n29736,n29497,n30777 );
   nand U31997 ( n30777,n29326,n29278 );
   nand U31998 ( n29497,n29829,p3_instqueuewr_addr_reg_2_ );
   nor U31999 ( n29494,n30732,p3_instqueuewr_addr_reg_0_ );
   nor U32000 ( n30772,n29326,n30778 );
   nand U32001 ( n30778,p3_state2_reg_3_,n29278 );
   not U32002 ( n29326,n29829 );
   nor U32003 ( n29829,n30775,n29316 );
   nand U32004 ( n30780,n29579,p3_state2_reg_3_ );
   nor U32005 ( n30779,n30781,n30782 );
   nor U32006 ( n30782,n30783,n30784 );
   nor U32007 ( n30784,n30785,n30786 );
   nand U32008 ( n30786,n30787,n30788 );
   nand U32009 ( n30788,n30733,n30789 );
   or U32010 ( n30789,n29660,n29578 );
   nor U32011 ( n29578,n30775,n30732 );
   and U32012 ( n29660,n30732,n30775 );
   nor U32013 ( n30732,n29575,n29657 );
   nor U32014 ( n29657,n30740,n30775 );
   nor U32015 ( n29575,n30776,p3_instqueuewr_addr_reg_0_ );
   not U32016 ( n30733,n30743 );
   nand U32017 ( n30743,p3_statebs16_reg,n28795 );
   nand U32018 ( n30787,n30754,n30740 );
   not U32019 ( n30740,n30776 );
   nor U32020 ( n30776,n29572,n29655 );
   nor U32021 ( n29655,n30383,p3_instqueuewr_addr_reg_0_ );
   not U32022 ( n30383,n29735 );
   nor U32023 ( n29572,n30775,n29735 );
   nor U32024 ( n29735,n29661,n29579 );
   nor U32025 ( n29579,n29316,p3_instqueuewr_addr_reg_0_ );
   nand U32026 ( n30754,n28791,n30734 );
   nand U32027 ( n30734,n28795,n28806 );
   not U32028 ( n28791,n28866 );
   and U32029 ( n30785,p3_state2_reg_3_,n29661 );
   nor U32030 ( n29661,n30775,p3_instqueuewr_addr_reg_1_ );
   not U32031 ( n30783,n30744 );
   nor U32032 ( n30781,n29316,n30744 );
   nand U32033 ( n30791,n30792,n30744 );
   nand U32034 ( n30792,n30793,n30794 );
   nand U32035 ( n30794,n28793,n29171 );
   nand U32036 ( n30793,p3_state2_reg_3_,n30775 );
   nand U32037 ( n30790,p3_instqueuewr_addr_reg_0_,n30795 );
   nand U32038 ( n30795,n30796,n30744 );
   nand U32039 ( n30744,n30797,n30798 );
   or U32040 ( n30798,n29171,n29170 );
   nand U32041 ( n29171,n30799,n30800 );
   nand U32042 ( n30799,n29197,n30801 );
   nand U32043 ( n30801,n28883,n30802 );
   nor U32044 ( n30797,n29487,n28886 );
   nor U32045 ( n28886,n30800,n29170 );
   nand U32046 ( n29170,n28793,p3_state2_reg_0_ );
   not U32047 ( n30800,p3_flush_reg );
   not U32048 ( n29487,n29574 );
   nand U32049 ( n29574,n30803,n28790 );
   nand U32050 ( n30803,n30804,n30805 );
   nand U32051 ( n30805,p3_state2_reg_2_,n28856 );
   nor U32052 ( n30804,n28850,n29149 );
   nor U32053 ( n28850,n30726,p3_instqueuerd_addr_reg_4_ );
   nor U32054 ( n30807,n30808,n30809 );
   nor U32055 ( n30809,n30810,n28839 );
   nor U32056 ( n30810,n30811,n30812 );
   nor U32057 ( n30808,p3_instaddrpointer_reg_0_,n30813 );
   nor U32058 ( n30806,n30814,n30815 );
   nand U32059 ( n30815,n30816,n30817 );
   nand U32060 ( n30817,n30818,n30819 );
   nand U32061 ( n30816,n30820,n30821 );
   nor U32062 ( n30814,n28823,n30822 );
   nor U32063 ( n30824,n30825,n30826 );
   nor U32064 ( n30826,n30827,n30828 );
   nor U32065 ( n30825,n30829,n28337 );
   nor U32066 ( n30823,n30831,n30832 );
   nand U32067 ( n30832,n30833,n30834 );
   nand U32068 ( n30834,p3_instaddrpointer_reg_1_,n30835 );
   nand U32069 ( n30835,n30836,n30837 );
   nand U32070 ( n30837,n30838,n28839 );
   nand U32071 ( n30833,n30839,n30840 );
   nand U32072 ( n30839,n28351,n30842 );
   nand U32073 ( n30842,n30838,p3_instaddrpointer_reg_0_ );
   nor U32074 ( n30831,n29064,n28125 );
   nor U32075 ( n30844,n30845,n30846 );
   nand U32076 ( n30846,n30847,n30848 );
   nand U32077 ( n30848,n30849,n30821 );
   not U32078 ( n30821,n30827 );
   nor U32079 ( n30827,n28222,n30851 );
   nand U32080 ( n30847,n30852,n30853 );
   nand U32081 ( n30853,n30854,n30855 );
   nand U32082 ( n30855,n30856,n30857 );
   or U32083 ( n30856,n30858,n30859 );
   nor U32084 ( n30854,n30860,n30861 );
   nor U32085 ( n30861,p3_instaddrpointer_reg_2_,n30862 );
   nand U32086 ( n30862,n30863,p3_instaddrpointer_reg_0_ );
   nor U32087 ( n30863,n30864,n30840 );
   nor U32088 ( n30860,n30865,n30866 );
   nor U32089 ( n30865,n30867,n30868 );
   nor U32090 ( n30868,p3_instaddrpointer_reg_0_,n30864 );
   nor U32091 ( n30867,p3_instaddrpointer_reg_1_,n30869 );
   nor U32092 ( n30869,n30870,n30871 );
   nor U32093 ( n30845,n30872,n28337 );
   nor U32094 ( n30843,n30873,n30874 );
   nand U32095 ( n30874,n30875,n30876 );
   nand U32096 ( n30876,n30877,n30866 );
   nor U32097 ( n30877,n30840,n28351 );
   nand U32098 ( n30875,n30812,p3_instaddrpointer_reg_2_ );
   nor U32099 ( n30873,n29059,n30822 );
   nor U32100 ( n30879,n30880,n30881 );
   nand U32101 ( n30881,n30882,n30883 );
   or U32102 ( n30883,n30884,n30885 );
   nand U32103 ( n30882,n30850,n30886 );
   nor U32104 ( n30880,n30830,n30887 );
   nor U32105 ( n30878,n30888,n30889 );
   nand U32106 ( n30889,n30890,n30891 );
   nand U32107 ( n30891,p3_instaddrpointer_reg_3_,n30892 );
   nand U32108 ( n30892,n30893,n30894 );
   nand U32109 ( n30894,n30811,n30895 );
   nand U32110 ( n30890,n30896,n30897 );
   nand U32111 ( n30896,n30898,n30899 );
   or U32112 ( n30899,n30841,n30895 );
   nand U32113 ( n30898,n30852,n30900 );
   nor U32114 ( n30888,n29054,n28126 );
   nor U32115 ( n30902,n30903,n30904 );
   nand U32116 ( n30904,n30905,n30906 );
   nand U32117 ( n30906,n30907,n30850 );
   or U32118 ( n30905,n30908,n28240 );
   and U32119 ( n30903,n30909,n30818 );
   nor U32120 ( n30901,n30910,n30911 );
   nand U32121 ( n30911,n30912,n30913 );
   nand U32122 ( n30913,p3_instaddrpointer_reg_4_,n30914 );
   nand U32123 ( n30914,n30915,n30893 );
   and U32124 ( n30893,n30916,n30917 );
   nand U32125 ( n30917,n30918,n30858 );
   nor U32126 ( n30916,n30812,n30919 );
   nor U32127 ( n30919,n30859,n30920 );
   nor U32128 ( n30915,n30921,n30922 );
   nor U32129 ( n30922,n30923,n28351 );
   nor U32130 ( n30921,p3_instaddrpointer_reg_3_,n30813 );
   nand U32131 ( n30912,n30924,n30925 );
   nand U32132 ( n30924,n30926,n30927 );
   nand U32133 ( n30927,n30928,p3_instaddrpointer_reg_3_ );
   nor U32134 ( n30928,n30929,n28266 );
   nand U32135 ( n30926,n30923,n28235 );
   nor U32136 ( n30910,n29049,n28125 );
   nor U32137 ( n30932,n30933,n30934 );
   nand U32138 ( n30934,n30935,n30936 );
   nand U32139 ( n30936,n30851,n30937 );
   nand U32140 ( n30935,n30938,n30850 );
   nor U32141 ( n30933,n30830,n30939 );
   nor U32142 ( n30931,n30940,n30941 );
   nand U32143 ( n30941,n30942,n30943 );
   nand U32144 ( n30943,p3_instaddrpointer_reg_5_,n30944 );
   nand U32145 ( n30944,n30945,n30946 );
   nand U32146 ( n30946,n30811,n30947 );
   nand U32147 ( n30947,n30923,p3_instaddrpointer_reg_4_ );
   nand U32148 ( n30942,n30948,n30949 );
   nand U32149 ( n30948,n30950,n30951 );
   nand U32150 ( n30951,n30952,n30923 );
   nor U32151 ( n30952,n30841,n30925 );
   nand U32152 ( n30950,n30953,n30852 );
   nor U32153 ( n30940,n29044,n28126 );
   nor U32154 ( n30955,n30956,n30957 );
   nand U32155 ( n30957,n30958,n30959 );
   nand U32156 ( n30959,n30851,n30960 );
   nand U32157 ( n30958,n30850,n30961 );
   nor U32158 ( n30956,n30830,n30962 );
   nor U32159 ( n30954,n30963,n30964 );
   nand U32160 ( n30964,n30965,n30966 );
   nand U32161 ( n30966,p3_instaddrpointer_reg_6_,n30967 );
   nand U32162 ( n30967,n30968,n30945 );
   and U32163 ( n30945,n30969,n30836 );
   nand U32164 ( n30969,n30838,n30970 );
   nand U32165 ( n30970,n30971,n30972 );
   nor U32166 ( n30972,n30858,n30973 );
   nor U32167 ( n30973,n30864,n30859 );
   not U32168 ( n30858,n30974 );
   nor U32169 ( n30968,n30975,n30976 );
   nor U32170 ( n30976,n30977,n28351 );
   nor U32171 ( n30975,p3_instaddrpointer_reg_5_,n30813 );
   nand U32172 ( n30965,n30978,n30979 );
   nand U32173 ( n30978,n30980,n30981 );
   nand U32174 ( n30981,n30982,n30953 );
   and U32175 ( n30953,n30983,p3_instaddrpointer_reg_4_ );
   nor U32176 ( n30983,n30929,n30897 );
   not U32177 ( n30929,n30900 );
   nand U32178 ( n30900,n30984,n30985 );
   nand U32179 ( n30985,n30859,n30870 );
   nand U32180 ( n30984,n30974,n30857 );
   nor U32181 ( n30982,n30930,n30949 );
   nand U32182 ( n30980,n30977,n28235 );
   nor U32183 ( n30963,n29039,n30822 );
   nor U32184 ( n30987,n30988,n30989 );
   nand U32185 ( n30989,n30990,n30991 );
   or U32186 ( n30991,n30992,n28240 );
   nand U32187 ( n30990,n30850,n30993 );
   nor U32188 ( n30988,n28337,n30994 );
   nor U32189 ( n30986,n30995,n30996 );
   nand U32190 ( n30996,n30997,n30998 );
   nand U32191 ( n30998,p3_instaddrpointer_reg_7_,n30999 );
   nand U32192 ( n30999,n31000,n31001 );
   nand U32193 ( n31001,n30811,n31002 );
   nand U32194 ( n30997,n31003,n31004 );
   nand U32195 ( n31003,n31005,n31006 );
   or U32196 ( n31006,n31002,n28351 );
   nand U32197 ( n31005,n30852,n31007 );
   nor U32198 ( n30995,n29034,n28125 );
   nor U32199 ( n31009,n31010,n31011 );
   nand U32200 ( n31011,n31012,n31013 );
   nand U32201 ( n31013,n31014,n30851 );
   nand U32202 ( n31012,n30850,n31015 );
   nor U32203 ( n31010,n31016,n28337 );
   nor U32204 ( n31008,n31017,n31018 );
   nand U32205 ( n31018,n31019,n31020 );
   nand U32206 ( n31020,p3_instaddrpointer_reg_8_,n31021 );
   nand U32207 ( n31021,n31022,n31000 );
   and U32208 ( n31000,n31023,n31024 );
   nand U32209 ( n31024,n30918,n31025 );
   nor U32210 ( n31023,n30812,n31026 );
   nor U32211 ( n31026,n31027,n30920 );
   nor U32212 ( n31022,n31028,n31029 );
   nor U32213 ( n31029,n31030,n28351 );
   nor U32214 ( n31028,p3_instaddrpointer_reg_7_,n30813 );
   nand U32215 ( n31019,n31031,n31032 );
   nand U32216 ( n31031,n31033,n31034 );
   nand U32217 ( n31034,n31035,p3_instaddrpointer_reg_7_ );
   nand U32218 ( n31033,n31030,n28235 );
   nor U32219 ( n31017,n29029,n28126 );
   nor U32220 ( n31037,n31038,n31039 );
   nand U32221 ( n31039,n31040,n31041 );
   nand U32222 ( n31041,n31042,n30818 );
   nand U32223 ( n31040,n30851,n31043 );
   nor U32224 ( n31038,n31044,n31045 );
   nor U32225 ( n31036,n31046,n31047 );
   nand U32226 ( n31047,n31048,n31049 );
   nand U32227 ( n31049,n31050,n31051 );
   nand U32228 ( n31048,p3_instaddrpointer_reg_9_,n31052 );
   nand U32229 ( n31052,n31053,n31054 );
   or U32230 ( n31054,n30841,n31055 );
   nor U32231 ( n31046,n29024,n30822 );
   nor U32232 ( n31057,n31058,n31059 );
   nand U32233 ( n31059,n31060,n31061 );
   nand U32234 ( n31061,n31062,n30818 );
   nand U32235 ( n31060,n30851,n31063 );
   nor U32236 ( n31058,n31045,n31064 );
   nor U32237 ( n31056,n31065,n31066 );
   nand U32238 ( n31066,n31067,n31068 );
   nand U32239 ( n31068,p3_instaddrpointer_reg_10_,n31069 );
   nand U32240 ( n31069,n31070,n31053 );
   and U32241 ( n31053,n31071,n30836 );
   nand U32242 ( n31071,n30838,n31072 );
   nand U32243 ( n31072,n31073,n31074 );
   nor U32244 ( n31074,n31075,n31004 );
   nor U32245 ( n31075,n30864,n31027 );
   nor U32246 ( n31073,n31025,n31032 );
   nor U32247 ( n31070,n31076,n31077 );
   nor U32248 ( n31077,p3_instaddrpointer_reg_9_,n30813 );
   nand U32249 ( n31067,n31078,n31079 );
   and U32250 ( n31078,n31050,p3_instaddrpointer_reg_9_ );
   nand U32251 ( n31050,n31080,n31081 );
   nand U32252 ( n31081,n31082,n31035 );
   nor U32253 ( n31035,n31083,n28266 );
   not U32254 ( n31083,n31007 );
   nand U32255 ( n31007,n31084,n31085 );
   nand U32256 ( n31085,n31027,n30870 );
   not U32257 ( n31027,n31086 );
   or U32258 ( n31084,n31025,n31087 );
   nor U32259 ( n31082,n31004,n31032 );
   nand U32260 ( n31080,n31055,n28235 );
   nor U32261 ( n31065,n29019,n28125 );
   nor U32262 ( n31089,n31090,n31091 );
   nand U32263 ( n31091,n31092,n31093 );
   nand U32264 ( n31093,n30850,n31094 );
   nand U32265 ( n31092,n30818,n31095 );
   nor U32266 ( n31090,n31096,n28240 );
   nor U32267 ( n31088,n31097,n31098 );
   nand U32268 ( n31098,n31099,n31100 );
   nand U32269 ( n31100,p3_instaddrpointer_reg_11_,n31101 );
   nand U32270 ( n31101,n31102,n31103 );
   nor U32271 ( n31102,n31076,n31104 );
   nor U32272 ( n31104,p3_instaddrpointer_reg_10_,n28351 );
   and U32273 ( n31076,n30811,n31105 );
   nand U32274 ( n31105,n31055,p3_instaddrpointer_reg_9_ );
   nor U32275 ( n31055,n31106,n31032 );
   nand U32276 ( n31099,n31107,n31108 );
   nand U32277 ( n31107,n31109,n31110 );
   nand U32278 ( n31110,n31111,n31112 );
   nor U32279 ( n31111,n30841,n31106 );
   nand U32280 ( n31109,n30852,n31113 );
   nor U32281 ( n31097,n29014,n28126 );
   nor U32282 ( n31115,n31116,n31117 );
   nand U32283 ( n31117,n31118,n31119 );
   nand U32284 ( n31119,n31120,n30818 );
   nand U32285 ( n31118,n31121,n30850 );
   nor U32286 ( n31116,n30884,n31122 );
   nor U32287 ( n31114,n31123,n31124 );
   nand U32288 ( n31124,n31125,n31126 );
   nand U32289 ( n31126,p3_instaddrpointer_reg_12_,n31127 );
   nand U32290 ( n31127,n31128,n31103 );
   and U32291 ( n31103,n31129,n31130 );
   nand U32292 ( n31130,n30918,n31131 );
   nor U32293 ( n31129,n30812,n31132 );
   nor U32294 ( n31132,n31133,n30920 );
   not U32295 ( n30920,n31134 );
   nor U32296 ( n31128,n31135,n31136 );
   nor U32297 ( n31136,n31137,n28351 );
   nor U32298 ( n31135,p3_instaddrpointer_reg_11_,n30813 );
   nand U32299 ( n31125,n31138,n31139 );
   nand U32300 ( n31138,n31140,n31141 );
   nand U32301 ( n31141,n31142,p3_instaddrpointer_reg_11_ );
   nand U32302 ( n31140,n31137,n28235 );
   nor U32303 ( n31123,n29009,n28126 );
   nor U32304 ( n31144,n31145,n31146 );
   nand U32305 ( n31146,n31147,n31148 );
   nand U32306 ( n31148,n31149,n31150 );
   nand U32307 ( n31147,n31151,n31152 );
   nor U32308 ( n31145,n30884,n31153 );
   nor U32309 ( n31143,n31154,n31155 );
   nand U32310 ( n31155,n31156,n31157 );
   nand U32311 ( n31157,n31158,n31159 );
   nand U32312 ( n31156,p3_instaddrpointer_reg_13_,n31160 );
   nand U32313 ( n31160,n31161,n31162 );
   nand U32314 ( n31162,n30811,n31163 );
   not U32315 ( n31161,n31164 );
   nor U32316 ( n31154,n29004,n28125 );
   nor U32317 ( n31166,n31167,n31168 );
   nor U32318 ( n31168,p3_instaddrpointer_reg_14_,n31169 );
   nor U32319 ( n31169,n31170,n31171 );
   nand U32320 ( n31171,n31172,n31173 );
   nand U32321 ( n31173,p3_instaddrpointer_reg_13_,n31158 );
   nand U32322 ( n31158,n31174,n31175 );
   nand U32323 ( n31175,n31142,n31176 );
   nor U32324 ( n31142,n31177,n30930 );
   not U32325 ( n31177,n31113 );
   nand U32326 ( n31113,n31178,n31179 );
   nand U32327 ( n31179,n31133,n30870 );
   nand U32328 ( n31178,n31180,n30857 );
   nand U32329 ( n31174,n31181,n30811 );
   nand U32330 ( n31172,n31182,n30850 );
   nor U32331 ( n31170,n30830,n31183 );
   nor U32332 ( n31167,n31184,n31185 );
   nor U32333 ( n31184,n31164,n31186 );
   nand U32334 ( n31186,n31187,n31188 );
   nand U32335 ( n31187,n30838,n31159 );
   nand U32336 ( n31164,n31189,n31190 );
   nor U32337 ( n31190,n28221,n31191 );
   nor U32338 ( n31191,n31192,n30813 );
   nor U32339 ( n31192,n31193,n31194 );
   nand U32340 ( n31194,n31180,n31195 );
   nand U32341 ( n31195,n31196,n30870 );
   nor U32342 ( n31189,n31149,n31151 );
   nor U32343 ( n31151,n31197,n28337 );
   nor U32344 ( n31149,n31182,n31045 );
   nor U32345 ( n31165,n31198,n31199 );
   nor U32346 ( n31199,n28999,n30822 );
   and U32347 ( n31198,n31200,n30851 );
   nor U32348 ( n31202,n31203,n31204 );
   and U32349 ( n31204,n31205,n30851 );
   nor U32350 ( n31203,n31206,n31185 );
   nor U32351 ( n31206,n31207,n31208 );
   nand U32352 ( n31208,n31209,n31210 );
   nand U32353 ( n31210,n31211,n31212 );
   nor U32354 ( n31212,p3_instaddrpointer_reg_15_,n30841 );
   nand U32355 ( n31209,n31213,n31182 );
   nor U32356 ( n31207,n31183,n31214 );
   nand U32357 ( n31214,n30818,n31215 );
   nor U32358 ( n31201,n31216,n31217 );
   nand U32359 ( n31217,n31218,n31219 );
   nand U32360 ( n31219,p3_instaddrpointer_reg_15_,n31220 );
   nand U32361 ( n31220,n31221,n31222 );
   not U32362 ( n31222,n31223 );
   nor U32363 ( n31221,n31224,n31225 );
   nor U32364 ( n31225,p3_instaddrpointer_reg_14_,n28351 );
   not U32365 ( n31224,n31188 );
   nand U32366 ( n31188,n30811,n31226 );
   nand U32367 ( n31226,n31181,p3_instaddrpointer_reg_13_ );
   not U32368 ( n31181,n31163 );
   nand U32369 ( n31218,n31227,n31228 );
   nor U32370 ( n31216,n28994,n30822 );
   nor U32371 ( n31230,n31231,n31232 );
   nor U32372 ( n31232,p3_instaddrpointer_reg_16_,n31233 );
   nor U32373 ( n31233,n31234,n31235 );
   nand U32374 ( n31235,n31236,n31237 );
   nand U32375 ( n31237,n31238,n30850 );
   nand U32376 ( n31236,n31239,n30818 );
   nand U32377 ( n31234,n31240,n31241 );
   nand U32378 ( n31241,n31227,p3_instaddrpointer_reg_15_ );
   or U32379 ( n31240,n31242,n28351 );
   nor U32380 ( n31231,n31243,n31244 );
   nor U32381 ( n31243,n31223,n31245 );
   nand U32382 ( n31245,n31246,n31247 );
   nand U32383 ( n31247,n30838,n31228 );
   nand U32384 ( n31246,n30811,n31242 );
   nand U32385 ( n31223,n31248,n31249 );
   nor U32386 ( n31249,n31250,n31251 );
   nand U32387 ( n31251,n31252,n30836 );
   nand U32388 ( n31252,n31134,n31253 );
   nor U32389 ( n31250,n31254,n31255 );
   nor U32390 ( n31248,n31213,n31256 );
   nor U32391 ( n31256,n31239,n28337 );
   nor U32392 ( n31213,n31238,n31045 );
   nor U32393 ( n31229,n31257,n31258 );
   nor U32394 ( n31258,n28989,n28125 );
   and U32395 ( n31257,n31259,n30851 );
   nor U32396 ( n31261,n31262,n31263 );
   nand U32397 ( n31263,n31264,n31265 );
   nand U32398 ( n31265,n31266,n30818 );
   nand U32399 ( n31264,n31267,n30850 );
   nor U32400 ( n31262,n30884,n31268 );
   nor U32401 ( n31260,n31269,n31270 );
   nand U32402 ( n31270,n31271,n31272 );
   nand U32403 ( n31272,n31273,n31274 );
   nand U32404 ( n31271,p3_instaddrpointer_reg_17_,n31275 );
   nand U32405 ( n31275,n31276,n31277 );
   or U32406 ( n31277,n30841,n31278 );
   not U32407 ( n31276,n31279 );
   nor U32408 ( n31269,n28984,n28126 );
   nor U32409 ( n31281,n31282,n31283 );
   nor U32410 ( n31283,p3_instaddrpointer_reg_18_,n31284 );
   nor U32411 ( n31284,n31285,n31286 );
   nand U32412 ( n31286,n31287,n31288 );
   nand U32413 ( n31288,p3_instaddrpointer_reg_17_,n31273 );
   nand U32414 ( n31273,n31289,n31290 );
   nand U32415 ( n31290,n31227,n31291 );
   nor U32416 ( n31227,n31292,n30930 );
   and U32417 ( n31292,n31293,n31294 );
   nand U32418 ( n31294,n31295,n30870 );
   nand U32419 ( n31293,n31254,n30857 );
   nand U32420 ( n31289,n31278,n30811 );
   nor U32421 ( n31278,n31242,n31244 );
   nand U32422 ( n31287,n31296,n30850 );
   nor U32423 ( n31285,n30830,n31297 );
   nor U32424 ( n31282,n31298,n31299 );
   nor U32425 ( n31298,n31279,n31300 );
   nand U32426 ( n31300,n31301,n31302 );
   not U32427 ( n31302,n31303 );
   nand U32428 ( n31301,n30838,n31274 );
   nand U32429 ( n31279,n31304,n31305 );
   nor U32430 ( n31305,n30812,n31306 );
   nor U32431 ( n31306,n31307,n30930 );
   nor U32432 ( n31307,n31308,n31309 );
   nor U32433 ( n31309,n31310,n30864 );
   nor U32434 ( n31310,n31253,n31311 );
   nor U32435 ( n31308,n31312,n31087 );
   nor U32436 ( n31312,n31313,n31311 );
   not U32437 ( n31311,n31291 );
   nor U32438 ( n31291,n31244,n31228 );
   nor U32439 ( n31304,n31314,n31315 );
   nor U32440 ( n31315,n31316,n28337 );
   nor U32441 ( n31314,n31296,n31045 );
   nor U32442 ( n31280,n31317,n31318 );
   nor U32443 ( n31318,n28979,n28126 );
   and U32444 ( n31317,n30851,n31319 );
   nor U32445 ( n31321,n31322,n31323 );
   nor U32446 ( n31323,n30884,n31324 );
   nor U32447 ( n31322,n31325,n31299 );
   nor U32448 ( n31325,n31326,n31327 );
   nand U32449 ( n31327,n31328,n31329 );
   nand U32450 ( n31329,n31330,n31331 );
   nor U32451 ( n31330,p3_instaddrpointer_reg_19_,n28351 );
   nand U32452 ( n31328,n31332,n31296 );
   nor U32453 ( n31326,n31297,n31333 );
   nand U32454 ( n31333,n30818,n31334 );
   nor U32455 ( n31320,n31335,n31336 );
   nand U32456 ( n31336,n31337,n31338 );
   nand U32457 ( n31338,p3_instaddrpointer_reg_19_,n31339 );
   nand U32458 ( n31339,n31340,n31341 );
   not U32459 ( n31341,n31342 );
   nor U32460 ( n31340,n31303,n31343 );
   nor U32461 ( n31343,p3_instaddrpointer_reg_18_,n28351 );
   nor U32462 ( n31303,n30841,n31331 );
   nand U32463 ( n31337,n31344,n31345 );
   and U32464 ( n31344,n31346,n30852 );
   nor U32465 ( n31335,n28974,n28125 );
   nor U32466 ( n31348,n31349,n31350 );
   nor U32467 ( n31350,p3_instaddrpointer_reg_20_,n31351 );
   nor U32468 ( n31351,n31352,n31353 );
   nand U32469 ( n31353,n31354,n31355 );
   nand U32470 ( n31355,n30852,n31356 );
   nand U32471 ( n31356,n31357,n31358 );
   nand U32472 ( n31358,p3_instaddrpointer_reg_19_,n31346 );
   nand U32473 ( n31346,n31359,n31360 );
   or U32474 ( n31360,n31361,n30864 );
   nand U32475 ( n31359,n31362,n30857 );
   nand U32476 ( n31354,n31363,n30850 );
   nor U32477 ( n31352,n30830,n31334 );
   nor U32478 ( n31349,n31364,n31365 );
   nor U32479 ( n31364,n31342,n31366 );
   nand U32480 ( n31366,n31367,n31368 );
   not U32481 ( n31368,n31369 );
   nand U32482 ( n31367,n30838,n31345 );
   nand U32483 ( n31342,n31370,n31371 );
   nor U32484 ( n31371,n31372,n31373 );
   nand U32485 ( n31373,n31374,n30836 );
   nand U32486 ( n31374,n31134,n31361 );
   nor U32487 ( n31134,n30930,n30864 );
   nor U32488 ( n31372,n31362,n31255 );
   not U32489 ( n31255,n30918 );
   nor U32490 ( n30918,n30930,n31087 );
   not U32491 ( n31362,n31375 );
   nor U32492 ( n31370,n31332,n31376 );
   nor U32493 ( n31376,n31377,n28337 );
   nor U32494 ( n31332,n31363,n31045 );
   nor U32495 ( n31347,n31378,n31379 );
   nor U32496 ( n31379,n28969,n30822 );
   nor U32497 ( n31378,n30884,n31380 );
   nor U32498 ( n31382,n31383,n31384 );
   nand U32499 ( n31384,n31385,n31386 );
   nand U32500 ( n31386,n31387,n30818 );
   nand U32501 ( n31385,n31388,n30850 );
   and U32502 ( n31383,n31389,n30851 );
   nor U32503 ( n31381,n31390,n31391 );
   nand U32504 ( n31391,n31392,n31393 );
   nand U32505 ( n31393,p3_instaddrpointer_reg_21_,n31394 );
   nand U32506 ( n31394,n31395,n31396 );
   not U32507 ( n31396,n31397 );
   nor U32508 ( n31395,n31369,n31398 );
   nor U32509 ( n31398,p3_instaddrpointer_reg_20_,n28351 );
   nor U32510 ( n31369,n30841,n31399 );
   nand U32511 ( n31392,n31400,n31401 );
   nor U32512 ( n31400,n31402,n30930 );
   nor U32513 ( n31402,n31403,n31404 );
   nor U32514 ( n31403,n31365,n31357 );
   nand U32515 ( n31357,n31399,n30871 );
   nor U32516 ( n31390,n28964,n30822 );
   nor U32517 ( n31406,n31407,n31408 );
   nor U32518 ( n31408,n31409,n31410 );
   nor U32519 ( n31409,n31397,n31411 );
   nand U32520 ( n31411,n31412,n31413 );
   nand U32521 ( n31412,n30838,n31401 );
   nand U32522 ( n31397,n31414,n31415 );
   nand U32523 ( n31415,n30818,n31416 );
   nor U32524 ( n31414,n31417,n31418 );
   nor U32525 ( n31418,n31419,n31045 );
   nor U32526 ( n31417,n31420,n31421 );
   nor U32527 ( n31420,n31422,n31423 );
   nand U32528 ( n31423,n31424,n31425 );
   nand U32529 ( n31425,n31426,n31427 );
   nor U32530 ( n31424,n31428,n31429 );
   nor U32531 ( n31429,n31430,n31431 );
   nor U32532 ( n31428,n31432,n31433 );
   nand U32533 ( n31422,n31434,n31435 );
   nand U32534 ( n31435,n29208,n31436 );
   nor U32535 ( n31434,n30812,n31437 );
   nor U32536 ( n31437,n31432,n31438 );
   nor U32537 ( n31407,p3_instaddrpointer_reg_22_,n31439 );
   nor U32538 ( n31439,n31440,n31441 );
   nand U32539 ( n31441,n31442,n31443 );
   nand U32540 ( n31443,n30852,n31444 );
   nand U32541 ( n31444,n31445,n31446 );
   nand U32542 ( n31446,p3_instaddrpointer_reg_21_,n31404 );
   nand U32543 ( n31404,n31447,n31448 );
   nand U32544 ( n31448,n31432,n30870 );
   nand U32545 ( n31447,n31430,n30857 );
   nand U32546 ( n31442,n31419,n30850 );
   nor U32547 ( n31440,n30830,n31416 );
   nor U32548 ( n31405,n31449,n31450 );
   nor U32549 ( n31450,n28959,n28125 );
   and U32550 ( n31449,n30851,n31451 );
   nor U32551 ( n31453,n31454,n31455 );
   nand U32552 ( n31455,n31456,n31457 );
   nand U32553 ( n31457,n31458,n30818 );
   nand U32554 ( n31456,n31459,n30850 );
   and U32555 ( n31454,n31460,n30851 );
   nor U32556 ( n31452,n31461,n31462 );
   nand U32557 ( n31462,n31463,n31464 );
   nand U32558 ( n31464,p3_instaddrpointer_reg_23_,n31465 );
   nand U32559 ( n31465,n31466,n31467 );
   not U32560 ( n31467,n31468 );
   nor U32561 ( n31466,n31469,n31470 );
   nor U32562 ( n31470,p3_instaddrpointer_reg_22_,n28351 );
   not U32563 ( n31469,n31413 );
   nand U32564 ( n31413,n30811,n31471 );
   nand U32565 ( n31463,n31472,n31473 );
   nor U32566 ( n31472,n31474,n30930 );
   nor U32567 ( n31474,n31475,n31476 );
   nor U32568 ( n31475,n31410,n31445 );
   or U32569 ( n31445,n31471,n31477 );
   nor U32570 ( n31461,n28954,n28126 );
   nor U32571 ( n31479,n31480,n31481 );
   nor U32572 ( n31481,n31482,n31483 );
   nor U32573 ( n31482,n31468,n31484 );
   nand U32574 ( n31484,n31485,n31486 );
   not U32575 ( n31486,n31487 );
   nand U32576 ( n31485,n30838,n31473 );
   not U32577 ( n30838,n30813 );
   nand U32578 ( n31468,n31488,n31489 );
   nand U32579 ( n31489,n30818,n31490 );
   nor U32580 ( n31488,n31491,n31492 );
   nor U32581 ( n31492,n31493,n31045 );
   nor U32582 ( n31491,n31494,n31421 );
   nor U32583 ( n31494,n31495,n31496 );
   nand U32584 ( n31496,n31497,n31498 );
   nand U32585 ( n31498,n31499,n31427 );
   nor U32586 ( n31497,n31500,n31501 );
   nor U32587 ( n31501,n31502,n31431 );
   not U32588 ( n31431,n29221 );
   nor U32589 ( n31500,n31433,n31503 );
   nand U32590 ( n31495,n31504,n31505 );
   nand U32591 ( n31505,n29208,n31506 );
   nor U32592 ( n31504,n30812,n31507 );
   nor U32593 ( n31507,n31438,n31503 );
   not U32594 ( n31438,n31508 );
   nor U32595 ( n31480,p3_instaddrpointer_reg_24_,n31509 );
   nor U32596 ( n31509,n31510,n31511 );
   nand U32597 ( n31511,n31512,n31513 );
   nand U32598 ( n31513,n30852,n31514 );
   nand U32599 ( n31514,n31515,n31516 );
   nand U32600 ( n31516,p3_instaddrpointer_reg_23_,n31476 );
   nand U32601 ( n31476,n31517,n31518 );
   nand U32602 ( n31518,n31503,n30870 );
   not U32603 ( n31503,n31499 );
   nand U32604 ( n31517,n31502,n30857 );
   not U32605 ( n31502,n31506 );
   nand U32606 ( n31512,n31493,n30850 );
   nor U32607 ( n31510,n30830,n31490 );
   nor U32608 ( n31478,n31519,n31520 );
   nor U32609 ( n31520,n28949,n30822 );
   nor U32610 ( n31519,n31521,n28240 );
   nor U32611 ( n31523,n31524,n31525 );
   nand U32612 ( n31525,n31526,n31527 );
   nand U32613 ( n31527,n31528,n30818 );
   nand U32614 ( n31526,n31529,n30850 );
   nor U32615 ( n31524,n30884,n31530 );
   nor U32616 ( n31522,n31531,n31532 );
   nand U32617 ( n31532,n31533,n31534 );
   nand U32618 ( n31534,p3_instaddrpointer_reg_25_,n31535 );
   nand U32619 ( n31535,n31536,n31537 );
   nand U32620 ( n31537,n30811,n31483 );
   nor U32621 ( n31536,n31487,n31538 );
   nor U32622 ( n31487,n30841,n31539 );
   nand U32623 ( n31533,n31540,n31541 );
   nor U32624 ( n31540,n31542,n28266 );
   nor U32625 ( n31542,n31543,n31544 );
   nor U32626 ( n31543,n31483,n31515 );
   nand U32627 ( n31515,n31539,n30871 );
   nor U32628 ( n31531,n28944,n28125 );
   nor U32629 ( n31546,n31547,n31548 );
   nand U32630 ( n31548,n31549,n31550 );
   nand U32631 ( n31550,n31551,n31552 );
   nand U32632 ( n31549,n31553,n31554 );
   nor U32633 ( n31553,n31555,n28337 );
   nor U32634 ( n31547,n30884,n31556 );
   nor U32635 ( n31545,n31557,n31558 );
   nand U32636 ( n31558,n31559,n31560 );
   nand U32637 ( n31560,p3_instaddrpointer_reg_26_,n31561 );
   nand U32638 ( n31561,n31562,n31563 );
   not U32639 ( n31563,n31564 );
   nor U32640 ( n31562,n31538,n31565 );
   nor U32641 ( n31565,p3_instaddrpointer_reg_25_,n30813 );
   and U32642 ( n31538,n31566,n31567 );
   nand U32643 ( n31567,n31568,n31569 );
   nor U32644 ( n31569,n31570,n31571 );
   nand U32645 ( n31571,n31572,n30836 );
   nand U32646 ( n31572,n31573,n31508 );
   nor U32647 ( n31570,n31574,n29373 );
   nor U32648 ( n31568,n31575,n31576 );
   nand U32649 ( n31576,n31577,n31578 );
   nand U32650 ( n31578,n31573,n31579 );
   nand U32651 ( n31577,n29221,n31580 );
   nor U32652 ( n31575,n31581,n31582 );
   nand U32653 ( n31559,n31583,n31584 );
   nor U32654 ( n31583,n31585,n28266 );
   nor U32655 ( n31585,n31586,n31587 );
   and U32656 ( n31586,n31544,p3_instaddrpointer_reg_25_ );
   nand U32657 ( n31544,n31588,n31589 );
   nand U32658 ( n31589,n31582,n30870 );
   not U32659 ( n31582,n31573 );
   nand U32660 ( n31588,n31574,n30857 );
   not U32661 ( n31574,n31580 );
   nor U32662 ( n31557,n28939,n28126 );
   nor U32663 ( n31591,n31592,n31593 );
   nor U32664 ( n31593,n31594,n31595 );
   nor U32665 ( n31594,n31564,n31596 );
   nand U32666 ( n31596,n31597,n31598 );
   nand U32667 ( n31597,n30811,n31584 );
   nand U32668 ( n31564,n31599,n31600 );
   nand U32669 ( n31600,n30818,n31601 );
   nor U32670 ( n31599,n31602,n31551 );
   nor U32671 ( n31551,n31603,n31045 );
   and U32672 ( n31602,n31604,n30811 );
   nor U32673 ( n31592,p3_instaddrpointer_reg_27_,n31605 );
   nor U32674 ( n31605,n31606,n31607 );
   nand U32675 ( n31607,n31608,n31609 );
   nand U32676 ( n31609,n30852,n31610 );
   nand U32677 ( n31610,n31611,n31612 );
   nand U32678 ( n31612,n31587,p3_instaddrpointer_reg_26_ );
   nor U32679 ( n31587,n31604,n31477 );
   nand U32680 ( n31608,n31603,n30850 );
   nor U32681 ( n31606,n30830,n31601 );
   nor U32682 ( n31590,n31613,n31614 );
   nor U32683 ( n31614,n28934,n30822 );
   and U32684 ( n31613,n31615,n30851 );
   nor U32685 ( n31617,n31618,n31619 );
   nand U32686 ( n31619,n31620,n31621 );
   nand U32687 ( n31621,n31622,n30818 );
   nand U32688 ( n31620,n31623,n30850 );
   nor U32689 ( n31618,n28240,n31624 );
   nor U32690 ( n31616,n31625,n31626 );
   nand U32691 ( n31626,n31627,n31628 );
   nand U32692 ( n31628,p3_instaddrpointer_reg_28_,n31629 );
   nand U32693 ( n31629,n31630,n31631 );
   nand U32694 ( n31631,n31632,n30852 );
   nor U32695 ( n31630,n31633,n31634 );
   nor U32696 ( n31634,p3_instaddrpointer_reg_27_,n30813 );
   nand U32697 ( n30813,n30852,n31635 );
   nand U32698 ( n31635,n31087,n30864 );
   not U32699 ( n31633,n31598 );
   nand U32700 ( n31598,n31566,n31636 );
   nand U32701 ( n31636,n31637,n31638 );
   nor U32702 ( n31638,n31639,n31640 );
   nand U32703 ( n31640,n31641,n30836 );
   nand U32704 ( n31641,n31642,n31508 );
   nor U32705 ( n31639,n31643,n29373 );
   not U32706 ( n29373,n29208 );
   nor U32707 ( n31637,n31644,n31645 );
   nand U32708 ( n31645,n31646,n31647 );
   nand U32709 ( n31647,n31642,n31579 );
   not U32710 ( n31579,n31433 );
   nand U32711 ( n31646,n29221,n31648 );
   nor U32712 ( n31644,n31581,n31649 );
   not U32713 ( n31581,n31427 );
   nand U32714 ( n31627,n31650,n31651 );
   nor U32715 ( n31650,n31652,n28266 );
   nor U32716 ( n31652,n31653,n31654 );
   nor U32717 ( n31653,n31611,n31595 );
   and U32718 ( n31611,n31655,n31656 );
   nand U32719 ( n31656,n31649,n30870 );
   nand U32720 ( n31655,n31643,n30857 );
   nor U32721 ( n31625,n28929,n28125 );
   nor U32722 ( n31658,n31659,n31660 );
   nand U32723 ( n31660,n31661,n31662 );
   nand U32724 ( n31662,n31663,n31664 );
   nor U32725 ( n31663,n31665,n31045 );
   nand U32726 ( n31661,n31666,n31667 );
   nor U32727 ( n31666,n31668,n28337 );
   nor U32728 ( n31659,n30884,n31669 );
   nor U32729 ( n31657,n31670,n31671 );
   nand U32730 ( n31671,n31672,n31673 );
   nand U32731 ( n31673,p3_instaddrpointer_reg_29_,n31674 );
   nand U32732 ( n31674,n31675,n31676 );
   nor U32733 ( n31676,n30812,n31677 );
   nor U32734 ( n31677,n31678,n28266 );
   nor U32735 ( n31678,n31632,n31679 );
   and U32736 ( n31632,n31680,n30871 );
   not U32737 ( n30871,n31477 );
   nor U32738 ( n31675,n31681,n31682 );
   nor U32739 ( n31681,p3_instaddrpointer_reg_28_,n28351 );
   not U32740 ( n30841,n30811 );
   nor U32741 ( n30811,n30930,n31477 );
   nand U32742 ( n31672,n31683,n31684 );
   nor U32743 ( n31683,n31685,n30930 );
   nor U32744 ( n31685,n31686,n31687 );
   and U32745 ( n31686,p3_instaddrpointer_reg_28_,n31654 );
   nor U32746 ( n31654,n31680,n31477 );
   nor U32747 ( n31670,n28924,n30822 );
   nor U32748 ( n31689,n31690,n31691 );
   nor U32749 ( n31691,n28919,n28126 );
   and U32750 ( n31690,n31692,n30851 );
   not U32751 ( n30851,n30884 );
   nand U32752 ( n30884,n31693,n30852 );
   nor U32753 ( n31693,n31694,n31695 );
   nor U32754 ( n31688,n31696,n31697 );
   nand U32755 ( n31697,n31698,n31699 );
   nand U32756 ( n31699,n31700,n31701 );
   nand U32757 ( n31700,n31702,n31703 );
   nand U32758 ( n31703,n31668,n30818 );
   nor U32759 ( n31702,n31704,n31705 );
   nor U32760 ( n31705,n31045,n31706 );
   nor U32761 ( n31704,n31707,n30930 );
   nor U32762 ( n31707,n31708,n31709 );
   and U32763 ( n31709,n31687,p3_instaddrpointer_reg_29_ );
   nand U32764 ( n31687,n31710,n31711 );
   nand U32765 ( n31711,n31712,n30870 );
   nand U32766 ( n31710,n31713,n30857 );
   nor U32767 ( n31708,n31477,n31714 );
   nand U32768 ( n31698,p3_instaddrpointer_reg_30_,n31682 );
   nand U32769 ( n31682,n31715,n31716 );
   nand U32770 ( n31716,n30850,n31706 );
   not U32771 ( n30850,n31045 );
   nand U32772 ( n31045,n31717,n31694 );
   nor U32773 ( n31717,n31695,n28266 );
   not U32774 ( n30930,n30852 );
   nand U32775 ( n31715,n30818,n31718 );
   not U32776 ( n30818,n28337 );
   nand U32777 ( n30830,n30852,n29214 );
   nor U32778 ( n31696,n31701,n31719 );
   nand U32779 ( n31719,n31720,n31566 );
   not U32780 ( n31566,n31421 );
   nor U32781 ( n31421,n30812,n30852 );
   nand U32782 ( n31720,n31721,n31722 );
   nor U32783 ( n31722,n31723,n31724 );
   nand U32784 ( n31724,n31725,n30836 );
   nand U32785 ( n31725,n29222,n31714 );
   nor U32786 ( n31723,p3_instaddrpointer_reg_29_,n31726 );
   nor U32787 ( n31726,n30870,n30857 );
   nor U32788 ( n31721,n31679,n31727 );
   nand U32789 ( n31727,n31728,n31729 );
   nand U32790 ( n31729,n29210,n31714 );
   not U32791 ( n29210,n29352 );
   nand U32792 ( n31728,n31714,n31730 );
   nand U32793 ( n31730,n29223,n29351 );
   nor U32794 ( n29223,n31731,n28878 );
   nand U32795 ( n31679,n31732,n31733 );
   nand U32796 ( n31733,n31734,n30870 );
   nand U32797 ( n31732,n31735,n30857 );
   nor U32798 ( n31737,n30852,n31738 );
   nor U32799 ( n30852,n28808,n30812 );
   nor U32800 ( n31736,n31739,n31740 );
   nand U32801 ( n31740,n31741,n31742 );
   not U32802 ( n31742,n31738 );
   nand U32803 ( n31738,n31743,n31744 );
   or U32804 ( n31744,n28125,n28917 );
   nand U32805 ( n30822,n28808,n30836 );
   nand U32806 ( n31743,n30812,p3_instaddrpointer_reg_31_ );
   not U32807 ( n30812,n30836 );
   nand U32808 ( n30836,n31745,n31746 );
   nand U32809 ( n31746,n31747,n31748 );
   nand U32810 ( n31748,n31749,n31750 );
   nor U32811 ( n31750,n31751,n31752 );
   nor U32812 ( n31752,n30702,n31753 );
   nand U32813 ( n31753,n31754,n31755 );
   nand U32814 ( n31755,n31756,n29366 );
   nand U32815 ( n31756,n31757,n30659 );
   nand U32816 ( n31754,n29304,n31758 );
   nand U32817 ( n31758,n31759,n31760 );
   nor U32818 ( n31751,n31761,n29211 );
   nor U32819 ( n31761,n31762,n31763 );
   nor U32820 ( n31762,n30670,n31764 );
   nor U32821 ( n31749,n31765,n29376 );
   nand U32822 ( n29376,n31766,n31767 );
   nor U32823 ( n31767,n31768,n31769 );
   nor U32824 ( n31769,n29308,n31770 );
   nor U32825 ( n31770,n29350,n31771 );
   nor U32826 ( n31768,n31772,n30702 );
   nor U32827 ( n31772,n31773,n31774 );
   nand U32828 ( n31774,n31775,n31776 );
   nand U32829 ( n31776,n31777,n28771 );
   nor U32830 ( n31775,n31778,n31779 );
   nand U32831 ( n31773,n31780,n30646 );
   and U32832 ( n31780,n28810,n31781 );
   nor U32833 ( n31766,n31782,n31783 );
   nor U32834 ( n31783,n31784,n31777 );
   not U32835 ( n31782,n31785 );
   nor U32836 ( n31765,n31777,n29209 );
   nand U32837 ( n31745,n28775,n28790 );
   nor U32838 ( n31741,n31786,n31787 );
   nor U32839 ( n31787,n31477,n31788 );
   nor U32840 ( n31788,n31789,n31790 );
   nand U32841 ( n31790,n31791,n31792 );
   nand U32842 ( n31792,p3_instaddrpointer_reg_31_,n31714 );
   or U32843 ( n31791,n31793,n31714 );
   nand U32844 ( n31714,n31794,p3_instaddrpointer_reg_29_ );
   nor U32845 ( n31794,n31651,n31680 );
   nand U32846 ( n31680,n31795,p3_instaddrpointer_reg_27_ );
   nor U32847 ( n31795,n31584,n31604 );
   nand U32848 ( n31604,n31796,n31539 );
   nor U32849 ( n31539,n31797,n31471 );
   nand U32850 ( n31471,n31798,n31399 );
   and U32851 ( n31399,n31799,n31331 );
   nor U32852 ( n31331,n31800,n31242 );
   nand U32853 ( n31242,n31801,n31211 );
   nor U32854 ( n31211,n31159,n31163 );
   nand U32855 ( n31163,n31137,p3_instaddrpointer_reg_12_ );
   and U32856 ( n31137,n31802,p3_instaddrpointer_reg_11_ );
   nor U32857 ( n31802,n31106,n31803 );
   not U32858 ( n31106,n31030 );
   nor U32859 ( n31030,n31002,n31004 );
   nand U32860 ( n31002,n30977,p3_instaddrpointer_reg_6_ );
   and U32861 ( n30977,n31804,p3_instaddrpointer_reg_5_ );
   and U32862 ( n31804,p3_instaddrpointer_reg_4_,n30923 );
   nor U32863 ( n30923,n30897,n30895 );
   nor U32864 ( n31801,n31185,n31228 );
   nor U32865 ( n31477,n29271,n31805 );
   nand U32866 ( n31805,n29260,n29352 );
   nand U32867 ( n29271,n31806,n29351 );
   nand U32868 ( n29351,n31807,n29346 );
   not U32869 ( n29346,n31808 );
   nor U32870 ( n31807,n31809,n31810 );
   nor U32871 ( n31806,n31731,n29222 );
   nor U32872 ( n31786,n30864,n31811 );
   nor U32873 ( n31811,n31812,n31813 );
   nand U32874 ( n31813,n31814,n31815 );
   nand U32875 ( n31815,p3_instaddrpointer_reg_31_,n31734 );
   nand U32876 ( n31814,n31816,n31712 );
   not U32877 ( n31712,n31734 );
   nand U32878 ( n31734,n31817,n31649 );
   not U32879 ( n31649,n31642 );
   nand U32880 ( n31642,n31818,p3_instaddrpointer_reg_26_ );
   nor U32881 ( n31818,n31541,n31573 );
   nand U32882 ( n31573,n31819,p3_instaddrpointer_reg_24_ );
   nor U32883 ( n31819,n31473,n31499 );
   nand U32884 ( n31499,n31820,p3_instaddrpointer_reg_22_ );
   nor U32885 ( n31820,n31401,n31426 );
   not U32886 ( n31426,n31432 );
   nor U32887 ( n31432,n31821,n31361 );
   nand U32888 ( n31361,n31822,n31295 );
   not U32889 ( n31295,n31253 );
   nand U32890 ( n31253,n31823,n31133 );
   not U32891 ( n31133,n31196 );
   nand U32892 ( n31196,n31824,n31112 );
   nor U32893 ( n31824,n31004,n31086 );
   nand U32894 ( n31086,n31825,n30859 );
   nor U32895 ( n30859,n30895,n28839 );
   nand U32896 ( n30895,p3_instaddrpointer_reg_2_,p3_instaddrpointer_reg_1_ );
   not U32897 ( n30864,n30870 );
   nand U32898 ( n30870,n31826,n31433 );
   nor U32899 ( n31433,n29272,n29334 );
   nand U32900 ( n29272,n31827,n31828 );
   nor U32901 ( n31828,n31829,n31830 );
   nand U32902 ( n31830,n31831,n31781 );
   nand U32903 ( n31781,n31832,n31784 );
   nor U32904 ( n31832,n29304,n29309 );
   nand U32905 ( n31831,n31809,n31833 );
   nand U32906 ( n31833,n31834,n31777 );
   nor U32907 ( n31834,n31835,n31836 );
   nor U32908 ( n31836,n31837,n29366 );
   nor U32909 ( n31835,n29304,n30659 );
   nand U32910 ( n31829,n31838,n31839 );
   nand U32911 ( n31839,n31840,n30691 );
   and U32912 ( n31840,n31841,n31837 );
   nand U32913 ( n31838,n31842,n31778 );
   nor U32914 ( n31842,n28771,n31837 );
   nor U32915 ( n31827,n31843,n31844 );
   nand U32916 ( n31844,n31845,n31846 );
   nand U32917 ( n31846,n31847,n31848 );
   nand U32918 ( n31845,n31760,n29309 );
   nand U32919 ( n31843,n31849,n31850 );
   nand U32920 ( n31850,n29308,n31851 );
   nand U32921 ( n31851,n31852,n31853 );
   nor U32922 ( n31853,n31854,n31855 );
   nand U32923 ( n31855,n31856,n31785 );
   nand U32924 ( n31785,n31857,n31858 );
   nand U32925 ( n31858,n31859,n31860 );
   not U32926 ( n31860,n31779 );
   nand U32927 ( n31856,n31861,n29366 );
   nor U32928 ( n31861,n31862,n31863 );
   nor U32929 ( n31854,n29350,n31841 );
   nor U32930 ( n31852,n31864,n31865 );
   nor U32931 ( n31865,n31848,n31810 );
   nor U32932 ( n31864,n30691,n28804 );
   nand U32933 ( n31849,n31866,n30702 );
   nor U32934 ( n31866,n31867,n31868 );
   nor U32935 ( n31868,n30691,n31848 );
   nor U32936 ( n31867,n30646,n29302 );
   not U32937 ( n29302,n31869 );
   nor U32938 ( n31826,n31508,n31427 );
   nand U32939 ( n31427,n31870,n31871 );
   nor U32940 ( n31871,n31872,n31873 );
   nand U32941 ( n31873,n29363,n31874 );
   nand U32942 ( n29363,n31875,n31876 );
   nor U32943 ( n31876,n29308,n31877 );
   nor U32944 ( n31875,n28810,n30646 );
   not U32945 ( n28810,n31847 );
   nor U32946 ( n31872,n29306,n31878 );
   nand U32947 ( n31878,n31869,n29315 );
   nor U32948 ( n31870,n31879,n31880 );
   nor U32949 ( n31880,n29306,n31881 );
   nand U32950 ( n31881,n31869,n31857 );
   nand U32951 ( n29306,n31863,n31882 );
   nor U32952 ( n31882,n29308,n29309 );
   nor U32953 ( n31863,n30670,n30646 );
   nor U32954 ( n31879,n29362,n31883 );
   nand U32955 ( n31883,n31869,n31837 );
   nor U32956 ( n31869,n30659,n30691 );
   nand U32957 ( n31508,n31884,n31885 );
   nand U32958 ( n31885,n29335,n31778 );
   nor U32959 ( n29335,n29362,n31886 );
   nand U32960 ( n29362,n31887,n31888 );
   nor U32961 ( n31888,n31809,n31777 );
   nor U32962 ( n31887,n30702,n31810 );
   nand U32963 ( n31884,n29365,n31847 );
   nand U32964 ( n31739,n31889,n31890 );
   nand U32965 ( n31890,n31891,n30857 );
   not U32966 ( n30857,n31087 );
   nor U32967 ( n31087,n29221,n29208 );
   nand U32968 ( n31891,n31892,n31893 );
   not U32969 ( n31893,n31812 );
   nand U32970 ( n31812,n31894,n31895 );
   nand U32971 ( n31895,p3_instaddrpointer_reg_31_,n31684 );
   nor U32972 ( n31892,n31896,n31897 );
   and U32973 ( n31897,n31713,n31816 );
   nor U32974 ( n31816,n31793,n31684 );
   nor U32975 ( n31896,n31713,n31898 );
   not U32976 ( n31713,n31735 );
   nand U32977 ( n31735,n31817,n31643 );
   not U32978 ( n31643,n31648 );
   nand U32979 ( n31648,n31899,p3_instaddrpointer_reg_26_ );
   nor U32980 ( n31899,n31541,n31580 );
   nand U32981 ( n31580,n31900,p3_instaddrpointer_reg_24_ );
   nor U32982 ( n31900,n31473,n31506 );
   nand U32983 ( n31506,n31901,p3_instaddrpointer_reg_22_ );
   nor U32984 ( n31901,n31401,n31436 );
   not U32985 ( n31436,n31430 );
   nor U32986 ( n31430,n31821,n31375 );
   nand U32987 ( n31375,n31822,n31254 );
   not U32988 ( n31254,n31313 );
   nand U32989 ( n31313,n31823,n31180 );
   not U32990 ( n31180,n31131 );
   nand U32991 ( n31131,n31902,n31112 );
   not U32992 ( n31112,n31803 );
   nor U32993 ( n31902,n31004,n31025 );
   nand U32994 ( n31025,n31825,n30974 );
   nand U32995 ( n30974,n30866,n31903 );
   nand U32996 ( n31903,p3_instaddrpointer_reg_0_,p3_instaddrpointer_reg_1_ );
   and U32997 ( n31825,n31904,n30971 );
   nor U32998 ( n30971,n30897,n30925 );
   nor U32999 ( n31904,n30949,n30979 );
   and U33000 ( n31823,n31905,p3_instaddrpointer_reg_14_ );
   nor U33001 ( n31905,n31193,n31159 );
   and U33002 ( n31822,n31906,p3_instaddrpointer_reg_18_ );
   nor U33003 ( n31906,n31228,n31800 );
   not U33004 ( n31228,p3_instaddrpointer_reg_15_ );
   nor U33005 ( n31889,n31907,n31908 );
   and U33006 ( n31908,n31909,n29214 );
   nor U33007 ( n31907,n31695,n31910 );
   nand U33008 ( n31910,n31911,n31912 );
   nand U33009 ( n31912,n31913,n31694 );
   nand U33010 ( n31911,n31914,n31915 );
   nand U33011 ( n31914,n31916,n31917 );
   nor U33012 ( n31919,n31920,n31921 );
   nor U33013 ( n31921,n31922,n30819 );
   nor U33014 ( n31920,n30820,n31923 );
   not U33015 ( n30820,n30819 );
   nand U33016 ( n30819,n31924,n31925 );
   nand U33017 ( n31925,n31926,n28839 );
   nor U33018 ( n31918,n31927,n31928 );
   nor U33019 ( n31928,n28823,n31929 );
   nor U33020 ( n31927,n31930,n31931 );
   nor U33021 ( n31930,n31932,n31933 );
   nor U33022 ( n31935,n31936,n31937 );
   nor U33023 ( n31937,n30829,n31923 );
   xor U33024 ( n30829,n31938,n31939 );
   xor U33025 ( n31938,n31940,n30840 );
   nor U33026 ( n31936,n31922,n30828 );
   xor U33027 ( n30828,n31941,n31942 );
   xor U33028 ( n31941,n31924,n30840 );
   nor U33029 ( n31934,n31943,n31944 );
   nand U33030 ( n31944,n31945,n31946 );
   nand U33031 ( n31946,n31933,n31947 );
   nand U33032 ( n31945,p3_phyaddrpointer_reg_1_,n31932 );
   nor U33033 ( n31943,n29064,n31929 );
   nor U33034 ( n31949,n31950,n31951 );
   nand U33035 ( n31951,n31952,n31953 );
   nand U33036 ( n31953,n30849,n31954 );
   not U33037 ( n31954,n31922 );
   nor U33038 ( n31922,n31955,n31956 );
   xor U33039 ( n30849,n31957,n31958 );
   nand U33040 ( n31958,n31959,n31960 );
   or U33041 ( n31952,n31923,n30872 );
   xor U33042 ( n30872,n31961,n31962 );
   nand U33043 ( n31962,n31963,n31964 );
   nor U33044 ( n31950,n31965,n31966 );
   nor U33045 ( n31948,n31967,n31968 );
   nand U33046 ( n31968,n31969,n31970 );
   nand U33047 ( n31969,n31971,p3_phyaddrpointer_reg_2_ );
   nor U33048 ( n31967,n29059,n31929 );
   nor U33049 ( n31973,n31974,n31975 );
   nand U33050 ( n31975,n31976,n31977 );
   or U33051 ( n31977,n31923,n30887 );
   nand U33052 ( n30887,n31978,n31979 );
   nand U33053 ( n31979,n31980,n31981 );
   and U33054 ( n31981,n31982,n31964 );
   nor U33055 ( n31980,n31983,n31984 );
   nor U33056 ( n31984,n31985,n31961 );
   not U33057 ( n31985,n31963 );
   nand U33058 ( n31978,n31986,n31987 );
   nand U33059 ( n31987,n31988,n31982 );
   nand U33060 ( n31976,n31955,n30886 );
   and U33061 ( n30886,n31989,n31990 );
   nand U33062 ( n31990,n31991,n31992 );
   nand U33063 ( n31989,n31993,n31994 );
   nor U33064 ( n31974,n30885,n28263 );
   xor U33065 ( n30885,n31992,n31996 );
   nand U33066 ( n31996,n31960,n31997 );
   nand U33067 ( n31997,n31998,n31959 );
   not U33068 ( n31998,n31957 );
   nand U33069 ( n31992,n31994,n31999 );
   not U33070 ( n31994,n32000 );
   nor U33071 ( n31972,n32001,n32002 );
   nand U33072 ( n32002,n32003,n32004 );
   nand U33073 ( n32004,n32005,n31933 );
   nand U33074 ( n32003,n32006,p3_reip_reg_3_ );
   nand U33075 ( n32001,n32007,n32008 );
   nand U33076 ( n32008,p3_phyaddrpointer_reg_3_,n32009 );
   nand U33077 ( n32007,n32010,n32011 );
   nor U33078 ( n32010,n32012,n28133 );
   nor U33079 ( n32015,n32016,n32017 );
   nand U33080 ( n32017,n32018,n32019 );
   nand U33081 ( n32019,n30907,n28359 );
   nor U33082 ( n30907,n32020,n32021 );
   nor U33083 ( n32021,n32022,n32023 );
   and U33084 ( n32020,n32023,n32022 );
   nand U33085 ( n32018,n32024,n30909 );
   xor U33086 ( n30909,n32025,n32026 );
   nor U33087 ( n32025,n32027,n32028 );
   nor U33088 ( n32016,n30908,n28263 );
   xor U33089 ( n30908,n32029,n32022 );
   nand U33090 ( n32022,n32030,n32031 );
   nor U33091 ( n32014,n32032,n32033 );
   nand U33092 ( n32033,n32034,n32035 );
   nand U33093 ( n32035,n32036,n31933 );
   nand U33094 ( n32034,n32006,p3_reip_reg_4_ );
   nand U33095 ( n32032,n32037,n32038 );
   or U33096 ( n32038,n32039,n32040 );
   nand U33097 ( n32037,n32041,n32039 );
   and U33098 ( n32041,n32042,n32043 );
   nor U33099 ( n32045,n32046,n32047 );
   nand U33100 ( n32047,n32048,n32049 );
   nand U33101 ( n32049,n31955,n30938 );
   and U33102 ( n30938,n32050,n32051 );
   nand U33103 ( n32051,n32052,n32053 );
   nand U33104 ( n32050,n32054,n32055 );
   nand U33105 ( n32048,n31956,n30937 );
   nand U33106 ( n30937,n32056,n32057 );
   nand U33107 ( n32057,n32058,n32053 );
   nand U33108 ( n32053,n32059,n32060 );
   nand U33109 ( n32056,n32055,n32061 );
   xor U33110 ( n32055,p3_instaddrpointer_reg_5_,n32062 );
   nor U33111 ( n32046,n30939,n31923 );
   nand U33112 ( n30939,n32063,n32064 );
   nand U33113 ( n32064,n32065,n32066 );
   nor U33114 ( n32066,n32067,n32027 );
   not U33115 ( n32067,n32068 );
   nor U33116 ( n32065,n32069,n32070 );
   nor U33117 ( n32070,n32028,n32026 );
   not U33118 ( n32026,n32071 );
   not U33119 ( n32028,n32072 );
   not U33120 ( n32069,n32073 );
   nand U33121 ( n32063,n32074,n32075 );
   nand U33122 ( n32075,n32073,n32068 );
   nor U33123 ( n32044,n32076,n32077 );
   nand U33124 ( n32077,n32078,n32079 );
   nand U33125 ( n32079,n32080,n31933 );
   nand U33126 ( n32078,n28349,p3_reip_reg_5_ );
   nand U33127 ( n32076,n32081,n32082 );
   nand U33128 ( n32082,p3_phyaddrpointer_reg_5_,n32083 );
   nand U33129 ( n32081,n32084,n32085 );
   nor U33130 ( n32084,n28133,n32086 );
   nor U33131 ( n32088,n32089,n32090 );
   nand U33132 ( n32090,n32091,n32092 );
   nand U33133 ( n32092,n31956,n30960 );
   xor U33134 ( n30960,n32093,n32094 );
   nand U33135 ( n32091,n31955,n30961 );
   xor U33136 ( n30961,n32093,n32095 );
   nand U33137 ( n32093,n32096,n32097 );
   nor U33138 ( n32089,n30962,n31923 );
   xor U33139 ( n30962,n32098,n32099 );
   xor U33140 ( n32098,n32100,n30979 );
   nor U33141 ( n32087,n32101,n32102 );
   nand U33142 ( n32102,n32103,n32104 );
   nand U33143 ( n32104,n32105,n31933 );
   nand U33144 ( n32103,n32006,p3_reip_reg_6_ );
   nand U33145 ( n32101,n32106,n32107 );
   nand U33146 ( n32107,p3_phyaddrpointer_reg_6_,n32108 );
   nand U33147 ( n32108,n32109,n32110 );
   nand U33148 ( n32110,n32042,n32085 );
   not U33149 ( n32109,n32083 );
   nand U33150 ( n32083,n32040,n32111 );
   nand U33151 ( n32111,n32042,n32039 );
   nor U33152 ( n32040,n32009,n32112 );
   nor U33153 ( n32112,n32013,p3_phyaddrpointer_reg_3_ );
   nand U33154 ( n32009,n32113,n31970 );
   nand U33155 ( n31970,n32042,n32012 );
   nand U33156 ( n32106,n32114,n32115 );
   nor U33157 ( n32114,n32085,n32116 );
   or U33158 ( n32116,n32086,n28133 );
   nor U33159 ( n32118,n32119,n32120 );
   nand U33160 ( n32120,n32121,n32122 );
   nand U33161 ( n32122,n31955,n30993 );
   xor U33162 ( n30993,n32123,n32124 );
   xor U33163 ( n32123,p3_instaddrpointer_reg_7_,n32125 );
   or U33164 ( n32121,n31923,n30994 );
   xor U33165 ( n30994,n32126,n32127 );
   xor U33166 ( n32126,n32128,n31004 );
   nor U33167 ( n32119,n30992,n28263 );
   xor U33168 ( n30992,n32129,n32130 );
   xor U33169 ( n32129,n28175,p3_instaddrpointer_reg_7_ );
   nor U33170 ( n32117,n32132,n32133 );
   nand U33171 ( n32133,n32134,n32135 );
   nand U33172 ( n32135,n32136,n31933 );
   nand U33173 ( n32134,n28349,p3_reip_reg_7_ );
   nand U33174 ( n32132,n32137,n32138 );
   nand U33175 ( n32138,p3_phyaddrpointer_reg_7_,n32139 );
   nand U33176 ( n32137,n32140,n32141 );
   nor U33177 ( n32140,n32013,n32142 );
   nor U33178 ( n32144,n32145,n32146 );
   nand U33179 ( n32146,n32147,n32148 );
   nand U33180 ( n32148,n31956,n31014 );
   xor U33181 ( n31014,n32149,n32150 );
   nand U33182 ( n32147,n31955,n31015 );
   xor U33183 ( n31015,n32150,n32151 );
   xor U33184 ( n32150,n31032,n28169 );
   nor U33185 ( n32145,n31016,n31923 );
   not U33186 ( n31016,n32153 );
   xor U33187 ( n32153,n32154,n32155 );
   xor U33188 ( n32155,p3_instaddrpointer_reg_8_,n32156 );
   nor U33189 ( n32143,n32157,n32158 );
   nand U33190 ( n32158,n32159,n32160 );
   nand U33191 ( n32160,n32161,n31933 );
   nand U33192 ( n32159,n28349,p3_reip_reg_8_ );
   nand U33193 ( n32157,n32162,n32163 );
   nand U33194 ( n32163,n32164,n32165 );
   or U33195 ( n32162,n32165,n32166 );
   nor U33196 ( n32168,n32169,n32170 );
   nand U33197 ( n32170,n32171,n32172 );
   nand U33198 ( n32172,n32024,n31042 );
   xor U33199 ( n31042,p3_instaddrpointer_reg_9_,n32173 );
   nand U33200 ( n32171,n31956,n31043 );
   xor U33201 ( n31043,n32174,n32175 );
   or U33202 ( n32174,n32176,n32177 );
   nor U33203 ( n32169,n31044,n32178 );
   xor U33204 ( n31044,p3_instaddrpointer_reg_9_,n32179 );
   nand U33205 ( n32179,n32151,p3_instaddrpointer_reg_8_ );
   not U33206 ( n32151,n32180 );
   nor U33207 ( n32167,n32181,n32182 );
   nand U33208 ( n32182,n32183,n32184 );
   nand U33209 ( n32184,n32185,n31933 );
   nand U33210 ( n32183,n28349,p3_reip_reg_9_ );
   nand U33211 ( n32181,n32186,n32187 );
   nand U33212 ( n32187,p3_phyaddrpointer_reg_9_,n32188 );
   nand U33213 ( n32186,n32189,n32190 );
   nor U33214 ( n32189,n32165,n32191 );
   nor U33215 ( n32193,n32194,n32195 );
   nand U33216 ( n32195,n32196,n32197 );
   nand U33217 ( n32197,n31062,n28356 );
   nor U33218 ( n31062,n32198,n32199 );
   and U33219 ( n32199,n31079,n32200 );
   nand U33220 ( n32200,p3_instaddrpointer_reg_9_,n32173 );
   nand U33221 ( n32196,n31956,n31063 );
   xor U33222 ( n31063,n32152,n32201 );
   xor U33223 ( n32201,p3_instaddrpointer_reg_10_,n32202 );
   or U33224 ( n32202,n32203,n32176 );
   nor U33225 ( n32194,n31064,n32178 );
   nand U33226 ( n31064,n32204,n32205 );
   nand U33227 ( n32204,n31079,n32206 );
   nand U33228 ( n32206,n32207,p3_instaddrpointer_reg_9_ );
   nor U33229 ( n32207,n31032,n32180 );
   nor U33230 ( n32192,n32208,n32209 );
   nand U33231 ( n32209,n32210,n32211 );
   nand U33232 ( n32211,n32212,n31933 );
   nand U33233 ( n32210,n32006,p3_reip_reg_10_ );
   nand U33234 ( n32208,n32213,n32214 );
   nand U33235 ( n32214,p3_phyaddrpointer_reg_10_,n32215 );
   nand U33236 ( n32215,n32216,n32217 );
   nand U33237 ( n32217,n32042,n32190 );
   not U33238 ( n32216,n32188 );
   nand U33239 ( n32188,n32166,n32218 );
   nand U33240 ( n32218,n32042,n32165 );
   nor U33241 ( n32166,n32139,n32219 );
   nor U33242 ( n32219,n28134,p3_phyaddrpointer_reg_7_ );
   nand U33243 ( n32139,n32113,n32220 );
   nand U33244 ( n32220,n32042,n32142 );
   nand U33245 ( n32213,n32221,n32222 );
   nor U33246 ( n32221,n32190,n32223 );
   nand U33247 ( n32223,n32164,p3_phyaddrpointer_reg_8_ );
   not U33248 ( n32164,n32191 );
   nand U33249 ( n32191,n32224,n32225 );
   nor U33250 ( n32224,n28134,n32141 );
   nor U33251 ( n32227,n32228,n32229 );
   nand U33252 ( n32229,n32230,n32231 );
   nand U33253 ( n32231,n28359,n31094 );
   xor U33254 ( n31094,n31108,n32205 );
   nand U33255 ( n32230,n32024,n31095 );
   xor U33256 ( n31095,p3_instaddrpointer_reg_11_,n32198 );
   nor U33257 ( n32228,n31096,n28263 );
   xor U33258 ( n31096,n32232,n32233 );
   nand U33259 ( n32233,n32234,n32235 );
   nand U33260 ( n32235,n32203,n32236 );
   nand U33261 ( n32236,n28177,n31079 );
   xor U33262 ( n32232,n28177,p3_instaddrpointer_reg_11_ );
   nor U33263 ( n32226,n32237,n32238 );
   nand U33264 ( n32238,n32239,n32240 );
   nand U33265 ( n32240,n32241,n31933 );
   nand U33266 ( n32239,n32006,p3_reip_reg_11_ );
   nand U33267 ( n32237,n32242,n32243 );
   nand U33268 ( n32243,p3_phyaddrpointer_reg_11_,n32244 );
   nand U33269 ( n32242,n32245,n32246 );
   nor U33270 ( n32248,n32249,n32250 );
   nand U33271 ( n32250,n32251,n32252 );
   nand U33272 ( n32252,n31120,n28356 );
   nor U33273 ( n31120,n31152,n32253 );
   and U33274 ( n32253,n31139,n32254 );
   nand U33275 ( n32254,n32198,p3_instaddrpointer_reg_11_ );
   not U33276 ( n31152,n32255 );
   nand U33277 ( n32251,n31121,n28359 );
   nor U33278 ( n31121,n31150,n32256 );
   and U33279 ( n32256,n31139,n32257 );
   nand U33280 ( n32257,n32258,p3_instaddrpointer_reg_11_ );
   nor U33281 ( n32249,n31122,n28263 );
   xor U33282 ( n31122,n32259,n32260 );
   nor U33283 ( n32259,n32261,n32262 );
   nor U33284 ( n32247,n32263,n32264 );
   nand U33285 ( n32264,n32265,n32266 );
   nand U33286 ( n32266,n32006,p3_reip_reg_12_ );
   nand U33287 ( n32265,n32267,n32268 );
   nand U33288 ( n32263,n32269,n32270 );
   nand U33289 ( n32270,p3_phyaddrpointer_reg_12_,n32271 );
   nand U33290 ( n32271,n32272,n32273 );
   not U33291 ( n32273,n32244 );
   nand U33292 ( n32244,n32113,n32274 );
   nand U33293 ( n32274,n32042,n32275 );
   nor U33294 ( n32272,n32276,n32277 );
   and U33295 ( n32277,n32278,n32279 );
   nor U33296 ( n32276,p3_phyaddrpointer_reg_11_,n32280 );
   nand U33297 ( n32269,n32281,n32282 );
   nor U33298 ( n32281,n32283,n32246 );
   nor U33299 ( n32283,n32245,n32284 );
   nor U33300 ( n32284,n32278,n32285 );
   nor U33301 ( n32245,n28133,n32275 );
   nor U33302 ( n32287,n32288,n32289 );
   nand U33303 ( n32289,n32290,n32291 );
   nand U33304 ( n32291,p3_instaddrpointer_reg_13_,n32292 );
   nand U33305 ( n32290,n32293,n31933 );
   nand U33306 ( n32288,n32294,n32295 );
   nand U33307 ( n32295,n32296,n28356 );
   nor U33308 ( n32296,n31197,n32255 );
   nand U33309 ( n32294,n32297,n28359 );
   nor U33310 ( n32297,n31182,n32298 );
   nor U33311 ( n32286,n32299,n32300 );
   nand U33312 ( n32300,n32301,n32302 );
   or U33313 ( n32302,n31995,n31153 );
   nand U33314 ( n31153,n32303,n32304 );
   nand U33315 ( n32304,n32305,n32306 );
   xor U33316 ( n32306,n28177,p3_instaddrpointer_reg_13_ );
   nor U33317 ( n32305,n32262,n32307 );
   nor U33318 ( n32307,n32260,n32261 );
   nor U33319 ( n32261,n32152,p3_instaddrpointer_reg_12_ );
   nand U33320 ( n32303,n32308,n32309 );
   nand U33321 ( n32309,n32260,n32310 );
   not U33322 ( n32310,n32262 );
   nor U33323 ( n32260,n32311,n32312 );
   not U33324 ( n32312,n32313 );
   nor U33325 ( n32308,n32314,n32315 );
   nor U33326 ( n32315,n32316,n31159 );
   nor U33327 ( n32316,n28169,n31139 );
   nor U33328 ( n32314,p3_instaddrpointer_reg_13_,n32152 );
   nand U33329 ( n32301,n32006,p3_reip_reg_13_ );
   nand U33330 ( n32299,n32317,n32318 );
   nand U33331 ( n32318,p3_phyaddrpointer_reg_13_,n32319 );
   nand U33332 ( n32317,n32320,n32321 );
   nor U33333 ( n32323,n32324,n32325 );
   nand U33334 ( n32325,n32326,n32327 );
   nand U33335 ( n32327,n31956,n31200 );
   xor U33336 ( n31200,n32328,n32329 );
   xor U33337 ( n32328,n28175,p3_instaddrpointer_reg_14_ );
   nand U33338 ( n32326,n32006,p3_reip_reg_14_ );
   nor U33339 ( n32324,n32330,n32331 );
   nor U33340 ( n32322,n32332,n32333 );
   nand U33341 ( n32333,n32334,n32335 );
   nand U33342 ( n32335,p3_instaddrpointer_reg_14_,n32292 );
   nand U33343 ( n32292,n32336,n32337 );
   nand U33344 ( n32337,n32024,n31183 );
   nand U33345 ( n32336,n31955,n32338 );
   nand U33346 ( n32334,n32339,n31185 );
   nand U33347 ( n32339,n32340,n32341 );
   nand U33348 ( n32341,n32024,n31197 );
   nand U33349 ( n32340,n31955,n31182 );
   nand U33350 ( n32332,n32342,n32343 );
   nand U33351 ( n32343,p3_phyaddrpointer_reg_14_,n32344 );
   nand U33352 ( n32344,n32345,n32346 );
   not U33353 ( n32346,n32319 );
   nand U33354 ( n32319,n32113,n32347 );
   nand U33355 ( n32347,n32042,n32348 );
   nor U33356 ( n32345,n32349,n32350 );
   nor U33357 ( n32350,n32351,n32285 );
   nor U33358 ( n32349,p3_phyaddrpointer_reg_13_,n32280 );
   nand U33359 ( n32342,n32352,n32353 );
   nor U33360 ( n32352,n32354,n32321 );
   nor U33361 ( n32354,n32320,n32355 );
   nor U33362 ( n32355,n32285,n32356 );
   nor U33363 ( n32320,n32013,n32348 );
   nor U33364 ( n32358,n32359,n32360 );
   nand U33365 ( n32360,n32361,n32362 );
   nand U33366 ( n32362,p3_instaddrpointer_reg_14_,n32363 );
   nand U33367 ( n32363,n32364,n32365 );
   nand U33368 ( n32365,n32366,n28356 );
   nor U33369 ( n32366,n31239,n31183 );
   nand U33370 ( n32364,n32367,n28359 );
   nor U33371 ( n32367,n31238,n32338 );
   nand U33372 ( n32361,p3_instaddrpointer_reg_15_,n32368 );
   nor U33373 ( n32359,n31965,n32369 );
   nor U33374 ( n32357,n32370,n32371 );
   nand U33375 ( n32371,n32372,n32373 );
   nand U33376 ( n32373,n31956,n31205 );
   xor U33377 ( n31205,n32374,n32375 );
   xor U33378 ( n32374,n32131,p3_instaddrpointer_reg_15_ );
   nand U33379 ( n32372,n32006,p3_reip_reg_15_ );
   nand U33380 ( n32370,n32376,n32377 );
   nand U33381 ( n32377,p3_phyaddrpointer_reg_15_,n32378 );
   nand U33382 ( n32376,n32379,n32380 );
   nor U33383 ( n32382,n32383,n32384 );
   nand U33384 ( n32384,n32385,n32386 );
   nand U33385 ( n32386,n31956,n31259 );
   nand U33386 ( n31259,n32387,n32388 );
   nand U33387 ( n32388,n32389,n32152 );
   nand U33388 ( n32389,n32390,n32391 );
   nand U33389 ( n32387,n32392,n28177 );
   xor U33390 ( n32392,n31244,n32393 );
   nand U33391 ( n32385,n32006,p3_reip_reg_16_ );
   nor U33392 ( n32383,n32330,n32394 );
   nor U33393 ( n32381,n32395,n32396 );
   nand U33394 ( n32396,n32397,n32398 );
   nand U33395 ( n32398,p3_instaddrpointer_reg_16_,n32368 );
   nand U33396 ( n32368,n32399,n32400 );
   nand U33397 ( n32400,n32024,n31215 );
   nand U33398 ( n32399,n31955,n32401 );
   nand U33399 ( n32397,n32402,n31244 );
   nand U33400 ( n32402,n32403,n32404 );
   nand U33401 ( n32404,n32024,n31239 );
   nand U33402 ( n32403,n28359,n31238 );
   nand U33403 ( n32395,n32405,n32406 );
   nand U33404 ( n32406,p3_phyaddrpointer_reg_16_,n32407 );
   nand U33405 ( n32407,n32408,n32409 );
   not U33406 ( n32409,n32378 );
   nand U33407 ( n32378,n32113,n32410 );
   nand U33408 ( n32410,n32042,n32411 );
   nor U33409 ( n32408,n32412,n32413 );
   nor U33410 ( n32413,n32414,n32285 );
   nor U33411 ( n32412,p3_phyaddrpointer_reg_15_,n32280 );
   nand U33412 ( n32405,n32415,n32416 );
   nor U33413 ( n32415,n32417,n32380 );
   nor U33414 ( n32417,n32379,n32418 );
   nor U33415 ( n32418,n32285,n32419 );
   nor U33416 ( n32379,n28133,n32411 );
   nor U33417 ( n32421,n32422,n32423 );
   nand U33418 ( n32423,n32424,n32425 );
   nand U33419 ( n32425,p3_instaddrpointer_reg_17_,n32426 );
   nand U33420 ( n32424,n32427,n31933 );
   nand U33421 ( n32422,n32428,n32429 );
   nand U33422 ( n32429,n28356,n31266 );
   and U33423 ( n31266,n32430,n31239 );
   not U33424 ( n31239,n31215 );
   nor U33425 ( n32430,n31316,n31244 );
   nand U33426 ( n32428,n31955,n31267 );
   and U33427 ( n31267,n32431,n31238 );
   not U33428 ( n31238,n32401 );
   nor U33429 ( n32431,n31296,n31244 );
   nor U33430 ( n32420,n32432,n32433 );
   nand U33431 ( n32433,n32434,n32435 );
   or U33432 ( n32435,n31995,n31268 );
   nand U33433 ( n31268,n32436,n32437 );
   nand U33434 ( n32437,n32438,n32391 );
   nor U33435 ( n32438,n32439,n32440 );
   nor U33436 ( n32440,n32131,n32441 );
   nor U33437 ( n32441,n31274,n32390 );
   nor U33438 ( n32439,n32152,n31274 );
   nand U33439 ( n32436,n32442,n32390 );
   nor U33440 ( n32442,n32443,n32444 );
   nor U33441 ( n32444,n32445,n32152 );
   nor U33442 ( n32445,n32393,n31800 );
   nor U33443 ( n32443,n28175,n31274 );
   not U33444 ( n31274,p3_instaddrpointer_reg_17_ );
   nand U33445 ( n32434,n32006,p3_reip_reg_17_ );
   nand U33446 ( n32432,n32446,n32447 );
   nand U33447 ( n32447,p3_phyaddrpointer_reg_17_,n32448 );
   nand U33448 ( n32446,n32449,n32450 );
   nor U33449 ( n32449,n32013,n32451 );
   nor U33450 ( n32453,n32454,n32455 );
   nand U33451 ( n32455,n32456,n32457 );
   nand U33452 ( n32457,n31956,n31319 );
   xor U33453 ( n31319,n32458,n32459 );
   nor U33454 ( n32458,n32460,n32461 );
   nand U33455 ( n32456,n28349,p3_reip_reg_18_ );
   nor U33456 ( n32454,n32330,n32462 );
   nor U33457 ( n32452,n32463,n32464 );
   nand U33458 ( n32464,n32465,n32466 );
   nand U33459 ( n32466,p3_phyaddrpointer_reg_18_,n32467 );
   nand U33460 ( n32467,n32468,n32469 );
   not U33461 ( n32469,n32448 );
   nand U33462 ( n32448,n32113,n32470 );
   nand U33463 ( n32470,n32042,n32451 );
   nor U33464 ( n32468,n32471,n32472 );
   nor U33465 ( n32472,n32473,n32285 );
   nor U33466 ( n32471,p3_phyaddrpointer_reg_17_,n32013 );
   nand U33467 ( n32465,n32474,n32475 );
   not U33468 ( n32475,p3_phyaddrpointer_reg_18_ );
   nand U33469 ( n32474,n32476,n32477 );
   nand U33470 ( n32477,n32478,n32479 );
   not U33471 ( n32479,n32451 );
   nor U33472 ( n32478,n32013,n32450 );
   nand U33473 ( n32476,n32473,n32279 );
   nand U33474 ( n32463,n32480,n32481 );
   nand U33475 ( n32481,p3_instaddrpointer_reg_18_,n32426 );
   nand U33476 ( n32426,n32482,n32483 );
   nand U33477 ( n32483,n32024,n31297 );
   nand U33478 ( n32482,n31955,n32484 );
   nand U33479 ( n32480,n32485,n31299 );
   nand U33480 ( n32485,n32486,n32487 );
   nand U33481 ( n32487,n32024,n31316 );
   nand U33482 ( n32486,n28359,n31296 );
   nor U33483 ( n32489,n32490,n32491 );
   nand U33484 ( n32491,n32492,n32493 );
   nand U33485 ( n32493,p3_instaddrpointer_reg_18_,n32494 );
   nand U33486 ( n32494,n32495,n32496 );
   nand U33487 ( n32496,n32497,n28356 );
   nor U33488 ( n32497,n31377,n31297 );
   not U33489 ( n31297,n31316 );
   nand U33490 ( n32495,n32498,n28359 );
   nor U33491 ( n32498,n31363,n32484 );
   not U33492 ( n32484,n31296 );
   nand U33493 ( n32492,p3_instaddrpointer_reg_19_,n32499 );
   nor U33494 ( n32490,n31965,n32500 );
   nor U33495 ( n32488,n32501,n32502 );
   nand U33496 ( n32502,n32503,n32504 );
   or U33497 ( n32504,n31995,n31324 );
   xor U33498 ( n31324,n32505,n32506 );
   xor U33499 ( n32506,n31345,n32131 );
   nand U33500 ( n32503,n32006,p3_reip_reg_19_ );
   nand U33501 ( n32501,n32507,n32508 );
   nand U33502 ( n32508,p3_phyaddrpointer_reg_19_,n32509 );
   nand U33503 ( n32507,n32510,n32511 );
   nor U33504 ( n32510,n28134,n32512 );
   nor U33505 ( n32514,n32515,n32516 );
   nand U33506 ( n32516,n32517,n32518 );
   or U33507 ( n32518,n31995,n31380 );
   nand U33508 ( n31380,n32519,n32520 );
   nand U33509 ( n32520,n32521,n32522 );
   nand U33510 ( n32522,n32523,p3_instaddrpointer_reg_19_ );
   nor U33511 ( n32521,n32524,n32525 );
   nor U33512 ( n32525,n32131,n32526 );
   nor U33513 ( n32526,n31365,n32527 );
   nand U33514 ( n32527,n32505,n31345 );
   nor U33515 ( n32524,n28168,n31365 );
   nand U33516 ( n32519,n32528,n32529 );
   nand U33517 ( n32529,n32530,n31345 );
   nand U33518 ( n32530,n32523,n31365 );
   nor U33519 ( n32528,n32531,n32532 );
   nor U33520 ( n32532,n32533,n32152 );
   nor U33521 ( n32533,n32505,n31365 );
   not U33522 ( n32505,n32523 );
   nand U33523 ( n32517,n32006,p3_reip_reg_20_ );
   nor U33524 ( n32515,n32330,n32534 );
   nor U33525 ( n32513,n32535,n32536 );
   nand U33526 ( n32536,n32537,n32538 );
   nand U33527 ( n32538,p3_phyaddrpointer_reg_20_,n32539 );
   nand U33528 ( n32539,n32540,n32541 );
   not U33529 ( n32541,n32509 );
   nand U33530 ( n32509,n32113,n32542 );
   nand U33531 ( n32542,n32042,n32512 );
   nor U33532 ( n32540,n32543,n32544 );
   nor U33533 ( n32544,n32545,n32285 );
   nor U33534 ( n32543,p3_phyaddrpointer_reg_19_,n28133 );
   nand U33535 ( n32537,n32546,n32547 );
   not U33536 ( n32547,p3_phyaddrpointer_reg_20_ );
   nand U33537 ( n32546,n32548,n32549 );
   nand U33538 ( n32549,n32550,n32551 );
   not U33539 ( n32551,n32512 );
   nor U33540 ( n32550,n28133,n32511 );
   nand U33541 ( n32548,n32545,n32279 );
   nand U33542 ( n32535,n32552,n32553 );
   nand U33543 ( n32553,p3_instaddrpointer_reg_20_,n32499 );
   nand U33544 ( n32499,n32554,n32555 );
   nand U33545 ( n32555,n32024,n31334 );
   nand U33546 ( n32554,n31955,n32556 );
   nand U33547 ( n32552,n32557,n31365 );
   nand U33548 ( n32557,n32558,n32559 );
   nand U33549 ( n32559,n28356,n31377 );
   nand U33550 ( n32558,n28359,n31363 );
   nor U33551 ( n32561,n32562,n32563 );
   nand U33552 ( n32563,n32564,n32565 );
   nand U33553 ( n32565,p3_instaddrpointer_reg_21_,n32566 );
   nand U33554 ( n32564,n32567,n31933 );
   nand U33555 ( n32562,n32568,n32569 );
   nand U33556 ( n32569,n28356,n31387 );
   and U33557 ( n31387,n32570,n31377 );
   nor U33558 ( n32570,n32571,n31365 );
   nand U33559 ( n32568,n28359,n31388 );
   and U33560 ( n31388,n32572,n31363 );
   nor U33561 ( n32572,n31419,n31365 );
   nor U33562 ( n32560,n32573,n32574 );
   nand U33563 ( n32574,n32575,n32576 );
   nand U33564 ( n32576,n31956,n31389 );
   xor U33565 ( n31389,n28168,n32577 );
   xor U33566 ( n32577,p3_instaddrpointer_reg_21_,n32578 );
   nand U33567 ( n32578,n32579,n32580 );
   nand U33568 ( n32580,n32523,n32581 );
   nand U33569 ( n32581,n28175,n31821 );
   nand U33570 ( n31821,p3_instaddrpointer_reg_20_,p3_instaddrpointer_reg_19_ );
   nor U33571 ( n32523,n32460,n32582 );
   nor U33572 ( n32582,n32459,n32461 );
   nor U33573 ( n32460,n28168,p3_instaddrpointer_reg_18_ );
   nand U33574 ( n32579,n32152,n32583 );
   nand U33575 ( n32583,n31345,n31365 );
   nand U33576 ( n32575,n32006,p3_reip_reg_21_ );
   nand U33577 ( n32573,n32584,n32585 );
   nand U33578 ( n32585,p3_phyaddrpointer_reg_21_,n32586 );
   nand U33579 ( n32584,n32587,n32588 );
   nor U33580 ( n32587,n28134,n32589 );
   nor U33581 ( n32591,n32592,n32593 );
   nand U33582 ( n32593,n32594,n32595 );
   nand U33583 ( n32595,n31956,n31451 );
   xor U33584 ( n31451,n32596,n32597 );
   nand U33585 ( n32597,n32598,n32599 );
   nor U33586 ( n32596,n32600,n32601 );
   nor U33587 ( n32600,n28175,n31410 );
   nand U33588 ( n32594,n32006,p3_reip_reg_22_ );
   nor U33589 ( n32592,n32330,n32602 );
   nor U33590 ( n32590,n32603,n32604 );
   nand U33591 ( n32604,n32605,n32606 );
   nand U33592 ( n32606,p3_phyaddrpointer_reg_22_,n32607 );
   nand U33593 ( n32607,n32608,n32609 );
   not U33594 ( n32609,n32586 );
   nand U33595 ( n32586,n32113,n32610 );
   nand U33596 ( n32610,n32042,n32589 );
   nor U33597 ( n32608,n32611,n32612 );
   nor U33598 ( n32612,n32613,n32285 );
   nor U33599 ( n32611,p3_phyaddrpointer_reg_21_,n28134 );
   nand U33600 ( n32605,n32614,n32615 );
   not U33601 ( n32615,p3_phyaddrpointer_reg_22_ );
   nand U33602 ( n32614,n32616,n32617 );
   nand U33603 ( n32617,n32618,n32619 );
   not U33604 ( n32619,n32589 );
   nor U33605 ( n32618,n28133,n32588 );
   nand U33606 ( n32616,n32613,n32279 );
   nand U33607 ( n32603,n32620,n32621 );
   nand U33608 ( n32621,p3_instaddrpointer_reg_22_,n32566 );
   nand U33609 ( n32566,n32622,n32623 );
   nand U33610 ( n32623,n28356,n31416 );
   nand U33611 ( n32622,n28359,n32624 );
   nand U33612 ( n32620,n32625,n31410 );
   nand U33613 ( n32625,n32626,n32627 );
   nand U33614 ( n32627,n28356,n32571 );
   nand U33615 ( n32626,n28359,n31419 );
   nor U33616 ( n32629,n32630,n32631 );
   nand U33617 ( n32631,n32632,n32633 );
   nand U33618 ( n32633,p3_instaddrpointer_reg_23_,n32634 );
   nand U33619 ( n32632,n32635,n31933 );
   nand U33620 ( n32630,n32636,n32637 );
   nand U33621 ( n32637,n28356,n31458 );
   and U33622 ( n31458,n32638,n32571 );
   not U33623 ( n32571,n31416 );
   nor U33624 ( n32638,n32639,n31410 );
   nand U33625 ( n32636,n28359,n31459 );
   and U33626 ( n31459,n32640,n31419 );
   not U33627 ( n31419,n32624 );
   nor U33628 ( n32640,n31493,n31410 );
   nor U33629 ( n32628,n32641,n32642 );
   nand U33630 ( n32642,n32643,n32644 );
   nand U33631 ( n32644,n31956,n31460 );
   nand U33632 ( n31460,n32645,n32646 );
   nand U33633 ( n32646,n32647,p3_instaddrpointer_reg_23_ );
   nor U33634 ( n32647,n28177,n32648 );
   nor U33635 ( n32648,p3_instaddrpointer_reg_22_,n32649 );
   nor U33636 ( n32645,n32650,n32651 );
   nor U33637 ( n32651,n32652,n32653 );
   nand U33638 ( n32653,n32654,n32655 );
   and U33639 ( n32650,n32649,n32652 );
   nor U33640 ( n32652,n28169,p3_instaddrpointer_reg_23_ );
   nand U33641 ( n32649,n32598,n32655 );
   or U33642 ( n32655,n32599,n32601 );
   nor U33643 ( n32601,n32152,p3_instaddrpointer_reg_22_ );
   nand U33644 ( n32643,n28349,p3_reip_reg_23_ );
   nand U33645 ( n32641,n32656,n32657 );
   nand U33646 ( n32657,p3_phyaddrpointer_reg_23_,n32658 );
   nand U33647 ( n32656,n32659,n32660 );
   nor U33648 ( n32659,n28134,n32661 );
   nor U33649 ( n32663,n32664,n32665 );
   nand U33650 ( n32665,n32666,n32667 );
   or U33651 ( n32667,n31995,n31521 );
   xor U33652 ( n31521,n32668,n32669 );
   xor U33653 ( n32669,n31483,n28176 );
   nor U33654 ( n32668,n32670,n32671 );
   nor U33655 ( n32670,n32672,n32599 );
   nand U33656 ( n32666,n28349,p3_reip_reg_24_ );
   nor U33657 ( n32664,n32330,n32673 );
   nor U33658 ( n32662,n32674,n32675 );
   nand U33659 ( n32675,n32676,n32677 );
   nand U33660 ( n32677,p3_phyaddrpointer_reg_24_,n32678 );
   nand U33661 ( n32678,n32679,n32680 );
   not U33662 ( n32680,n32658 );
   nand U33663 ( n32658,n32113,n32681 );
   nand U33664 ( n32681,n32042,n32661 );
   nor U33665 ( n32679,n32682,n32683 );
   nor U33666 ( n32683,n32684,n32285 );
   nor U33667 ( n32682,p3_phyaddrpointer_reg_23_,n32013 );
   nand U33668 ( n32676,n32685,n32686 );
   not U33669 ( n32686,p3_phyaddrpointer_reg_24_ );
   nand U33670 ( n32685,n32687,n32688 );
   nand U33671 ( n32688,n32689,n32690 );
   not U33672 ( n32690,n32661 );
   nor U33673 ( n32689,n28133,n32660 );
   nand U33674 ( n32687,n32684,n32279 );
   nand U33675 ( n32674,n32691,n32692 );
   nand U33676 ( n32692,p3_instaddrpointer_reg_24_,n32634 );
   nand U33677 ( n32634,n32693,n32694 );
   nand U33678 ( n32694,n28356,n31490 );
   not U33679 ( n31490,n32639 );
   or U33680 ( n32693,n32178,n31493 );
   nand U33681 ( n32691,n32695,n31483 );
   nand U33682 ( n32695,n32696,n32697 );
   nand U33683 ( n32697,n28356,n32639 );
   nand U33684 ( n32696,n31955,n31493 );
   nor U33685 ( n32699,n32700,n32701 );
   nand U33686 ( n32701,n32702,n32703 );
   nand U33687 ( n32703,n31528,n28356 );
   nor U33688 ( n31528,n31554,n32704 );
   and U33689 ( n32704,n31541,n32705 );
   nand U33690 ( n32705,n32639,p3_instaddrpointer_reg_24_ );
   not U33691 ( n31554,n32706 );
   nand U33692 ( n32702,n31529,n28359 );
   nor U33693 ( n31529,n31552,n32707 );
   and U33694 ( n32707,n31541,n32708 );
   nand U33695 ( n32708,n31493,p3_instaddrpointer_reg_24_ );
   not U33696 ( n31552,n32709 );
   nor U33697 ( n32700,n31965,n32710 );
   not U33698 ( n32710,n32711 );
   nor U33699 ( n32698,n32712,n32713 );
   nand U33700 ( n32713,n32714,n32715 );
   or U33701 ( n32715,n31995,n31530 );
   xor U33702 ( n31530,n32716,n32717 );
   nor U33703 ( n32716,n32718,n32719 );
   nand U33704 ( n32714,n32006,p3_reip_reg_25_ );
   nand U33705 ( n32712,n32720,n32721 );
   nand U33706 ( n32721,p3_phyaddrpointer_reg_25_,n32722 );
   nand U33707 ( n32720,n32723,n32724 );
   nor U33708 ( n32723,n32013,n32725 );
   nor U33709 ( n32727,n32728,n32729 );
   nand U33710 ( n32729,n32730,n32731 );
   nand U33711 ( n32731,p3_instaddrpointer_reg_26_,n32732 );
   or U33712 ( n32730,n31995,n31556 );
   nand U33713 ( n31556,n32733,n32734 );
   nand U33714 ( n32734,n32735,n32736 );
   xor U33715 ( n32736,n28176,p3_instaddrpointer_reg_26_ );
   nor U33716 ( n32735,n32719,n32737 );
   nor U33717 ( n32737,n32717,n32718 );
   nor U33718 ( n32718,n28169,p3_instaddrpointer_reg_25_ );
   nand U33719 ( n32733,n32738,n32739 );
   or U33720 ( n32739,n32740,n32719 );
   nor U33721 ( n32738,n32741,n32742 );
   nor U33722 ( n32742,n32743,n31584 );
   nor U33723 ( n32743,n28168,n31541 );
   nor U33724 ( n32741,p3_instaddrpointer_reg_26_,n28168 );
   nand U33725 ( n32728,n32744,n32745 );
   nand U33726 ( n32745,n32746,n28356 );
   nor U33727 ( n32746,n31555,n32706 );
   nand U33728 ( n32744,n32747,n28359 );
   nor U33729 ( n32747,n31603,n32709 );
   nor U33730 ( n32726,n32748,n32749 );
   nand U33731 ( n32749,n32750,n32751 );
   nand U33732 ( n32751,n28349,p3_reip_reg_26_ );
   nand U33733 ( n32750,n32752,n32267 );
   nand U33734 ( n32748,n32753,n32754 );
   nand U33735 ( n32754,p3_phyaddrpointer_reg_26_,n32755 );
   nand U33736 ( n32755,n32756,n32757 );
   not U33737 ( n32757,n32722 );
   nand U33738 ( n32722,n32113,n32758 );
   nand U33739 ( n32758,n32042,n32725 );
   nor U33740 ( n32756,n32759,n32760 );
   nor U33741 ( n32760,n32761,n32285 );
   nor U33742 ( n32759,p3_phyaddrpointer_reg_25_,n28134 );
   nand U33743 ( n32753,n32762,n32763 );
   not U33744 ( n32763,p3_phyaddrpointer_reg_26_ );
   nand U33745 ( n32762,n32764,n32765 );
   nand U33746 ( n32765,n32766,n32767 );
   not U33747 ( n32767,n32725 );
   nor U33748 ( n32766,n28133,n32724 );
   nand U33749 ( n32764,n32761,n32279 );
   nor U33750 ( n32769,n32770,n32771 );
   nand U33751 ( n32771,n32772,n32773 );
   nand U33752 ( n32773,n32774,n31933 );
   not U33753 ( n31933,n31965 );
   nand U33754 ( n32772,n31956,n31615 );
   nand U33755 ( n31615,n32775,n32776 );
   nand U33756 ( n32776,n32777,n28168 );
   nand U33757 ( n32777,n32778,n32779 );
   nand U33758 ( n32775,n32780,n28175 );
   xor U33759 ( n32780,n32781,p3_instaddrpointer_reg_27_ );
   nor U33760 ( n32770,n28934,n31929 );
   not U33761 ( n31929,n32006 );
   nor U33762 ( n32768,n32782,n32783 );
   nand U33763 ( n32783,n32784,n32785 );
   nand U33764 ( n32785,p3_instaddrpointer_reg_27_,n32732 );
   nand U33765 ( n32732,n32786,n32787 );
   nand U33766 ( n32787,n32024,n31601 );
   not U33767 ( n31601,n31555 );
   or U33768 ( n32786,n32178,n31603 );
   nand U33769 ( n32784,n32788,n31595 );
   nand U33770 ( n32788,n32789,n32790 );
   nand U33771 ( n32790,n32024,n31555 );
   nand U33772 ( n32789,n31955,n31603 );
   nand U33773 ( n32782,n32791,n32792 );
   nand U33774 ( n32792,p3_phyaddrpointer_reg_27_,n32793 );
   nand U33775 ( n32791,n32794,n32795 );
   nor U33776 ( n32794,n28134,n32796 );
   nor U33777 ( n32798,n32799,n32800 );
   nand U33778 ( n32800,n32801,n32802 );
   nand U33779 ( n32802,n31622,n28356 );
   nor U33780 ( n31622,n31667,n32803 );
   and U33781 ( n32803,n31651,n32804 );
   nand U33782 ( n32804,n31555,p3_instaddrpointer_reg_27_ );
   not U33783 ( n31667,n32805 );
   nand U33784 ( n32801,n31623,n28359 );
   nor U33785 ( n31623,n31664,n32806 );
   and U33786 ( n32806,n31651,n32807 );
   nand U33787 ( n32807,n31603,p3_instaddrpointer_reg_27_ );
   not U33788 ( n31664,n32808 );
   nor U33789 ( n32799,n31624,n28263 );
   nand U33790 ( n31624,n32809,n32810 );
   nand U33791 ( n32810,n32811,n32779 );
   nor U33792 ( n32811,n32812,n32813 );
   nor U33793 ( n32813,n28176,n32814 );
   nor U33794 ( n32814,n31651,n32778 );
   nor U33795 ( n32812,n28168,n31651 );
   nand U33796 ( n32809,n32815,n32778 );
   nor U33797 ( n32815,n32816,n32817 );
   nor U33798 ( n32817,n32818,n28169 );
   and U33799 ( n32818,n32781,n31817 );
   nor U33800 ( n32816,n28176,n31651 );
   nor U33801 ( n32797,n32819,n32820 );
   nand U33802 ( n32820,n32821,n32822 );
   nand U33803 ( n32822,n28349,p3_reip_reg_28_ );
   nand U33804 ( n32821,n32823,n32267 );
   nand U33805 ( n32819,n32824,n32825 );
   nand U33806 ( n32825,p3_phyaddrpointer_reg_28_,n32826 );
   nand U33807 ( n32826,n32827,n32828 );
   not U33808 ( n32828,n32793 );
   nand U33809 ( n32793,n32113,n32829 );
   nand U33810 ( n32829,n32042,n32796 );
   nor U33811 ( n32827,n32830,n32831 );
   nor U33812 ( n32831,n32832,n32285 );
   nor U33813 ( n32830,p3_phyaddrpointer_reg_27_,n28134 );
   nand U33814 ( n32824,n32833,n32834 );
   not U33815 ( n32834,p3_phyaddrpointer_reg_28_ );
   nand U33816 ( n32833,n32835,n32836 );
   nand U33817 ( n32836,n32837,n32838 );
   not U33818 ( n32838,n32796 );
   nor U33819 ( n32837,n28134,n32795 );
   nand U33820 ( n32835,n32832,n32279 );
   nor U33821 ( n32840,n32841,n32842 );
   nand U33822 ( n32842,n32843,n32844 );
   nand U33823 ( n32844,p3_instaddrpointer_reg_29_,n32845 );
   or U33824 ( n32843,n32846,n31965 );
   nor U33825 ( n31965,n32267,n32279 );
   not U33826 ( n32267,n32330 );
   nand U33827 ( n32841,n32847,n32848 );
   nand U33828 ( n32848,n32849,n28356 );
   nor U33829 ( n32849,n31668,n32805 );
   nand U33830 ( n32847,n32850,n28359 );
   nor U33831 ( n32850,n31665,n32808 );
   nor U33832 ( n32839,n32851,n32852 );
   nand U33833 ( n32852,n32853,n32854 );
   or U33834 ( n32854,n31995,n31669 );
   xor U33835 ( n31669,n32855,n32856 );
   nor U33836 ( n32855,n32857,n32858 );
   nand U33837 ( n32853,n28349,p3_reip_reg_29_ );
   nand U33838 ( n32851,n32859,n32860 );
   nand U33839 ( n32860,n32861,n32862 );
   nor U33840 ( n32861,n32013,n32863 );
   nand U33841 ( n32859,n32864,p3_phyaddrpointer_reg_29_ );
   nor U33842 ( n32866,n32867,n32868 );
   nand U33843 ( n32868,n32869,n32870 );
   nand U33844 ( n32870,n31956,n31692 );
   xor U33845 ( n31692,n32871,n32872 );
   xor U33846 ( n32871,n28176,p3_instaddrpointer_reg_30_ );
   nand U33847 ( n32869,n28349,p3_reip_reg_30_ );
   nor U33848 ( n32867,n32330,n32873 );
   nor U33849 ( n32865,n32874,n32875 );
   nand U33850 ( n32875,n32876,n32877 );
   nand U33851 ( n32877,n32878,n32879 );
   nand U33852 ( n32876,p3_phyaddrpointer_reg_30_,n32880 );
   nand U33853 ( n32874,n32881,n32882 );
   nand U33854 ( n32882,p3_instaddrpointer_reg_30_,n32845 );
   nand U33855 ( n32845,n32883,n32884 );
   nand U33856 ( n32884,n32024,n31718 );
   nand U33857 ( n32883,n31955,n31706 );
   nand U33858 ( n32881,n32885,n31701 );
   nand U33859 ( n32885,n32886,n32887 );
   nand U33860 ( n32887,n32024,n31668 );
   nand U33861 ( n32886,n31955,n31665 );
   not U33862 ( n31955,n32178 );
   nor U33863 ( n32889,n32890,n32891 );
   nand U33864 ( n32891,n32892,n32893 );
   nand U33865 ( n32893,n32894,n31956 );
   not U33866 ( n31956,n31995 );
   nand U33867 ( n31995,n32895,n32896 );
   nor U33868 ( n32896,n29304,n31694 );
   and U33869 ( n32894,n31917,n31916 );
   nand U33870 ( n31916,n32897,n32898 );
   nand U33871 ( n32898,n32872,n31701 );
   not U33872 ( n32872,n32899 );
   nor U33873 ( n32897,n32900,n32901 );
   nor U33874 ( n32901,n32902,n28169 );
   nor U33875 ( n32902,n31701,n32903 );
   nand U33876 ( n32903,p3_instaddrpointer_reg_31_,n32899 );
   not U33877 ( n31701,p3_instaddrpointer_reg_30_ );
   nor U33878 ( n32900,n28177,n31898 );
   nand U33879 ( n31917,n32904,n32905 );
   nand U33880 ( n32905,p3_instaddrpointer_reg_30_,n32899 );
   nand U33881 ( n32899,n32906,n32907 );
   or U33882 ( n32907,n32857,n32856 );
   nor U33883 ( n32857,n32152,p3_instaddrpointer_reg_29_ );
   nor U33884 ( n32904,n32908,n32909 );
   nor U33885 ( n32909,n32131,n32910 );
   nor U33886 ( n32910,n31894,n32911 );
   nand U33887 ( n32911,n32856,n32906 );
   not U33888 ( n32906,n32858 );
   nor U33889 ( n32858,n31684,n28177 );
   and U33890 ( n32856,n32912,n32913 );
   nand U33891 ( n32913,p3_instaddrpointer_reg_28_,n32914 );
   nand U33892 ( n32914,n32131,n32779 );
   nand U33893 ( n32779,p3_instaddrpointer_reg_27_,n32781 );
   nand U33894 ( n32912,n32778,n28168 );
   nand U33895 ( n32778,n32915,n31595 );
   not U33896 ( n32915,n32781 );
   nand U33897 ( n32781,n32916,n32917 );
   nand U33898 ( n32917,n32740,n32152 );
   nor U33899 ( n32916,n32719,n32918 );
   nor U33900 ( n32918,n32919,n31584 );
   nor U33901 ( n32919,n32920,n28168 );
   nor U33902 ( n32920,n32717,n31541 );
   not U33903 ( n32717,n32740 );
   nand U33904 ( n32740,n32921,n32654 );
   not U33905 ( n32654,n32671 );
   nand U33906 ( n32671,n32598,n32922 );
   nand U33907 ( n32922,n28168,n32923 );
   nand U33908 ( n32923,n31410,n31473 );
   and U33909 ( n32598,n32924,n32925 );
   nand U33910 ( n32925,n28169,n32926 );
   nand U33911 ( n32926,n31345,n31401 );
   nor U33912 ( n32924,n32461,n32531 );
   nor U33913 ( n32531,n31365,n28175 );
   nor U33914 ( n32461,n31299,n28176 );
   nor U33915 ( n32921,n32927,n32928 );
   nor U33916 ( n32928,n28175,n31483 );
   nor U33917 ( n32927,n32599,n32929 );
   nand U33918 ( n32929,n32930,n32931 );
   not U33919 ( n32931,n32672 );
   nor U33920 ( n32672,n28168,n32932 );
   nand U33921 ( n32930,n28176,n31483 );
   nand U33922 ( n32599,n32933,n32459 );
   nand U33923 ( n32459,n32934,n32935 );
   nand U33924 ( n32935,p3_instaddrpointer_reg_17_,n32936 );
   nand U33925 ( n32936,n28176,n32391 );
   nand U33926 ( n32391,p3_instaddrpointer_reg_16_,n32937 );
   nand U33927 ( n32934,n32390,n28168 );
   nand U33928 ( n32390,n32393,n31244 );
   not U33929 ( n31244,p3_instaddrpointer_reg_16_ );
   not U33930 ( n32393,n32937 );
   nand U33931 ( n32937,n32938,n32939 );
   nand U33932 ( n32939,p3_instaddrpointer_reg_15_,n32940 );
   nand U33933 ( n32940,n32375,n28175 );
   not U33934 ( n32375,n32941 );
   nand U33935 ( n32938,n32941,n28169 );
   nand U33936 ( n32941,n32942,n32943 );
   nand U33937 ( n32943,p3_instaddrpointer_reg_14_,n32944 );
   nand U33938 ( n32944,n32329,n28176 );
   not U33939 ( n32329,n32945 );
   nand U33940 ( n32942,n32945,n28169 );
   nand U33941 ( n32945,n32946,n32947 );
   nor U33942 ( n32947,n32262,n32948 );
   nor U33943 ( n32948,n32949,n31159 );
   nor U33944 ( n32949,n32950,n28169 );
   nor U33945 ( n32950,n31139,n32313 );
   nor U33946 ( n32262,n31139,n28176 );
   nor U33947 ( n32946,n32951,n32311 );
   nand U33948 ( n32311,n32234,n32952 );
   nand U33949 ( n32952,p3_instaddrpointer_reg_11_,n28169 );
   nor U33950 ( n32234,n32176,n32953 );
   nor U33951 ( n32953,n31079,n28175 );
   not U33952 ( n31079,p3_instaddrpointer_reg_10_ );
   nor U33953 ( n32176,n31051,n32131 );
   nor U33954 ( n32951,n28177,n32313 );
   nand U33955 ( n32313,n32203,n32954 );
   nand U33956 ( n32954,n32131,n32955 );
   nand U33957 ( n32955,p3_instaddrpointer_reg_11_,p3_instaddrpointer_reg_10_ );
   nor U33958 ( n32203,n32175,n32177 );
   nor U33959 ( n32177,n28169,p3_instaddrpointer_reg_9_ );
   nand U33960 ( n32175,n32956,n32957 );
   nand U33961 ( n32957,n32958,n31032 );
   or U33962 ( n32958,n32149,n28176 );
   nand U33963 ( n32956,n28177,n32149 );
   nand U33964 ( n32149,n32959,n32960 );
   nand U33965 ( n32960,n32961,n31004 );
   nand U33966 ( n32961,n32130,n32152 );
   not U33967 ( n32130,n32962 );
   nand U33968 ( n32959,n28175,n32962 );
   nand U33969 ( n32962,n32096,n32963 );
   nand U33970 ( n32963,n32094,n32097 );
   nand U33971 ( n32094,n32060,n32964 );
   nand U33972 ( n32964,n32059,n32061 );
   not U33973 ( n32061,n32058 );
   nor U33974 ( n32058,n32965,n32966 );
   and U33975 ( n32965,n32967,n32968 );
   nand U33976 ( n32933,n32131,n32969 );
   nand U33977 ( n32969,n31798,n31799 );
   nor U33978 ( n32719,n31541,n28177 );
   not U33979 ( n32131,n32152 );
   nor U33980 ( n32908,n31898,n28168 );
   nand U33981 ( n32152,n32970,n32966 );
   nand U33982 ( n32892,n32024,n31909 );
   nand U33983 ( n31909,n32971,n31894 );
   nor U33984 ( n32971,n32972,n32973 );
   nor U33985 ( n32973,n31718,n31793 );
   not U33986 ( n31718,n31668 );
   nor U33987 ( n32972,n31668,n31898 );
   nor U33988 ( n31668,n32805,n31684 );
   nand U33989 ( n32805,n31817,n31555 );
   nor U33990 ( n31555,n32706,n31584 );
   nand U33991 ( n32706,n31796,n32639 );
   nor U33992 ( n32639,n31797,n31416 );
   nand U33993 ( n31416,n31798,n31377 );
   not U33994 ( n31377,n31334 );
   nand U33995 ( n31334,n31799,n31316 );
   nor U33996 ( n31316,n31800,n31215 );
   nand U33997 ( n31215,n32974,p3_instaddrpointer_reg_15_ );
   nor U33998 ( n32974,n31185,n31183 );
   not U33999 ( n31183,n31197 );
   nor U34000 ( n31197,n32255,n31159 );
   nand U34001 ( n32255,n31176,n32198 );
   and U34002 ( n32198,n32975,p3_instaddrpointer_reg_10_ );
   and U34003 ( n32975,n32173,p3_instaddrpointer_reg_9_ );
   nand U34004 ( n32173,n32976,n32977 );
   nand U34005 ( n32977,p3_instaddrpointer_reg_8_,n32978 );
   nand U34006 ( n32978,n32156,n32154 );
   or U34007 ( n32976,n32154,n32156 );
   nand U34008 ( n32156,n32979,n32980 );
   nand U34009 ( n32980,n32981,n31004 );
   nand U34010 ( n32981,n32127,n32128 );
   or U34011 ( n32979,n32128,n32127 );
   and U34012 ( n32127,n32982,n32983 );
   nand U34013 ( n32983,n32984,n30979 );
   or U34014 ( n32984,n32099,n32100 );
   nand U34015 ( n32982,n32099,n32100 );
   nand U34016 ( n32100,n32985,n32073 );
   nand U34017 ( n32073,n30949,n32986 );
   or U34018 ( n32986,n32987,n32988 );
   not U34019 ( n30949,p3_instaddrpointer_reg_5_ );
   nand U34020 ( n32985,n32074,n32068 );
   nand U34021 ( n32068,n32989,p3_instaddrpointer_reg_5_ );
   nor U34022 ( n32989,n32988,n32987 );
   and U34023 ( n32987,n32967,n32990 );
   and U34024 ( n32074,n32072,n32991 );
   or U34025 ( n32991,n32071,n32027 );
   nor U34026 ( n32027,n32992,p3_instaddrpointer_reg_4_ );
   nand U34027 ( n32071,n32993,n31988 );
   not U34028 ( n31988,n31983 );
   nor U34029 ( n31983,n32994,p3_instaddrpointer_reg_3_ );
   nand U34030 ( n32993,n31986,n31982 );
   nand U34031 ( n31982,p3_instaddrpointer_reg_3_,n32994 );
   xor U34032 ( n32994,n32995,n32996 );
   and U34033 ( n31986,n31963,n32997 );
   nand U34034 ( n32997,n31961,n31964 );
   or U34035 ( n31964,n32998,p3_instaddrpointer_reg_2_ );
   and U34036 ( n31961,n32999,n33000 );
   nand U34037 ( n33000,n33001,n30840 );
   nand U34038 ( n33001,n31940,n31939 );
   or U34039 ( n32999,n31939,n31940 );
   nor U34040 ( n31940,n33002,n28839 );
   not U34041 ( n28839,p3_instaddrpointer_reg_0_ );
   xor U34042 ( n31939,n31926,n33003 );
   nand U34043 ( n31963,p3_instaddrpointer_reg_2_,n32998 );
   nand U34044 ( n32998,n33004,n33005 );
   nand U34045 ( n33005,n33006,n33002 );
   nand U34046 ( n32072,n32992,p3_instaddrpointer_reg_4_ );
   xor U34047 ( n32992,n33007,n33008 );
   nand U34048 ( n33008,n33009,n33004 );
   xor U34049 ( n32099,n33010,n32988 );
   nand U34050 ( n32128,n33011,n33012 );
   nand U34051 ( n33012,n31915,n33013 );
   nand U34052 ( n33013,n32988,n33014 );
   nand U34053 ( n33011,n33015,n32988 );
   nand U34054 ( n32154,n32970,n32988 );
   nor U34055 ( n32988,n32990,n32967 );
   nand U34056 ( n32990,n33016,n33009 );
   nor U34057 ( n33016,n33007,n32996 );
   not U34058 ( n32996,n33004 );
   nand U34059 ( n33004,n33017,n33018 );
   nand U34060 ( n33018,n31942,n33002 );
   nor U34061 ( n32970,n31694,n33010 );
   not U34062 ( n32024,n31923 );
   nand U34063 ( n31923,n32895,n29304 );
   nor U34064 ( n32895,n31971,n28790 );
   nor U34065 ( n32890,n31913,n32178 );
   nand U34066 ( n32178,n33019,n33020 );
   nor U34067 ( n33020,n29304,n31971 );
   nor U34068 ( n33019,n28790,n31915 );
   and U34069 ( n31913,n33021,n31894 );
   not U34070 ( n31894,n31789 );
   nor U34071 ( n31789,n31898,p3_instaddrpointer_reg_30_ );
   nor U34072 ( n33021,n33022,n33023 );
   nor U34073 ( n33023,n31706,n31793 );
   nand U34074 ( n31793,p3_instaddrpointer_reg_30_,n31898 );
   not U34075 ( n31706,n31665 );
   nor U34076 ( n33022,n31665,n31898 );
   not U34077 ( n31898,p3_instaddrpointer_reg_31_ );
   nor U34078 ( n31665,n31684,n32808 );
   nand U34079 ( n32808,n31817,n31603 );
   nor U34080 ( n31603,n31584,n32709 );
   nand U34081 ( n32709,n31796,n31493 );
   nor U34082 ( n31493,n31797,n32624 );
   nand U34083 ( n32624,n31798,n31363 );
   not U34084 ( n31363,n32556 );
   nand U34085 ( n32556,n31799,n31296 );
   nor U34086 ( n31296,n31800,n32401 );
   nand U34087 ( n32401,n33024,p3_instaddrpointer_reg_15_ );
   nor U34088 ( n33024,n31185,n32338 );
   not U34089 ( n32338,n31182 );
   nor U34090 ( n31182,n31159,n32298 );
   not U34091 ( n32298,n31150 );
   nor U34092 ( n31150,n31193,n32205 );
   not U34093 ( n32205,n32258 );
   nor U34094 ( n32258,n31803,n32180 );
   nand U34095 ( n32180,n33025,n33026 );
   nand U34096 ( n33026,n33027,n31004 );
   not U34097 ( n31004,p3_instaddrpointer_reg_7_ );
   or U34098 ( n33027,n32124,n32125 );
   nand U34099 ( n33025,n32124,n32125 );
   nand U34100 ( n32125,n33015,n32966 );
   nor U34101 ( n33015,n31915,n33010 );
   nand U34102 ( n32124,n32096,n33028 );
   nand U34103 ( n33028,n32097,n32095 );
   nand U34104 ( n32095,n32060,n33029 );
   nand U34105 ( n33029,n32052,n32059 );
   nand U34106 ( n32059,p3_instaddrpointer_reg_5_,n32062 );
   not U34107 ( n32052,n32054 );
   xor U34108 ( n32054,n32967,n32968 );
   or U34109 ( n32060,n32062,p3_instaddrpointer_reg_5_ );
   nand U34110 ( n32062,n32031,n33030 );
   nand U34111 ( n33030,n32029,n32030 );
   nand U34112 ( n32030,n33031,n30925 );
   not U34113 ( n30925,p3_instaddrpointer_reg_4_ );
   not U34114 ( n32029,n32023 );
   nor U34115 ( n32023,n31993,n32000 );
   nor U34116 ( n32000,n30897,n33032 );
   nor U34117 ( n31993,n31991,n33033 );
   not U34118 ( n33033,n31999 );
   nand U34119 ( n31999,n33032,n30897 );
   not U34120 ( n30897,p3_instaddrpointer_reg_3_ );
   xor U34121 ( n33032,n32995,n33006 );
   nand U34122 ( n31991,n31959,n33034 );
   nand U34123 ( n33034,n31960,n31957 );
   nand U34124 ( n31957,n33035,n33036 );
   nand U34125 ( n33036,n33037,n30840 );
   not U34126 ( n30840,p3_instaddrpointer_reg_1_ );
   or U34127 ( n33037,n31924,n31942 );
   nand U34128 ( n33035,n31942,n31924 );
   nand U34129 ( n31924,p3_instaddrpointer_reg_0_,n33002 );
   nand U34130 ( n31960,n33038,p3_instaddrpointer_reg_2_ );
   nor U34131 ( n33038,n33006,n33039 );
   nor U34132 ( n33039,n31942,n33040 );
   nand U34133 ( n31959,n30866,n33041 );
   nand U34134 ( n33041,n33042,n33043 );
   not U34135 ( n33043,n33006 );
   nand U34136 ( n33042,n33017,n33003 );
   not U34137 ( n30866,p3_instaddrpointer_reg_2_ );
   nand U34138 ( n32031,p3_instaddrpointer_reg_4_,n33044 );
   not U34139 ( n33044,n33031 );
   nand U34140 ( n33031,n33045,n32968 );
   nand U34141 ( n33045,n33007,n33046 );
   nand U34142 ( n33046,n33006,n33009 );
   nand U34143 ( n32097,n33047,p3_instaddrpointer_reg_6_ );
   xor U34144 ( n33047,n33014,n32966 );
   nand U34145 ( n32096,n33048,n30979 );
   not U34146 ( n30979,p3_instaddrpointer_reg_6_ );
   xor U34147 ( n33048,n33010,n32966 );
   nor U34148 ( n32966,n32968,n32967 );
   nand U34149 ( n32968,n33049,n33006 );
   nor U34150 ( n33006,n33003,n33017 );
   nor U34151 ( n33049,n33007,n32995 );
   nand U34152 ( n31803,n33050,p3_instaddrpointer_reg_10_ );
   nor U34153 ( n33050,n31032,n31051 );
   not U34154 ( n31051,p3_instaddrpointer_reg_9_ );
   not U34155 ( n31032,p3_instaddrpointer_reg_8_ );
   not U34156 ( n31193,n31176 );
   nor U34157 ( n31176,n31139,n31108 );
   not U34158 ( n31108,p3_instaddrpointer_reg_11_ );
   not U34159 ( n31139,p3_instaddrpointer_reg_12_ );
   not U34160 ( n31159,p3_instaddrpointer_reg_13_ );
   not U34161 ( n31185,p3_instaddrpointer_reg_14_ );
   nand U34162 ( n31800,p3_instaddrpointer_reg_17_,p3_instaddrpointer_reg_16_ );
   nor U34163 ( n31799,n31345,n31299 );
   not U34164 ( n31299,p3_instaddrpointer_reg_18_ );
   not U34165 ( n31345,p3_instaddrpointer_reg_19_ );
   nor U34166 ( n31798,n31401,n31365 );
   not U34167 ( n31365,p3_instaddrpointer_reg_20_ );
   not U34168 ( n31401,p3_instaddrpointer_reg_21_ );
   not U34169 ( n31797,n32932 );
   nor U34170 ( n32932,n31473,n31410 );
   not U34171 ( n31410,p3_instaddrpointer_reg_22_ );
   not U34172 ( n31473,p3_instaddrpointer_reg_23_ );
   nor U34173 ( n31796,n31541,n31483 );
   not U34174 ( n31483,p3_instaddrpointer_reg_24_ );
   not U34175 ( n31541,p3_instaddrpointer_reg_25_ );
   not U34176 ( n31584,p3_instaddrpointer_reg_26_ );
   nor U34177 ( n31817,n31651,n31595 );
   not U34178 ( n31595,p3_instaddrpointer_reg_27_ );
   not U34179 ( n31651,p3_instaddrpointer_reg_28_ );
   not U34180 ( n31684,p3_instaddrpointer_reg_29_ );
   nor U34181 ( n32888,n33051,n33052 );
   nand U34182 ( n33052,n33053,n33054 );
   nand U34183 ( n33054,n28349,p3_reip_reg_31_ );
   nor U34184 ( n32006,n28796,n31971 );
   or U34185 ( n33053,n32330,n33055 );
   nand U34186 ( n32330,n33056,p3_state2_reg_1_ );
   nor U34187 ( n33056,p3_statebs16_reg,n31971 );
   nand U34188 ( n33051,n33057,n33058 );
   nand U34189 ( n33058,p3_phyaddrpointer_reg_31_,n33059 );
   nand U34190 ( n33059,n33060,n33061 );
   or U34191 ( n33061,n32280,p3_phyaddrpointer_reg_30_ );
   not U34192 ( n33060,n32880 );
   nand U34193 ( n32880,n33062,n33063 );
   nand U34194 ( n33063,n32279,n33064 );
   nor U34195 ( n33062,n32864,n33065 );
   nor U34196 ( n33065,p3_phyaddrpointer_reg_29_,n32280 );
   nor U34197 ( n32280,n32279,n32042 );
   not U34198 ( n32042,n32013 );
   and U34199 ( n32864,n31932,n33066 );
   nand U34200 ( n33066,n33067,n32113 );
   nand U34201 ( n31932,n32113,n32013 );
   nand U34202 ( n33057,n33068,n33069 );
   and U34203 ( n33068,n32878,p3_phyaddrpointer_reg_30_ );
   nand U34204 ( n32878,n33070,n33071 );
   nand U34205 ( n33071,n33072,n33067 );
   not U34206 ( n33067,n32863 );
   nand U34207 ( n32863,n33073,p3_phyaddrpointer_reg_28_ );
   nor U34208 ( n33073,n32795,n32796 );
   nand U34209 ( n32796,n33074,p3_phyaddrpointer_reg_26_ );
   nor U34210 ( n33074,n32724,n32725 );
   nand U34211 ( n32725,n33075,p3_phyaddrpointer_reg_24_ );
   nor U34212 ( n33075,n32660,n32661 );
   nand U34213 ( n32661,n33076,p3_phyaddrpointer_reg_22_ );
   nor U34214 ( n33076,n32588,n32589 );
   nand U34215 ( n32589,n33077,p3_phyaddrpointer_reg_20_ );
   nor U34216 ( n33077,n32511,n32512 );
   nand U34217 ( n32512,n33078,p3_phyaddrpointer_reg_18_ );
   nor U34218 ( n33078,n32450,n32451 );
   nand U34219 ( n32451,n33079,p3_phyaddrpointer_reg_16_ );
   nor U34220 ( n33079,n32380,n32411 );
   nand U34221 ( n32411,n33080,p3_phyaddrpointer_reg_14_ );
   nor U34222 ( n33080,n32321,n32348 );
   nand U34223 ( n32348,n33081,p3_phyaddrpointer_reg_12_ );
   nor U34224 ( n33081,n32246,n32275 );
   nand U34225 ( n32275,n33082,n33083 );
   nor U34226 ( n33083,n32165,n33084 );
   nand U34227 ( n33084,n32225,p3_phyaddrpointer_reg_7_ );
   not U34228 ( n32225,n32142 );
   nand U34229 ( n32142,n33085,p3_phyaddrpointer_reg_6_ );
   nor U34230 ( n33085,n32086,n32085 );
   nor U34231 ( n33082,n32190,n32222 );
   not U34232 ( n32321,p3_phyaddrpointer_reg_13_ );
   nor U34233 ( n33072,n28133,n32862 );
   nand U34234 ( n32013,n33086,p3_statebs16_reg );
   nor U34235 ( n33086,n31971,n28856 );
   nand U34236 ( n33070,n33087,n32279 );
   not U34237 ( n32279,n32285 );
   nand U34238 ( n32285,n33088,p3_state2_reg_2_ );
   nor U34239 ( n33088,p3_state2_reg_0_,n31971 );
   not U34240 ( n31971,n32113 );
   nand U34241 ( n32113,n33089,n33090 );
   or U34242 ( n33090,n30796,p3_state2_reg_0_ );
   nor U34243 ( n30796,n28795,n28866 );
   nor U34244 ( n28866,p3_state2_reg_1_,p3_state2_reg_3_ );
   nand U34245 ( n33092,p3_lword_reg_15_,n28335 );
   nor U34246 ( n33091,n33094,n33095 );
   nor U34247 ( n33095,n28145,n33096 );
   nor U34248 ( n33094,n33097,n33098 );
   nand U34249 ( n33100,p3_lword_reg_14_,n28335 );
   nor U34250 ( n33099,n33101,n33102 );
   nor U34251 ( n33102,n28144,n33103 );
   nand U34252 ( n33105,p3_lword_reg_13_,n33093 );
   nor U34253 ( n33104,n33106,n33107 );
   nor U34254 ( n33107,n28144,n33108 );
   nand U34255 ( n33110,p3_lword_reg_12_,n33093 );
   nor U34256 ( n33109,n33111,n33112 );
   nor U34257 ( n33112,n28146,n33113 );
   nand U34258 ( n33115,p3_lword_reg_11_,n33093 );
   nor U34259 ( n33114,n33116,n33117 );
   nor U34260 ( n33117,n28146,n33118 );
   nand U34261 ( n33120,p3_lword_reg_10_,n33093 );
   nor U34262 ( n33119,n33121,n33122 );
   nor U34263 ( n33122,n28143,n33123 );
   nand U34264 ( n33125,p3_lword_reg_9_,n33093 );
   nor U34265 ( n33124,n33126,n33127 );
   nor U34266 ( n33127,n28143,n33128 );
   nand U34267 ( n33130,p3_lword_reg_8_,n33093 );
   nor U34268 ( n33129,n33131,n33132 );
   nor U34269 ( n33132,n28145,n33133 );
   nand U34270 ( n33135,p3_lword_reg_7_,n33093 );
   nor U34271 ( n33134,n33136,n33137 );
   nor U34272 ( n33137,n28145,n33138 );
   nand U34273 ( n33140,p3_lword_reg_6_,n33093 );
   nor U34274 ( n33139,n33141,n33142 );
   nor U34275 ( n33142,n28144,n33143 );
   nand U34276 ( n33145,p3_lword_reg_5_,n33093 );
   nor U34277 ( n33144,n33146,n33147 );
   nor U34278 ( n33147,n28144,n33148 );
   nand U34279 ( n33150,p3_lword_reg_4_,n33093 );
   nor U34280 ( n33149,n33151,n33152 );
   nor U34281 ( n33152,n28146,n33153 );
   nand U34282 ( n33155,p3_lword_reg_3_,n33093 );
   nor U34283 ( n33154,n33156,n33157 );
   nor U34284 ( n33157,n28143,n33158 );
   nand U34285 ( n33160,p3_lword_reg_2_,n33093 );
   nor U34286 ( n33159,n33161,n33162 );
   nor U34287 ( n33162,n28143,n33163 );
   nand U34288 ( n33165,p3_lword_reg_1_,n33093 );
   nor U34289 ( n33164,n33166,n33167 );
   nor U34290 ( n33167,n28145,n33168 );
   nand U34291 ( n33170,p3_lword_reg_0_,n33093 );
   nor U34292 ( n33169,n33171,n33172 );
   nor U34293 ( n33172,n28145,n33173 );
   nand U34294 ( n33175,p3_uword_reg_14_,n33093 );
   nor U34295 ( n33174,n33101,n33176 );
   nor U34296 ( n33176,n28143,n33177 );
   nor U34297 ( n33101,n33178,n28254 );
   nand U34298 ( n33180,p3_uword_reg_13_,n33093 );
   nor U34299 ( n33179,n33106,n33181 );
   nor U34300 ( n33181,n28143,n33182 );
   nor U34301 ( n33106,n33183,n28254 );
   nand U34302 ( n33185,p3_uword_reg_12_,n33093 );
   nor U34303 ( n33184,n33111,n33186 );
   nor U34304 ( n33186,n28145,n33187 );
   nor U34305 ( n33111,n33188,n28254 );
   nand U34306 ( n33190,p3_uword_reg_11_,n33093 );
   nor U34307 ( n33189,n33116,n33191 );
   nor U34308 ( n33191,n28144,n33192 );
   nor U34309 ( n33116,n33193,n33098 );
   nand U34310 ( n33195,p3_uword_reg_10_,n33093 );
   nor U34311 ( n33194,n33121,n33196 );
   nor U34312 ( n33196,n28144,n33197 );
   nor U34313 ( n33121,n33198,n33098 );
   nand U34314 ( n33200,p3_uword_reg_9_,n28335 );
   nor U34315 ( n33199,n33126,n33201 );
   nor U34316 ( n33201,n28146,n33202 );
   nor U34317 ( n33126,n33203,n33098 );
   nand U34318 ( n33205,p3_uword_reg_8_,n28335 );
   nor U34319 ( n33204,n33131,n33206 );
   nor U34320 ( n33206,n28146,n33207 );
   nor U34321 ( n33131,n33208,n33098 );
   nand U34322 ( n33210,p3_uword_reg_7_,n28335 );
   nor U34323 ( n33209,n33136,n33211 );
   nor U34324 ( n33211,n28143,n33212 );
   nor U34325 ( n33136,n30643,n33098 );
   nand U34326 ( n33214,p3_uword_reg_6_,n28335 );
   nor U34327 ( n33213,n33141,n33215 );
   nor U34328 ( n33215,n28143,n33216 );
   nor U34329 ( n33141,n30658,n33098 );
   nand U34330 ( n33218,p3_uword_reg_5_,n28335 );
   nor U34331 ( n33217,n33146,n33219 );
   nor U34332 ( n33219,n28145,n33220 );
   nor U34333 ( n33146,n30669,n33098 );
   nand U34334 ( n33222,p3_uword_reg_4_,n28335 );
   nor U34335 ( n33221,n33151,n33223 );
   nor U34336 ( n33223,n28145,n33224 );
   nor U34337 ( n33151,n30680,n33098 );
   nand U34338 ( n33226,p3_uword_reg_3_,n28335 );
   nor U34339 ( n33225,n33156,n33227 );
   nor U34340 ( n33227,n28144,n33228 );
   nor U34341 ( n33156,n30690,n33098 );
   nand U34342 ( n33230,p3_uword_reg_2_,n28335 );
   nor U34343 ( n33229,n33161,n33231 );
   nor U34344 ( n33231,n28144,n33232 );
   nor U34345 ( n33161,n30701,n33098 );
   nand U34346 ( n33234,p3_uword_reg_1_,n28335 );
   nor U34347 ( n33233,n33166,n33235 );
   nor U34348 ( n33235,n28146,n33236 );
   nor U34349 ( n33166,n30712,n28254 );
   nand U34350 ( n33238,p3_uword_reg_0_,n28335 );
   nor U34351 ( n33237,n33171,n33239 );
   nor U34352 ( n33239,n28146,n33240 );
   nor U34353 ( n33171,n30737,n33098 );
   nand U34354 ( n33098,n33241,n29366 );
   not U34355 ( n33241,n33093 );
   nand U34356 ( n33093,n33242,n31747 );
   nor U34357 ( n33242,n33243,n29211 );
   nor U34358 ( n33243,n31731,n33244 );
   nor U34359 ( n33244,n28801,n33245 );
   not U34360 ( n31731,n29187 );
   nand U34361 ( n33247,p3_datao_reg_0_,n28332 );
   nor U34362 ( n33246,n33249,n33250 );
   nor U34363 ( n33250,n33173,n33251 );
   nor U34364 ( n33249,n33252,n28111 );
   not U34365 ( n33252,p3_lword_reg_0_ );
   nand U34366 ( n33255,p3_datao_reg_1_,n28332 );
   nor U34367 ( n33254,n33256,n33257 );
   nor U34368 ( n33257,n33168,n33251 );
   nor U34369 ( n33256,n33258,n28111 );
   not U34370 ( n33258,p3_lword_reg_1_ );
   nand U34371 ( n33260,p3_datao_reg_2_,n33248 );
   nor U34372 ( n33259,n33261,n33262 );
   nor U34373 ( n33262,n33163,n33251 );
   nor U34374 ( n33261,n33263,n28112 );
   not U34375 ( n33263,p3_lword_reg_2_ );
   nand U34376 ( n33265,p3_datao_reg_3_,n33248 );
   nor U34377 ( n33264,n33266,n33267 );
   nor U34378 ( n33267,n33158,n33251 );
   nor U34379 ( n33266,n33268,n33253 );
   not U34380 ( n33268,p3_lword_reg_3_ );
   nand U34381 ( n33270,p3_datao_reg_4_,n33248 );
   nor U34382 ( n33269,n33271,n33272 );
   nor U34383 ( n33272,n33153,n28257 );
   nor U34384 ( n33271,n33273,n28111 );
   not U34385 ( n33273,p3_lword_reg_4_ );
   nand U34386 ( n33275,p3_datao_reg_5_,n33248 );
   nor U34387 ( n33274,n33276,n33277 );
   nor U34388 ( n33277,n33148,n28257 );
   nor U34389 ( n33276,n33278,n28112 );
   not U34390 ( n33278,p3_lword_reg_5_ );
   nand U34391 ( n33280,p3_datao_reg_6_,n33248 );
   nor U34392 ( n33279,n33281,n33282 );
   nor U34393 ( n33282,n33143,n33251 );
   nor U34394 ( n33281,n33283,n33253 );
   not U34395 ( n33283,p3_lword_reg_6_ );
   nand U34396 ( n33285,p3_datao_reg_7_,n33248 );
   nor U34397 ( n33284,n33286,n33287 );
   nor U34398 ( n33287,n33138,n33251 );
   nor U34399 ( n33286,n33288,n28111 );
   not U34400 ( n33288,p3_lword_reg_7_ );
   nand U34401 ( n33290,p3_datao_reg_8_,n33248 );
   nor U34402 ( n33289,n33291,n33292 );
   nor U34403 ( n33292,n33133,n33251 );
   nor U34404 ( n33291,n33293,n28112 );
   not U34405 ( n33293,p3_lword_reg_8_ );
   nand U34406 ( n33295,p3_datao_reg_9_,n33248 );
   nor U34407 ( n33294,n33296,n33297 );
   nor U34408 ( n33297,n33128,n28257 );
   nor U34409 ( n33296,n33298,n33253 );
   not U34410 ( n33298,p3_lword_reg_9_ );
   nand U34411 ( n33300,p3_datao_reg_10_,n33248 );
   nor U34412 ( n33299,n33301,n33302 );
   nor U34413 ( n33302,n33123,n33251 );
   nor U34414 ( n33301,n33303,n28111 );
   not U34415 ( n33303,p3_lword_reg_10_ );
   nand U34416 ( n33305,p3_datao_reg_11_,n33248 );
   nor U34417 ( n33304,n33306,n33307 );
   nor U34418 ( n33307,n33118,n33251 );
   nor U34419 ( n33306,n33308,n28112 );
   not U34420 ( n33308,p3_lword_reg_11_ );
   nand U34421 ( n33310,p3_datao_reg_12_,n33248 );
   nor U34422 ( n33309,n33311,n33312 );
   nor U34423 ( n33312,n33113,n33251 );
   nor U34424 ( n33311,n33313,n33253 );
   not U34425 ( n33313,p3_lword_reg_12_ );
   nand U34426 ( n33315,p3_datao_reg_13_,n33248 );
   nor U34427 ( n33314,n33316,n33317 );
   nor U34428 ( n33317,n33108,n28257 );
   nor U34429 ( n33316,n33318,n28111 );
   not U34430 ( n33318,p3_lword_reg_13_ );
   nand U34431 ( n33320,p3_datao_reg_14_,n33248 );
   nor U34432 ( n33319,n33321,n33322 );
   nor U34433 ( n33322,n33103,n33251 );
   nor U34434 ( n33321,n33323,n33253 );
   not U34435 ( n33323,p3_lword_reg_14_ );
   nand U34436 ( n33325,p3_datao_reg_15_,n33248 );
   nor U34437 ( n33324,n33326,n33327 );
   nor U34438 ( n33327,n33096,n28257 );
   nor U34439 ( n33326,n33328,n28112 );
   not U34440 ( n33328,p3_lword_reg_15_ );
   nand U34441 ( n33330,p3_datao_reg_16_,n33248 );
   nor U34442 ( n33329,n33331,n33332 );
   nor U34443 ( n33332,n33240,n28298 );
   nor U34444 ( n33331,n33333,n28111 );
   not U34445 ( n33333,p3_uword_reg_0_ );
   nand U34446 ( n33335,p3_datao_reg_17_,n33248 );
   nor U34447 ( n33334,n33336,n33337 );
   nor U34448 ( n33337,n33236,n28298 );
   nor U34449 ( n33336,n33338,n33253 );
   not U34450 ( n33338,p3_uword_reg_1_ );
   nand U34451 ( n33340,p3_datao_reg_18_,n33248 );
   nor U34452 ( n33339,n33341,n33342 );
   nor U34453 ( n33342,n33232,n28299 );
   nor U34454 ( n33341,n33343,n28112 );
   not U34455 ( n33343,p3_uword_reg_2_ );
   nand U34456 ( n33345,p3_datao_reg_19_,n33248 );
   nor U34457 ( n33344,n33346,n33347 );
   nor U34458 ( n33347,n33228,n28299 );
   nor U34459 ( n33346,n33348,n33253 );
   not U34460 ( n33348,p3_uword_reg_3_ );
   nand U34461 ( n33350,p3_datao_reg_20_,n33248 );
   nor U34462 ( n33349,n33351,n33352 );
   nor U34463 ( n33352,n33224,n28298 );
   nor U34464 ( n33351,n33353,n28111 );
   not U34465 ( n33353,p3_uword_reg_4_ );
   nand U34466 ( n33355,p3_datao_reg_21_,n33248 );
   nor U34467 ( n33354,n33356,n33357 );
   nor U34468 ( n33357,n33220,n28298 );
   nor U34469 ( n33356,n33358,n28112 );
   not U34470 ( n33358,p3_uword_reg_5_ );
   nand U34471 ( n33360,p3_datao_reg_22_,n33248 );
   nor U34472 ( n33359,n33361,n33362 );
   nor U34473 ( n33362,n33216,n28299 );
   nor U34474 ( n33361,n33363,n33253 );
   not U34475 ( n33363,p3_uword_reg_6_ );
   nand U34476 ( n33365,p3_datao_reg_23_,n33248 );
   nor U34477 ( n33364,n33366,n33367 );
   nor U34478 ( n33367,n33212,n28299 );
   nor U34479 ( n33366,n33368,n28111 );
   not U34480 ( n33368,p3_uword_reg_7_ );
   nand U34481 ( n33370,p3_datao_reg_24_,n28332 );
   nor U34482 ( n33369,n33371,n33372 );
   nor U34483 ( n33372,n33207,n28299 );
   nor U34484 ( n33371,n33373,n28112 );
   not U34485 ( n33373,p3_uword_reg_8_ );
   nand U34486 ( n33375,p3_datao_reg_25_,n28332 );
   nor U34487 ( n33374,n33376,n33377 );
   nor U34488 ( n33377,n33202,n28298 );
   nor U34489 ( n33376,n33378,n33253 );
   not U34490 ( n33378,p3_uword_reg_9_ );
   nand U34491 ( n33380,p3_datao_reg_26_,n28332 );
   nor U34492 ( n33379,n33381,n33382 );
   nor U34493 ( n33382,n33197,n28298 );
   nor U34494 ( n33381,n33383,n28111 );
   not U34495 ( n33383,p3_uword_reg_10_ );
   nand U34496 ( n33385,p3_datao_reg_27_,n28332 );
   nor U34497 ( n33384,n33386,n33387 );
   nor U34498 ( n33387,n33192,n28299 );
   nor U34499 ( n33386,n33388,n28112 );
   not U34500 ( n33388,p3_uword_reg_11_ );
   nand U34501 ( n33390,p3_datao_reg_28_,n28332 );
   nor U34502 ( n33389,n33391,n33392 );
   nor U34503 ( n33392,n33187,n28299 );
   nor U34504 ( n33391,n33393,n33253 );
   not U34505 ( n33393,p3_uword_reg_12_ );
   nand U34506 ( n33395,p3_datao_reg_29_,n28332 );
   nor U34507 ( n33394,n33396,n33397 );
   nor U34508 ( n33397,n33182,n28298 );
   nor U34509 ( n33396,n33398,n28111 );
   not U34510 ( n33398,p3_uword_reg_13_ );
   nand U34511 ( n33400,n33248,p3_datao_reg_30_ );
   not U34512 ( n33248,n33401 );
   nor U34513 ( n33399,n33402,n33403 );
   nor U34514 ( n33403,n33177,n28298 );
   nand U34515 ( n33251,p3_state2_reg_0_,n33401 );
   nor U34516 ( n33402,n33404,n28112 );
   nand U34517 ( n33253,n28790,n33401 );
   not U34518 ( n33404,p3_uword_reg_14_ );
   not U34519 ( n28475,p3_datao_reg_31_ );
   nand U34520 ( n33401,n33405,n33406 );
   nand U34521 ( n33406,n33407,n33408 );
   not U34522 ( n33408,n29374 );
   nor U34523 ( n33407,n28815,n28805 );
   not U34524 ( n28815,n31747 );
   nand U34525 ( n33405,n28793,n28790 );
   nor U34526 ( n28793,n28856,n28808 );
   nor U34527 ( n33410,n33411,n33412 );
   nor U34528 ( n33412,p3_eax_reg_0_,n28367 );
   nor U34529 ( n33411,n33414,n33173 );
   nor U34530 ( n33409,n33415,n33416 );
   nor U34531 ( n33416,n30737,n33417 );
   nor U34532 ( n33415,n31926,n28129 );
   not U34533 ( n31926,n33002 );
   nand U34534 ( n33002,n33419,n33420 );
   nor U34535 ( n33420,n33421,n33422 );
   nand U34536 ( n33422,n33423,n33424 );
   nor U34537 ( n33424,n33425,n33426 );
   nor U34538 ( n33426,n33427,n33428 );
   nor U34539 ( n33425,n33429,n33430 );
   nor U34540 ( n33423,n33431,n33432 );
   nor U34541 ( n33432,n33433,n33434 );
   nor U34542 ( n33431,n33435,n33436 );
   nand U34543 ( n33421,n33437,n33438 );
   nor U34544 ( n33438,n33439,n33440 );
   nor U34545 ( n33440,n33441,n33442 );
   nor U34546 ( n33439,n33443,n33444 );
   nor U34547 ( n33437,n33445,n33446 );
   nor U34548 ( n33446,n33447,n33448 );
   nor U34549 ( n33445,n33449,n33450 );
   nor U34550 ( n33419,n33451,n33452 );
   nand U34551 ( n33452,n33453,n33454 );
   nor U34552 ( n33454,n33455,n33456 );
   nor U34553 ( n33456,n33457,n33458 );
   nor U34554 ( n33455,n33459,n33460 );
   nor U34555 ( n33453,n33461,n33462 );
   nor U34556 ( n33462,n33463,n33464 );
   nor U34557 ( n33461,n33465,n33466 );
   nand U34558 ( n33451,n33467,n33468 );
   nor U34559 ( n33468,n33469,n33470 );
   nor U34560 ( n33470,n33471,n33472 );
   nor U34561 ( n33469,n33473,n33474 );
   nor U34562 ( n33467,n33475,n33476 );
   nor U34563 ( n33476,n33477,n33478 );
   nor U34564 ( n33475,n33479,n33480 );
   nor U34565 ( n33482,n33483,n33484 );
   nor U34566 ( n33484,p3_eax_reg_1_,n33485 );
   nand U34567 ( n33485,n28291,p3_eax_reg_0_ );
   and U34568 ( n33483,n33487,p3_eax_reg_1_ );
   nor U34569 ( n33481,n33488,n33489 );
   nor U34570 ( n33489,n30712,n28302 );
   nor U34571 ( n33488,n33003,n28129 );
   not U34572 ( n33003,n31942 );
   nand U34573 ( n31942,n33490,n33491 );
   nor U34574 ( n33491,n33492,n33493 );
   nand U34575 ( n33493,n33494,n33495 );
   nor U34576 ( n33495,n33496,n33497 );
   nor U34577 ( n33497,n33498,n33428 );
   nor U34578 ( n33496,n33499,n33430 );
   nor U34579 ( n33494,n33500,n33501 );
   nor U34580 ( n33501,n33502,n33434 );
   nor U34581 ( n33500,n33503,n33436 );
   nand U34582 ( n33492,n33504,n33505 );
   nor U34583 ( n33505,n33506,n33507 );
   nor U34584 ( n33507,n33508,n33442 );
   nor U34585 ( n33506,n33509,n33444 );
   nor U34586 ( n33504,n33510,n33511 );
   nor U34587 ( n33511,n33512,n33448 );
   nor U34588 ( n33510,n33513,n33450 );
   nor U34589 ( n33490,n33514,n33515 );
   nand U34590 ( n33515,n33516,n33517 );
   nor U34591 ( n33517,n33518,n33519 );
   nor U34592 ( n33519,n33520,n33458 );
   nor U34593 ( n33518,n33521,n33460 );
   nor U34594 ( n33516,n33522,n33523 );
   nor U34595 ( n33523,n33524,n33464 );
   nor U34596 ( n33522,n33525,n33466 );
   nand U34597 ( n33514,n33526,n33527 );
   nor U34598 ( n33527,n33528,n33529 );
   nor U34599 ( n33529,n33530,n33472 );
   nor U34600 ( n33528,n33531,n33474 );
   nor U34601 ( n33526,n33532,n33533 );
   nor U34602 ( n33533,n33534,n33478 );
   nor U34603 ( n33532,n30716,n33480 );
   nor U34604 ( n33536,n33537,n33538 );
   nor U34605 ( n33538,p3_eax_reg_2_,n33539 );
   nand U34606 ( n33539,n33540,n28291 );
   nor U34607 ( n33540,n33168,n33173 );
   nor U34608 ( n33537,n33541,n33163 );
   nor U34609 ( n33541,n33542,n33487 );
   nand U34610 ( n33487,n33414,n33543 );
   nand U34611 ( n33543,n33486,n33173 );
   not U34612 ( n33173,p3_eax_reg_0_ );
   nor U34613 ( n33542,p3_eax_reg_1_,n28366 );
   nor U34614 ( n33535,n33544,n33545 );
   nor U34615 ( n33545,n30701,n28302 );
   nor U34616 ( n33544,n33017,n28128 );
   not U34617 ( n33017,n33040 );
   nand U34618 ( n33040,n33546,n33547 );
   nor U34619 ( n33547,n33548,n33549 );
   nand U34620 ( n33549,n33550,n33551 );
   nor U34621 ( n33551,n33552,n33553 );
   nor U34622 ( n33553,n33554,n33472 );
   nor U34623 ( n33552,n33555,n33474 );
   nor U34624 ( n33550,n33556,n33557 );
   nor U34625 ( n33557,n33558,n33478 );
   nor U34626 ( n33556,n30705,n33480 );
   nand U34627 ( n33548,n33559,n33560 );
   nor U34628 ( n33560,n33561,n33562 );
   nor U34629 ( n33562,n33563,n33458 );
   nor U34630 ( n33561,n33564,n33460 );
   nor U34631 ( n33559,n33565,n33566 );
   nor U34632 ( n33566,n33567,n33464 );
   nor U34633 ( n33565,n33568,n33466 );
   nor U34634 ( n33546,n33569,n33570 );
   nand U34635 ( n33570,n33571,n33572 );
   nor U34636 ( n33572,n33573,n33574 );
   nor U34637 ( n33574,n33575,n33442 );
   nor U34638 ( n33573,n33576,n33444 );
   nor U34639 ( n33571,n33577,n33578 );
   nor U34640 ( n33578,n33579,n33448 );
   nor U34641 ( n33577,n33580,n33450 );
   nand U34642 ( n33569,n33581,n33582 );
   nor U34643 ( n33582,n33583,n33584 );
   nor U34644 ( n33584,n33585,n33428 );
   nor U34645 ( n33583,n33586,n33430 );
   nor U34646 ( n33581,n33587,n33588 );
   nor U34647 ( n33588,n33589,n33434 );
   nor U34648 ( n33587,n33590,n33436 );
   nor U34649 ( n33592,n33593,n33594 );
   nor U34650 ( n33594,p3_eax_reg_3_,n33595 );
   nand U34651 ( n33595,n33596,n28365 );
   and U34652 ( n33593,n33597,p3_eax_reg_3_ );
   nor U34653 ( n33591,n33598,n33599 );
   nor U34654 ( n33599,n30690,n28302 );
   nor U34655 ( n33598,n32995,n28128 );
   not U34656 ( n32995,n33009 );
   nand U34657 ( n33009,n33600,n33601 );
   nor U34658 ( n33601,n33602,n33603 );
   nand U34659 ( n33603,n33604,n33605 );
   nor U34660 ( n33605,n33606,n33607 );
   nor U34661 ( n33607,n33608,n33428 );
   nor U34662 ( n33606,n33609,n33430 );
   nor U34663 ( n33604,n33610,n33611 );
   nor U34664 ( n33611,n33612,n33434 );
   nor U34665 ( n33610,n33613,n33436 );
   nand U34666 ( n33602,n33614,n33615 );
   nor U34667 ( n33615,n33616,n33617 );
   nor U34668 ( n33617,n33618,n33442 );
   nor U34669 ( n33616,n33619,n33444 );
   nor U34670 ( n33614,n33620,n33621 );
   nor U34671 ( n33621,n33622,n33448 );
   nor U34672 ( n33620,n33623,n33450 );
   nor U34673 ( n33600,n33624,n33625 );
   nand U34674 ( n33625,n33626,n33627 );
   nor U34675 ( n33627,n33628,n33629 );
   nor U34676 ( n33629,n33630,n33458 );
   nor U34677 ( n33628,n33631,n33460 );
   nor U34678 ( n33626,n33632,n33633 );
   nor U34679 ( n33633,n33634,n33464 );
   nor U34680 ( n33632,n33635,n33466 );
   nand U34681 ( n33624,n33636,n33637 );
   nor U34682 ( n33637,n33638,n33639 );
   nor U34683 ( n33639,n33640,n33472 );
   nor U34684 ( n33638,n33641,n33474 );
   nor U34685 ( n33636,n33642,n33643 );
   nor U34686 ( n33643,n33644,n33478 );
   nor U34687 ( n33642,n30694,n33480 );
   nor U34688 ( n33646,n33647,n33648 );
   nor U34689 ( n33648,p3_eax_reg_4_,n33649 );
   nand U34690 ( n33649,n33650,n33596 );
   nor U34691 ( n33650,n33158,n28366 );
   nor U34692 ( n33647,n33651,n33153 );
   nor U34693 ( n33651,n33652,n33597 );
   nand U34694 ( n33597,n33414,n33653 );
   nand U34695 ( n33653,n28291,n33654 );
   nor U34696 ( n33652,p3_eax_reg_3_,n28366 );
   nor U34697 ( n33645,n33655,n33656 );
   nor U34698 ( n33656,n30680,n33417 );
   nor U34699 ( n33655,n33007,n33418 );
   and U34700 ( n33007,n33657,n33658 );
   nor U34701 ( n33658,n33659,n33660 );
   nand U34702 ( n33660,n33661,n33662 );
   nor U34703 ( n33662,n33663,n33664 );
   nor U34704 ( n33664,n33665,n33472 );
   nor U34705 ( n33663,n33666,n33474 );
   nor U34706 ( n33661,n33667,n33668 );
   nor U34707 ( n33668,n33669,n33478 );
   nor U34708 ( n33667,n30683,n33480 );
   nand U34709 ( n33659,n33670,n33671 );
   nor U34710 ( n33671,n33672,n33673 );
   nor U34711 ( n33673,n33674,n33458 );
   nor U34712 ( n33672,n33675,n33460 );
   nor U34713 ( n33670,n33676,n33677 );
   nor U34714 ( n33677,n33678,n33464 );
   nor U34715 ( n33676,n33679,n33466 );
   nor U34716 ( n33657,n33680,n33681 );
   nand U34717 ( n33681,n33682,n33683 );
   nor U34718 ( n33683,n33684,n33685 );
   nor U34719 ( n33685,n33686,n33442 );
   nor U34720 ( n33684,n33687,n33444 );
   nor U34721 ( n33682,n33688,n33689 );
   nor U34722 ( n33689,n33690,n33448 );
   nor U34723 ( n33688,n33691,n33450 );
   nand U34724 ( n33680,n33692,n33693 );
   nor U34725 ( n33693,n33694,n33695 );
   nor U34726 ( n33695,n33696,n33428 );
   nor U34727 ( n33694,n33697,n33430 );
   nor U34728 ( n33692,n33698,n33699 );
   nor U34729 ( n33699,n33700,n33434 );
   nor U34730 ( n33698,n33701,n33436 );
   nor U34731 ( n33703,n33704,n33705 );
   nor U34732 ( n33705,p3_eax_reg_5_,n33706 );
   nand U34733 ( n33706,n33707,n28291 );
   and U34734 ( n33704,n33708,p3_eax_reg_5_ );
   nor U34735 ( n33702,n33709,n33710 );
   nor U34736 ( n33710,n30669,n33417 );
   nor U34737 ( n33709,n32967,n28129 );
   and U34738 ( n32967,n33711,n33712 );
   nor U34739 ( n33712,n33713,n33714 );
   nand U34740 ( n33714,n33715,n33716 );
   nor U34741 ( n33716,n33717,n33718 );
   nor U34742 ( n33718,n33719,n33472 );
   nor U34743 ( n33717,n33720,n33474 );
   nor U34744 ( n33715,n33721,n33722 );
   nor U34745 ( n33722,n33723,n33478 );
   nor U34746 ( n33721,n30673,n33480 );
   nand U34747 ( n33713,n33724,n33725 );
   nor U34748 ( n33725,n33726,n33727 );
   nor U34749 ( n33727,n33728,n33458 );
   nor U34750 ( n33726,n33729,n33460 );
   nor U34751 ( n33724,n33730,n33731 );
   nor U34752 ( n33731,n33732,n33464 );
   nor U34753 ( n33730,n33733,n33466 );
   nor U34754 ( n33711,n33734,n33735 );
   nand U34755 ( n33735,n33736,n33737 );
   nor U34756 ( n33737,n33738,n33739 );
   nor U34757 ( n33739,n33740,n33442 );
   nor U34758 ( n33738,n33741,n33444 );
   nor U34759 ( n33736,n33742,n33743 );
   nor U34760 ( n33743,n33744,n33448 );
   nor U34761 ( n33742,n33745,n33450 );
   nand U34762 ( n33734,n33746,n33747 );
   nor U34763 ( n33747,n33748,n33749 );
   nor U34764 ( n33749,n33750,n33428 );
   nor U34765 ( n33748,n33751,n33430 );
   nor U34766 ( n33746,n33752,n33753 );
   nor U34767 ( n33753,n33754,n33434 );
   nor U34768 ( n33752,n33755,n33436 );
   nor U34769 ( n33757,n33758,n33759 );
   nor U34770 ( n33759,p3_eax_reg_6_,n33760 );
   nand U34771 ( n33760,n33761,n33707 );
   nor U34772 ( n33761,n33148,n28367 );
   nor U34773 ( n33758,n33762,n33143 );
   nor U34774 ( n33762,n33763,n33708 );
   nand U34775 ( n33708,n33414,n33764 );
   nand U34776 ( n33764,n28365,n33765 );
   nor U34777 ( n33763,p3_eax_reg_5_,n28366 );
   nor U34778 ( n33756,n33766,n33767 );
   nor U34779 ( n33767,n30658,n33417 );
   nor U34780 ( n33766,n33010,n28129 );
   not U34781 ( n33010,n33014 );
   nand U34782 ( n33014,n33768,n33769 );
   nor U34783 ( n33769,n33770,n33771 );
   nand U34784 ( n33771,n33772,n33773 );
   nor U34785 ( n33773,n33774,n33775 );
   nor U34786 ( n33775,n33776,n33428 );
   nor U34787 ( n33774,n33777,n33430 );
   nor U34788 ( n33772,n33778,n33779 );
   nor U34789 ( n33779,n33780,n33434 );
   nor U34790 ( n33778,n33781,n33436 );
   nand U34791 ( n33770,n33782,n33783 );
   nor U34792 ( n33783,n33784,n33785 );
   nor U34793 ( n33785,n33786,n33442 );
   nor U34794 ( n33784,n33787,n33444 );
   nor U34795 ( n33782,n33788,n33789 );
   nor U34796 ( n33789,n33790,n33448 );
   nor U34797 ( n33788,n33791,n33450 );
   nor U34798 ( n33768,n33792,n33793 );
   nand U34799 ( n33793,n33794,n33795 );
   nor U34800 ( n33795,n33796,n33797 );
   nor U34801 ( n33797,n33798,n33458 );
   nor U34802 ( n33796,n33799,n33460 );
   nor U34803 ( n33794,n33800,n33801 );
   nor U34804 ( n33801,n33802,n33464 );
   nor U34805 ( n33800,n33803,n33466 );
   nand U34806 ( n33792,n33804,n33805 );
   nor U34807 ( n33805,n33806,n33807 );
   nor U34808 ( n33807,n33808,n33472 );
   nor U34809 ( n33806,n33809,n33474 );
   nor U34810 ( n33804,n33810,n33811 );
   nor U34811 ( n33811,n33812,n33478 );
   nor U34812 ( n33810,n30662,n33480 );
   nor U34813 ( n33814,n33815,n33816 );
   nor U34814 ( n33816,p3_eax_reg_7_,n33817 );
   nand U34815 ( n33817,n33818,n33486 );
   and U34816 ( n33815,n33819,p3_eax_reg_7_ );
   nor U34817 ( n33813,n33820,n33821 );
   nor U34818 ( n33821,n30643,n33417 );
   nor U34819 ( n33820,n31694,n33418 );
   not U34820 ( n31694,n31915 );
   nand U34821 ( n31915,n33822,n33823 );
   nor U34822 ( n33823,n33824,n33825 );
   nand U34823 ( n33825,n33826,n33827 );
   nor U34824 ( n33827,n33828,n33829 );
   nor U34825 ( n33829,n33830,n33428 );
   nand U34826 ( n33428,n33831,n33832 );
   nor U34827 ( n33828,n33833,n33430 );
   nand U34828 ( n33430,n33831,n33834 );
   nor U34829 ( n33826,n33835,n33836 );
   nor U34830 ( n33836,n33837,n33434 );
   nand U34831 ( n33434,n33831,n33838 );
   nor U34832 ( n33835,n33839,n33436 );
   nand U34833 ( n33436,n33832,n33840 );
   nand U34834 ( n33824,n33841,n33842 );
   nor U34835 ( n33842,n33843,n33844 );
   nor U34836 ( n33844,n33845,n33442 );
   nand U34837 ( n33442,n33834,n33840 );
   nor U34838 ( n33843,n33846,n33444 );
   nand U34839 ( n33444,n33838,n33840 );
   nor U34840 ( n33841,n33847,n33848 );
   nor U34841 ( n33848,n33849,n33448 );
   nand U34842 ( n33448,n33832,n33850 );
   nor U34843 ( n33847,n33851,n33450 );
   nand U34844 ( n33450,n33850,n33834 );
   nor U34845 ( n33822,n33852,n33853 );
   nand U34846 ( n33853,n33854,n33855 );
   nor U34847 ( n33855,n33856,n33857 );
   nor U34848 ( n33857,n33858,n33458 );
   nand U34849 ( n33458,n33850,n33838 );
   nor U34850 ( n33856,n33859,n33460 );
   nand U34851 ( n33460,n33860,n33832 );
   nor U34852 ( n33854,n33861,n33862 );
   nor U34853 ( n33862,n33863,n33464 );
   nand U34854 ( n33464,n33860,n33834 );
   nor U34855 ( n33861,n33864,n33466 );
   nand U34856 ( n33466,n33860,n33838 );
   nand U34857 ( n33852,n33865,n33866 );
   nor U34858 ( n33866,n33867,n33868 );
   nor U34859 ( n33868,n33869,n33472 );
   nand U34860 ( n33472,n33870,n33840 );
   nor U34861 ( n33840,n28874,n33871 );
   nor U34862 ( n33867,n33872,n33474 );
   nand U34863 ( n33474,n33870,n33850 );
   nor U34864 ( n33850,n28862,n33873 );
   nor U34865 ( n33865,n33874,n33875 );
   nor U34866 ( n33875,n33876,n33478 );
   nand U34867 ( n33478,n33860,n33870 );
   nor U34868 ( n33860,n33871,n33873 );
   not U34869 ( n33873,n28874 );
   nor U34870 ( n33874,n30650,n33480 );
   nand U34871 ( n33480,n33870,n33831 );
   nor U34872 ( n33831,n28874,n28862 );
   nand U34873 ( n28874,n33877,n33878 );
   nand U34874 ( n33878,p3_instqueuerd_addr_reg_3_,n29274 );
   nor U34875 ( n33880,n33881,n33882 );
   nor U34876 ( n33882,p3_eax_reg_8_,n33883 );
   nand U34877 ( n33883,n33884,n33818 );
   nor U34878 ( n33884,n33138,n28367 );
   nor U34879 ( n33881,n33885,n33133 );
   nor U34880 ( n33885,n33886,n33819 );
   nand U34881 ( n33819,n33414,n33887 );
   nand U34882 ( n33887,n28291,n33888 );
   nor U34883 ( n33886,p3_eax_reg_7_,n28367 );
   nor U34884 ( n33879,n33889,n33890 );
   nor U34885 ( n33890,n33208,n33417 );
   nor U34886 ( n33889,n33891,n28128 );
   not U34887 ( n33891,n33892 );
   nor U34888 ( n33894,n33895,n33896 );
   nor U34889 ( n33896,p3_eax_reg_9_,n33897 );
   nand U34890 ( n33897,n33898,n28291 );
   and U34891 ( n33895,n33899,p3_eax_reg_9_ );
   nor U34892 ( n33893,n33900,n33901 );
   nor U34893 ( n33901,n33203,n33417 );
   nor U34894 ( n33900,n33902,n28129 );
   not U34895 ( n33902,n33903 );
   nor U34896 ( n33905,n33906,n33907 );
   nor U34897 ( n33907,p3_eax_reg_10_,n33908 );
   nand U34898 ( n33908,n33909,n33898 );
   nor U34899 ( n33909,n33128,n28366 );
   nor U34900 ( n33906,n33910,n33123 );
   nor U34901 ( n33910,n33911,n33899 );
   nand U34902 ( n33899,n33414,n33912 );
   nand U34903 ( n33912,n28365,n33913 );
   nor U34904 ( n33911,p3_eax_reg_9_,n33413 );
   nor U34905 ( n33904,n33914,n33915 );
   nor U34906 ( n33915,n33198,n33417 );
   nor U34907 ( n33914,n33916,n33418 );
   not U34908 ( n33916,n33917 );
   nor U34909 ( n33919,n33920,n33921 );
   nor U34910 ( n33921,p3_eax_reg_11_,n33922 );
   nand U34911 ( n33922,n33923,n33486 );
   and U34912 ( n33920,n33924,p3_eax_reg_11_ );
   nor U34913 ( n33918,n33925,n33926 );
   nor U34914 ( n33926,n33193,n33417 );
   nor U34915 ( n33925,n33927,n28128 );
   not U34916 ( n33927,n33928 );
   nor U34917 ( n33930,n33931,n33932 );
   nor U34918 ( n33932,p3_eax_reg_12_,n33933 );
   nand U34919 ( n33933,n33934,n33923 );
   nor U34920 ( n33934,n33118,n28367 );
   nor U34921 ( n33931,n33935,n33113 );
   nor U34922 ( n33935,n33936,n33924 );
   nand U34923 ( n33924,n33414,n33937 );
   nand U34924 ( n33937,n28291,n33938 );
   nor U34925 ( n33936,p3_eax_reg_11_,n28366 );
   nor U34926 ( n33929,n33939,n33940 );
   nor U34927 ( n33940,n33188,n33417 );
   nor U34928 ( n33939,n33941,n28129 );
   not U34929 ( n33941,n33942 );
   nor U34930 ( n33944,n33945,n33946 );
   nor U34931 ( n33946,p3_eax_reg_13_,n33947 );
   nand U34932 ( n33947,n33948,n33486 );
   and U34933 ( n33945,n33949,p3_eax_reg_13_ );
   nor U34934 ( n33943,n33950,n33951 );
   nor U34935 ( n33951,n33183,n33417 );
   nor U34936 ( n33950,n33952,n28128 );
   not U34937 ( n33952,n33953 );
   nor U34938 ( n33955,n33956,n33957 );
   nor U34939 ( n33957,p3_eax_reg_14_,n33958 );
   nand U34940 ( n33958,n33959,n33948 );
   nor U34941 ( n33959,n33108,n33413 );
   nor U34942 ( n33956,n33960,n33103 );
   nor U34943 ( n33960,n33961,n33949 );
   nand U34944 ( n33949,n33414,n33962 );
   nand U34945 ( n33962,n33486,n33963 );
   nor U34946 ( n33961,p3_eax_reg_13_,n28366 );
   nor U34947 ( n33954,n33964,n33965 );
   nor U34948 ( n33965,n33178,n28302 );
   nor U34949 ( n33964,n33966,n33418 );
   not U34950 ( n33966,n33967 );
   nor U34951 ( n33969,n33970,n33971 );
   nor U34952 ( n33971,p3_eax_reg_15_,n33972 );
   nand U34953 ( n33972,n33973,n28291 );
   nor U34954 ( n33970,n33974,n33096 );
   nor U34955 ( n33968,n33975,n33976 );
   nor U34956 ( n33976,n33097,n33417 );
   nand U34957 ( n33417,n31859,n27893 );
   nor U34958 ( n31859,n31784,n31809 );
   not U34959 ( n33097,buf2_reg_15_ );
   nor U34960 ( n33975,n33977,n28128 );
   not U34961 ( n33977,n33978 );
   nor U34962 ( n33980,n33981,n33982 );
   nor U34963 ( n33982,n30737,n33983 );
   nor U34964 ( n33981,n33984,n33418 );
   not U34965 ( n33984,n33985 );
   nor U34966 ( n33979,n33986,n33987 );
   nand U34967 ( n33987,n33988,n33989 );
   nand U34968 ( n33989,p3_eax_reg_16_,n33990 );
   nand U34969 ( n33990,n33974,n33991 );
   nand U34970 ( n33991,n28365,n33096 );
   and U34971 ( n33974,n33414,n33992 );
   nand U34972 ( n33992,n33486,n33993 );
   nand U34973 ( n33988,n33994,n33240 );
   nor U34974 ( n33994,n33993,n33995 );
   nand U34975 ( n33995,n28291,p3_eax_reg_15_ );
   and U34976 ( n33986,buf2_reg_16_,n33996 );
   nor U34977 ( n33998,n33999,n34000 );
   nor U34978 ( n34000,n30712,n28233 );
   nor U34979 ( n33999,n34001,n33418 );
   not U34980 ( n34001,n34002 );
   nor U34981 ( n33997,n34003,n34004 );
   nand U34982 ( n34004,n34005,n34006 );
   nand U34983 ( n34006,p3_eax_reg_17_,n34007 );
   nand U34984 ( n34005,n34008,n33236 );
   nor U34985 ( n34008,n28366,n34009 );
   and U34986 ( n34003,buf2_reg_17_,n33996 );
   nor U34987 ( n34011,n34012,n34013 );
   nor U34988 ( n34013,n30701,n28233 );
   nor U34989 ( n34012,n34014,n28129 );
   not U34990 ( n34014,n34015 );
   nor U34991 ( n34010,n34016,n34017 );
   nand U34992 ( n34017,n34018,n34019 );
   nand U34993 ( n34019,p3_eax_reg_18_,n34020 );
   nand U34994 ( n34020,n34021,n34022 );
   nand U34995 ( n34022,n28365,n33236 );
   not U34996 ( n33236,p3_eax_reg_17_ );
   not U34997 ( n34021,n34007 );
   nand U34998 ( n34007,n27893,n34023 );
   nand U34999 ( n34023,n33486,n34009 );
   nand U35000 ( n34018,n34024,n33232 );
   not U35001 ( n33232,p3_eax_reg_18_ );
   nor U35002 ( n34024,n34009,n34025 );
   nand U35003 ( n34025,n28291,p3_eax_reg_17_ );
   and U35004 ( n34016,buf2_reg_18_,n33996 );
   nor U35005 ( n34027,n34028,n34029 );
   nor U35006 ( n34029,n30690,n28233 );
   nor U35007 ( n34028,n34030,n28128 );
   not U35008 ( n34030,n34031 );
   nor U35009 ( n34026,n34032,n34033 );
   nand U35010 ( n34033,n34034,n34035 );
   nand U35011 ( n34035,p3_eax_reg_19_,n34036 );
   nand U35012 ( n34034,n34037,n33228 );
   nor U35013 ( n34037,n33413,n34038 );
   and U35014 ( n34032,buf2_reg_19_,n33996 );
   nor U35015 ( n34040,n34041,n34042 );
   nor U35016 ( n34042,n30680,n33983 );
   nor U35017 ( n34041,n34043,n28129 );
   not U35018 ( n34043,n34044 );
   nor U35019 ( n34039,n34045,n34046 );
   nand U35020 ( n34046,n34047,n34048 );
   nand U35021 ( n34048,p3_eax_reg_20_,n34049 );
   nand U35022 ( n34049,n34050,n34051 );
   nand U35023 ( n34051,n33486,n33228 );
   not U35024 ( n34050,n34036 );
   nand U35025 ( n34036,n27893,n34052 );
   nand U35026 ( n34052,n33486,n34038 );
   nand U35027 ( n34047,n34053,n33224 );
   nor U35028 ( n34053,n34038,n34054 );
   nand U35029 ( n34054,n28291,p3_eax_reg_19_ );
   not U35030 ( n34038,n34055 );
   and U35031 ( n34045,buf2_reg_20_,n33996 );
   nor U35032 ( n34057,n34058,n34059 );
   nor U35033 ( n34059,n30669,n33983 );
   nor U35034 ( n34058,n34060,n33418 );
   not U35035 ( n34060,n34061 );
   nor U35036 ( n34056,n34062,n34063 );
   nand U35037 ( n34063,n34064,n34065 );
   nand U35038 ( n34065,p3_eax_reg_21_,n34066 );
   nand U35039 ( n34064,n34067,n33220 );
   nor U35040 ( n34067,n28367,n34068 );
   and U35041 ( n34062,buf2_reg_21_,n33996 );
   nor U35042 ( n34070,n34071,n34072 );
   nor U35043 ( n34072,n30658,n33983 );
   nor U35044 ( n34071,n34073,n28129 );
   not U35045 ( n34073,n34074 );
   nor U35046 ( n34069,n34075,n34076 );
   nand U35047 ( n34076,n34077,n34078 );
   nand U35048 ( n34078,p3_eax_reg_22_,n34079 );
   nand U35049 ( n34079,n34080,n34081 );
   nand U35050 ( n34081,n33486,n33220 );
   not U35051 ( n33220,p3_eax_reg_21_ );
   not U35052 ( n34080,n34066 );
   nand U35053 ( n34066,n33414,n34082 );
   nand U35054 ( n34082,n28291,n34068 );
   nand U35055 ( n34077,n34083,n33216 );
   not U35056 ( n33216,p3_eax_reg_22_ );
   nor U35057 ( n34083,n34068,n34084 );
   nand U35058 ( n34084,n28365,p3_eax_reg_21_ );
   and U35059 ( n34075,buf2_reg_22_,n33996 );
   nor U35060 ( n34086,n34087,n34088 );
   nor U35061 ( n34088,n30643,n33983 );
   nor U35062 ( n34087,n34089,n28128 );
   not U35063 ( n34089,n34090 );
   nor U35064 ( n34085,n34091,n34092 );
   nand U35065 ( n34092,n34093,n34094 );
   nand U35066 ( n34094,p3_eax_reg_23_,n34095 );
   nand U35067 ( n34093,n34096,n33212 );
   nor U35068 ( n34096,n28366,n34097 );
   and U35069 ( n34091,buf2_reg_23_,n33996 );
   nor U35070 ( n34099,n34100,n34101 );
   nor U35071 ( n34101,n33208,n33983 );
   nor U35072 ( n34100,n28128,n34102 );
   nor U35073 ( n34098,n34103,n34104 );
   nand U35074 ( n34104,n34105,n34106 );
   nand U35075 ( n34106,p3_eax_reg_24_,n34107 );
   nand U35076 ( n34107,n34108,n34109 );
   nand U35077 ( n34109,n33486,n33212 );
   not U35078 ( n34108,n34095 );
   nand U35079 ( n34095,n33414,n34110 );
   nand U35080 ( n34110,n28291,n34097 );
   nand U35081 ( n34105,n34111,n33207 );
   nor U35082 ( n34111,n34097,n34112 );
   nand U35083 ( n34112,n33486,p3_eax_reg_23_ );
   not U35084 ( n34097,n34113 );
   and U35085 ( n34103,buf2_reg_24_,n33996 );
   nor U35086 ( n34115,n34116,n34117 );
   nor U35087 ( n34117,n33203,n33983 );
   nor U35088 ( n34116,n33418,n34118 );
   or U35089 ( n34118,n34119,n34120 );
   nor U35090 ( n34114,n34121,n34122 );
   nand U35091 ( n34122,n34123,n34124 );
   nand U35092 ( n34124,p3_eax_reg_25_,n34125 );
   nand U35093 ( n34123,n34126,n33202 );
   nor U35094 ( n34126,n28367,n34127 );
   and U35095 ( n34121,buf2_reg_25_,n33996 );
   nor U35096 ( n34129,n34130,n34131 );
   nor U35097 ( n34131,n33198,n33983 );
   nor U35098 ( n34130,n28129,n34132 );
   nor U35099 ( n34128,n34133,n34134 );
   nand U35100 ( n34134,n34135,n34136 );
   nand U35101 ( n34136,p3_eax_reg_26_,n34137 );
   nand U35102 ( n34137,n34138,n34139 );
   nand U35103 ( n34139,n28365,n33202 );
   not U35104 ( n33202,p3_eax_reg_25_ );
   not U35105 ( n34138,n34125 );
   nand U35106 ( n34125,n33414,n34140 );
   nand U35107 ( n34140,n33486,n34127 );
   nand U35108 ( n34135,n34141,n33197 );
   not U35109 ( n33197,p3_eax_reg_26_ );
   nor U35110 ( n34141,n34127,n34142 );
   nand U35111 ( n34142,n33486,p3_eax_reg_25_ );
   and U35112 ( n34133,buf2_reg_26_,n33996 );
   nor U35113 ( n34144,n34145,n34146 );
   nor U35114 ( n34146,n33193,n33983 );
   nor U35115 ( n34145,n28128,n34147 );
   nand U35116 ( n34147,n34148,n34149 );
   nor U35117 ( n34143,n34150,n34151 );
   nand U35118 ( n34151,n34152,n34153 );
   nand U35119 ( n34153,p3_eax_reg_27_,n34154 );
   nand U35120 ( n34152,n34155,n33192 );
   nor U35121 ( n34155,n28366,n34156 );
   and U35122 ( n34150,buf2_reg_27_,n33996 );
   nor U35123 ( n34158,n34159,n34160 );
   nor U35124 ( n34160,n33188,n33983 );
   nor U35125 ( n34159,n28129,n34161 );
   nor U35126 ( n34157,n34162,n34163 );
   nand U35127 ( n34163,n34164,n34165 );
   or U35128 ( n34165,n33187,n34166 );
   nand U35129 ( n34164,n34167,n33187 );
   nor U35130 ( n34167,n34156,n34168 );
   nand U35131 ( n34168,n28365,p3_eax_reg_27_ );
   and U35132 ( n34162,buf2_reg_28_,n33996 );
   nor U35133 ( n34170,n34171,n34172 );
   nand U35134 ( n34172,n34173,n34174 );
   nand U35135 ( n34174,p3_eax_reg_29_,n34175 );
   nand U35136 ( n34175,n34166,n34176 );
   nand U35137 ( n34176,n28365,n33187 );
   nor U35138 ( n34166,n34154,n34177 );
   nor U35139 ( n34177,n28367,p3_eax_reg_27_ );
   nand U35140 ( n34154,n33414,n34178 );
   nand U35141 ( n34178,n28291,n34156 );
   not U35142 ( n34156,n34179 );
   not U35143 ( n33486,n33413 );
   nand U35144 ( n34173,n34180,n34181 );
   nor U35145 ( n34171,n33418,n34182 );
   not U35146 ( n34182,n34183 );
   nor U35147 ( n34169,n34184,n34185 );
   and U35148 ( n34185,buf2_reg_29_,n33996 );
   nor U35149 ( n34184,n33183,n33983 );
   nor U35150 ( n34187,n34188,n34189 );
   nor U35151 ( n34189,n33178,n33983 );
   nand U35152 ( n33983,n34190,n27893 );
   nor U35153 ( n34190,n31809,n30670 );
   nor U35154 ( n34188,n28128,n34191 );
   not U35155 ( n34191,n34192 );
   nand U35156 ( n33418,n33414,n31784 );
   not U35157 ( n31784,n31886 );
   nor U35158 ( n34186,n34193,n34194 );
   nand U35159 ( n34194,n34195,n34196 );
   nand U35160 ( n34196,p3_eax_reg_30_,n34197 );
   nand U35161 ( n34195,n34198,n33177 );
   not U35162 ( n33177,p3_eax_reg_30_ );
   and U35163 ( n34193,buf2_reg_30_,n33996 );
   nand U35164 ( n34200,n33996,buf2_reg_31_ );
   and U35165 ( n33996,n34201,n27893 );
   nor U35166 ( n34201,n31809,n34202 );
   nor U35167 ( n34199,n34203,n34204 );
   nor U35168 ( n34204,p3_eax_reg_31_,n34205 );
   nand U35169 ( n34205,n34198,p3_eax_reg_30_ );
   and U35170 ( n34198,n34206,n34181 );
   nor U35171 ( n34206,n33182,n28367 );
   not U35172 ( n33182,p3_eax_reg_29_ );
   nor U35173 ( n34203,n34207,n34208 );
   not U35174 ( n34208,p3_eax_reg_31_ );
   nor U35175 ( n34207,n34209,n34197 );
   nand U35176 ( n34197,n34210,n27893 );
   nor U35177 ( n34210,n34180,n34211 );
   nor U35178 ( n34211,n34181,n33413 );
   and U35179 ( n34181,n34212,n34179 );
   nor U35180 ( n34179,n34213,n34127 );
   nand U35181 ( n34127,n34214,n34113 );
   nor U35182 ( n34113,n34215,n34068 );
   nand U35183 ( n34068,n34216,n34055 );
   nor U35184 ( n34055,n34217,n34009 );
   nand U35185 ( n34009,n34218,n33973 );
   not U35186 ( n33973,n33993 );
   nand U35187 ( n33993,n34219,n33948 );
   not U35188 ( n33948,n33963 );
   nand U35189 ( n33963,n34220,n33923 );
   not U35190 ( n33923,n33938 );
   nand U35191 ( n33938,n34221,n33898 );
   not U35192 ( n33898,n33913 );
   nand U35193 ( n33913,n34222,n33818 );
   not U35194 ( n33818,n33888 );
   nand U35195 ( n33888,n34223,n33707 );
   not U35196 ( n33707,n33765 );
   nand U35197 ( n33765,n34224,n33596 );
   not U35198 ( n33596,n33654 );
   nand U35199 ( n33654,n34225,p3_eax_reg_0_ );
   nor U35200 ( n34225,n33163,n33168 );
   not U35201 ( n33168,p3_eax_reg_1_ );
   not U35202 ( n33163,p3_eax_reg_2_ );
   nor U35203 ( n34224,n33153,n33158 );
   not U35204 ( n33158,p3_eax_reg_3_ );
   not U35205 ( n33153,p3_eax_reg_4_ );
   nor U35206 ( n34223,n33143,n33148 );
   not U35207 ( n33148,p3_eax_reg_5_ );
   not U35208 ( n33143,p3_eax_reg_6_ );
   nor U35209 ( n34222,n33133,n33138 );
   not U35210 ( n33138,p3_eax_reg_7_ );
   not U35211 ( n33133,p3_eax_reg_8_ );
   nor U35212 ( n34221,n33123,n33128 );
   not U35213 ( n33128,p3_eax_reg_9_ );
   not U35214 ( n33123,p3_eax_reg_10_ );
   nor U35215 ( n34220,n33113,n33118 );
   not U35216 ( n33118,p3_eax_reg_11_ );
   not U35217 ( n33113,p3_eax_reg_12_ );
   nor U35218 ( n34219,n33103,n33108 );
   not U35219 ( n33108,p3_eax_reg_13_ );
   not U35220 ( n33103,p3_eax_reg_14_ );
   nor U35221 ( n34218,n33096,n33240 );
   not U35222 ( n33240,p3_eax_reg_16_ );
   not U35223 ( n33096,p3_eax_reg_15_ );
   nand U35224 ( n34217,p3_eax_reg_18_,p3_eax_reg_17_ );
   nor U35225 ( n34216,n33224,n33228 );
   not U35226 ( n33228,p3_eax_reg_19_ );
   not U35227 ( n33224,p3_eax_reg_20_ );
   nand U35228 ( n34215,p3_eax_reg_22_,p3_eax_reg_21_ );
   nor U35229 ( n34214,n33207,n33212 );
   not U35230 ( n33212,p3_eax_reg_23_ );
   not U35231 ( n33207,p3_eax_reg_24_ );
   nand U35232 ( n34213,p3_eax_reg_26_,p3_eax_reg_25_ );
   nor U35233 ( n34212,n33187,n33192 );
   not U35234 ( n33192,p3_eax_reg_27_ );
   not U35235 ( n33187,p3_eax_reg_28_ );
   nor U35236 ( n34180,n33413,p3_eax_reg_29_ );
   nor U35237 ( n34209,p3_eax_reg_30_,n33413 );
   nand U35238 ( n33413,n33414,n31809 );
   and U35239 ( n33414,n31747,n34226 );
   or U35240 ( n34226,n29377,n29334 );
   nor U35241 ( n29334,n29301,n31810 );
   nand U35242 ( n29377,n34227,n34228 );
   nand U35243 ( n34228,n34229,n29224 );
   nor U35244 ( n34229,n34230,n28801 );
   nand U35245 ( n34227,n31759,n29221 );
   nor U35246 ( n29221,n29247,n31810 );
   not U35247 ( n31810,n29315 );
   nand U35248 ( n34232,n34233,p3_instqueue_reg_0__0_ );
   nor U35249 ( n34231,n34234,n34235 );
   nor U35250 ( n34235,n34236,n34237 );
   nor U35251 ( n34234,p3_ebx_reg_0_,n28172 );
   nand U35252 ( n34240,p3_ebx_reg_1_,n34241 );
   nor U35253 ( n34239,n34242,n34243 );
   and U35254 ( n34243,p3_instqueue_reg_0__1_,n28283 );
   and U35255 ( n34242,n34244,n28170 );
   nand U35256 ( n34247,n34233,p3_instqueue_reg_0__2_ );
   nor U35257 ( n34246,n34248,n34249 );
   nor U35258 ( n34249,p3_ebx_reg_2_,n34250 );
   nand U35259 ( n34250,n34251,n28170 );
   nor U35260 ( n34248,n34252,n34253 );
   nor U35261 ( n34252,n34254,n34241 );
   nor U35262 ( n34254,n34251,n28173 );
   nand U35263 ( n34256,n34233,p3_instqueue_reg_0__3_ );
   nor U35264 ( n34255,n34257,n34258 );
   nor U35265 ( n34258,p3_ebx_reg_3_,n34259 );
   or U35266 ( n34259,n34260,n28172 );
   and U35267 ( n34257,n34261,p3_ebx_reg_3_ );
   nand U35268 ( n34263,n34233,p3_instqueue_reg_0__4_ );
   nor U35269 ( n34262,n34264,n34265 );
   nor U35270 ( n34265,p3_ebx_reg_4_,n34266 );
   nand U35271 ( n34266,n34267,p3_ebx_reg_3_ );
   nor U35272 ( n34267,n28171,n34260 );
   nor U35273 ( n34264,n34268,n34269 );
   nor U35274 ( n34268,n34270,n34261 );
   nand U35275 ( n34261,n34236,n34271 );
   nand U35276 ( n34271,n34245,n34260 );
   nor U35277 ( n34270,p3_ebx_reg_3_,n28171 );
   nand U35278 ( n34273,n34233,p3_instqueue_reg_0__5_ );
   nor U35279 ( n34272,n34274,n34275 );
   nor U35280 ( n34275,p3_ebx_reg_5_,n34276 );
   or U35281 ( n34276,n34277,n28172 );
   and U35282 ( n34274,n34278,p3_ebx_reg_5_ );
   nand U35283 ( n34280,n34233,p3_instqueue_reg_0__6_ );
   nor U35284 ( n34279,n34281,n34282 );
   nor U35285 ( n34282,p3_ebx_reg_6_,n34283 );
   nand U35286 ( n34283,n34284,p3_ebx_reg_5_ );
   nor U35287 ( n34284,n28173,n34277 );
   nor U35288 ( n34281,n34285,n34286 );
   nor U35289 ( n34285,n34287,n34278 );
   nand U35290 ( n34278,n34236,n34288 );
   nand U35291 ( n34288,n34245,n34277 );
   nor U35292 ( n34287,p3_ebx_reg_5_,n28172 );
   nand U35293 ( n34290,n34233,p3_instqueue_reg_0__7_ );
   nor U35294 ( n34289,n34291,n34292 );
   nor U35295 ( n34292,p3_ebx_reg_7_,n34293 );
   or U35296 ( n34293,n34294,n28171 );
   and U35297 ( n34291,n34295,p3_ebx_reg_7_ );
   nand U35298 ( n34297,n34233,n33892 );
   nand U35299 ( n33892,n34298,n34299 );
   nor U35300 ( n34299,n34300,n34301 );
   nand U35301 ( n34301,n34302,n34303 );
   nor U35302 ( n34303,n34304,n34305 );
   nor U35303 ( n34305,n33463,n34306 );
   nor U35304 ( n34304,n33459,n34307 );
   nor U35305 ( n34302,n34308,n34309 );
   nor U35306 ( n34309,n33477,n34310 );
   nor U35307 ( n34308,n33449,n34311 );
   nand U35308 ( n34300,n34312,n34313 );
   nor U35309 ( n34313,n34314,n34315 );
   nor U35310 ( n34315,n33447,n34316 );
   nor U35311 ( n34314,n33473,n34317 );
   nor U35312 ( n34312,n34318,n34319 );
   nor U35313 ( n34319,n33441,n34320 );
   nor U35314 ( n34318,n33435,n34321 );
   nor U35315 ( n34298,n34322,n34323 );
   nand U35316 ( n34323,n34324,n34325 );
   nor U35317 ( n34325,n34326,n34327 );
   nor U35318 ( n34327,n33471,n34328 );
   nor U35319 ( n34326,n33429,n34329 );
   nor U35320 ( n34324,n34330,n34331 );
   nor U35321 ( n34331,n33427,n34332 );
   nor U35322 ( n34330,n33479,n34333 );
   nand U35323 ( n34322,n34334,n34335 );
   nor U35324 ( n34335,n34336,n34337 );
   nor U35325 ( n34337,n33443,n34338 );
   nor U35326 ( n34336,n33433,n34339 );
   nor U35327 ( n34334,n34340,n34341 );
   nor U35328 ( n34341,n33465,n34342 );
   nor U35329 ( n34340,n33457,n34343 );
   nor U35330 ( n34296,n34344,n34345 );
   nor U35331 ( n34345,p3_ebx_reg_8_,n34346 );
   nand U35332 ( n34346,n34347,p3_ebx_reg_7_ );
   nor U35333 ( n34347,n28172,n34294 );
   nor U35334 ( n34344,n34348,n34349 );
   nor U35335 ( n34348,n34350,n34295 );
   nand U35336 ( n34295,n34236,n34351 );
   nand U35337 ( n34351,n34245,n34294 );
   nor U35338 ( n34350,p3_ebx_reg_7_,n28172 );
   nand U35339 ( n34353,n34233,n33903 );
   nand U35340 ( n33903,n34354,n34355 );
   nor U35341 ( n34355,n34356,n34357 );
   nand U35342 ( n34357,n34358,n34359 );
   nor U35343 ( n34359,n34360,n34361 );
   nor U35344 ( n34361,n33524,n34306 );
   nor U35345 ( n34360,n33521,n34307 );
   nor U35346 ( n34358,n34362,n34363 );
   nor U35347 ( n34363,n33534,n34310 );
   nor U35348 ( n34362,n33513,n34311 );
   nand U35349 ( n34356,n34364,n34365 );
   nor U35350 ( n34365,n34366,n34367 );
   nor U35351 ( n34367,n33512,n34316 );
   nor U35352 ( n34366,n33531,n34317 );
   nor U35353 ( n34364,n34368,n34369 );
   nor U35354 ( n34369,n33508,n34320 );
   nor U35355 ( n34368,n33503,n34321 );
   nor U35356 ( n34354,n34370,n34371 );
   nand U35357 ( n34371,n34372,n34373 );
   nor U35358 ( n34373,n34374,n34375 );
   nor U35359 ( n34375,n33530,n34328 );
   nor U35360 ( n34374,n33499,n34329 );
   nor U35361 ( n34372,n34376,n34377 );
   nor U35362 ( n34377,n33498,n34332 );
   nor U35363 ( n34376,n30716,n34333 );
   nand U35364 ( n34370,n34378,n34379 );
   nor U35365 ( n34379,n34380,n34381 );
   nor U35366 ( n34381,n33509,n34338 );
   nor U35367 ( n34380,n33502,n34339 );
   nor U35368 ( n34378,n34382,n34383 );
   nor U35369 ( n34383,n33525,n34342 );
   nor U35370 ( n34382,n33520,n34343 );
   nor U35371 ( n34352,n34384,n34385 );
   nor U35372 ( n34385,p3_ebx_reg_9_,n34386 );
   or U35373 ( n34386,n34387,n28173 );
   and U35374 ( n34384,n34388,p3_ebx_reg_9_ );
   nand U35375 ( n34390,n34233,n33917 );
   nand U35376 ( n33917,n34391,n34392 );
   nor U35377 ( n34392,n34393,n34394 );
   nand U35378 ( n34394,n34395,n34396 );
   nor U35379 ( n34396,n34397,n34398 );
   nor U35380 ( n34398,n33567,n34306 );
   nor U35381 ( n34397,n33564,n34307 );
   nor U35382 ( n34395,n34399,n34400 );
   nor U35383 ( n34400,n33558,n34310 );
   nor U35384 ( n34399,n33580,n34311 );
   nand U35385 ( n34393,n34401,n34402 );
   nor U35386 ( n34402,n34403,n34404 );
   nor U35387 ( n34404,n33579,n34316 );
   nor U35388 ( n34403,n33555,n34317 );
   nor U35389 ( n34401,n34405,n34406 );
   nor U35390 ( n34406,n33575,n34320 );
   nor U35391 ( n34405,n33590,n34321 );
   nor U35392 ( n34391,n34407,n34408 );
   nand U35393 ( n34408,n34409,n34410 );
   nor U35394 ( n34410,n34411,n34412 );
   nor U35395 ( n34412,n33554,n34328 );
   nor U35396 ( n34411,n33586,n34329 );
   nor U35397 ( n34409,n34413,n34414 );
   nor U35398 ( n34414,n33585,n34332 );
   nor U35399 ( n34413,n30705,n34333 );
   nand U35400 ( n34407,n34415,n34416 );
   nor U35401 ( n34416,n34417,n34418 );
   nor U35402 ( n34418,n33576,n34338 );
   nor U35403 ( n34417,n33589,n34339 );
   nor U35404 ( n34415,n34419,n34420 );
   nor U35405 ( n34420,n33568,n34342 );
   nor U35406 ( n34419,n33563,n34343 );
   nor U35407 ( n34389,n34421,n34422 );
   nor U35408 ( n34422,p3_ebx_reg_10_,n34423 );
   nand U35409 ( n34423,n34424,p3_ebx_reg_9_ );
   nor U35410 ( n34424,n28172,n34387 );
   nor U35411 ( n34421,n34425,n34426 );
   nor U35412 ( n34425,n34427,n34388 );
   nand U35413 ( n34388,n34236,n34428 );
   nand U35414 ( n34428,n34245,n34387 );
   nor U35415 ( n34427,p3_ebx_reg_9_,n28172 );
   nand U35416 ( n34430,n34233,n33928 );
   nand U35417 ( n33928,n34431,n34432 );
   nor U35418 ( n34432,n34433,n34434 );
   nand U35419 ( n34434,n34435,n34436 );
   nor U35420 ( n34436,n34437,n34438 );
   nor U35421 ( n34438,n33634,n34306 );
   nor U35422 ( n34437,n33631,n34307 );
   nor U35423 ( n34435,n34439,n34440 );
   nor U35424 ( n34440,n33644,n34310 );
   nor U35425 ( n34439,n33623,n34311 );
   nand U35426 ( n34433,n34441,n34442 );
   nor U35427 ( n34442,n34443,n34444 );
   nor U35428 ( n34444,n33622,n34316 );
   nor U35429 ( n34443,n33641,n34317 );
   nor U35430 ( n34441,n34445,n34446 );
   nor U35431 ( n34446,n33618,n34320 );
   nor U35432 ( n34445,n33613,n34321 );
   nor U35433 ( n34431,n34447,n34448 );
   nand U35434 ( n34448,n34449,n34450 );
   nor U35435 ( n34450,n34451,n34452 );
   nor U35436 ( n34452,n33640,n34328 );
   nor U35437 ( n34451,n33609,n34329 );
   nor U35438 ( n34449,n34453,n34454 );
   nor U35439 ( n34454,n33608,n34332 );
   nor U35440 ( n34453,n30694,n34333 );
   nand U35441 ( n34447,n34455,n34456 );
   nor U35442 ( n34456,n34457,n34458 );
   nor U35443 ( n34458,n33619,n34338 );
   nor U35444 ( n34457,n33612,n34339 );
   nor U35445 ( n34455,n34459,n34460 );
   nor U35446 ( n34460,n33635,n34342 );
   nor U35447 ( n34459,n33630,n34343 );
   nor U35448 ( n34429,n34461,n34462 );
   nor U35449 ( n34462,p3_ebx_reg_11_,n34463 );
   or U35450 ( n34463,n34464,n28173 );
   and U35451 ( n34461,n34465,p3_ebx_reg_11_ );
   nand U35452 ( n34467,n28283,n33942 );
   nand U35453 ( n33942,n34468,n34469 );
   nor U35454 ( n34469,n34470,n34471 );
   nand U35455 ( n34471,n34472,n34473 );
   nor U35456 ( n34473,n34474,n34475 );
   nor U35457 ( n34475,n33678,n34306 );
   nor U35458 ( n34474,n33675,n34307 );
   nor U35459 ( n34472,n34476,n34477 );
   nor U35460 ( n34477,n33669,n34310 );
   nor U35461 ( n34476,n33691,n34311 );
   nand U35462 ( n34470,n34478,n34479 );
   nor U35463 ( n34479,n34480,n34481 );
   nor U35464 ( n34481,n33690,n34316 );
   nor U35465 ( n34480,n33666,n34317 );
   nor U35466 ( n34478,n34482,n34483 );
   nor U35467 ( n34483,n33686,n34320 );
   nor U35468 ( n34482,n33701,n34321 );
   nor U35469 ( n34468,n34484,n34485 );
   nand U35470 ( n34485,n34486,n34487 );
   nor U35471 ( n34487,n34488,n34489 );
   nor U35472 ( n34489,n33665,n34328 );
   nor U35473 ( n34488,n33697,n34329 );
   nor U35474 ( n34486,n34490,n34491 );
   nor U35475 ( n34491,n33696,n34332 );
   nor U35476 ( n34490,n30683,n34333 );
   nand U35477 ( n34484,n34492,n34493 );
   nor U35478 ( n34493,n34494,n34495 );
   nor U35479 ( n34495,n33687,n34338 );
   nor U35480 ( n34494,n33700,n34339 );
   nor U35481 ( n34492,n34496,n34497 );
   nor U35482 ( n34497,n33679,n34342 );
   nor U35483 ( n34496,n33674,n34343 );
   nor U35484 ( n34466,n34498,n34499 );
   nor U35485 ( n34499,p3_ebx_reg_12_,n34500 );
   nand U35486 ( n34500,n34501,p3_ebx_reg_11_ );
   nor U35487 ( n34501,n28172,n34464 );
   nor U35488 ( n34498,n34502,n34503 );
   nor U35489 ( n34502,n34504,n34465 );
   nand U35490 ( n34465,n34236,n34505 );
   nand U35491 ( n34505,n34245,n34464 );
   nor U35492 ( n34504,p3_ebx_reg_11_,n28171 );
   nand U35493 ( n34507,n28283,n33953 );
   nand U35494 ( n33953,n34508,n34509 );
   nor U35495 ( n34509,n34510,n34511 );
   nand U35496 ( n34511,n34512,n34513 );
   nor U35497 ( n34513,n34514,n34515 );
   nor U35498 ( n34515,n33732,n34306 );
   nor U35499 ( n34514,n33729,n34307 );
   nor U35500 ( n34512,n34516,n34517 );
   nor U35501 ( n34517,n33723,n34310 );
   nor U35502 ( n34516,n33745,n34311 );
   nand U35503 ( n34510,n34518,n34519 );
   nor U35504 ( n34519,n34520,n34521 );
   nor U35505 ( n34521,n33744,n34316 );
   nor U35506 ( n34520,n33720,n34317 );
   nor U35507 ( n34518,n34522,n34523 );
   nor U35508 ( n34523,n33740,n34320 );
   nor U35509 ( n34522,n33755,n34321 );
   nor U35510 ( n34508,n34524,n34525 );
   nand U35511 ( n34525,n34526,n34527 );
   nor U35512 ( n34527,n34528,n34529 );
   nor U35513 ( n34529,n33719,n34328 );
   nor U35514 ( n34528,n33751,n34329 );
   nor U35515 ( n34526,n34530,n34531 );
   nor U35516 ( n34531,n33750,n34332 );
   nor U35517 ( n34530,n30673,n34333 );
   nand U35518 ( n34524,n34532,n34533 );
   nor U35519 ( n34533,n34534,n34535 );
   nor U35520 ( n34535,n33741,n34338 );
   nor U35521 ( n34534,n33754,n34339 );
   nor U35522 ( n34532,n34536,n34537 );
   nor U35523 ( n34537,n33733,n34342 );
   nor U35524 ( n34536,n33728,n34343 );
   nor U35525 ( n34506,n34538,n34539 );
   nor U35526 ( n34539,p3_ebx_reg_13_,n34540 );
   or U35527 ( n34540,n34541,n28173 );
   and U35528 ( n34538,n34542,p3_ebx_reg_13_ );
   nand U35529 ( n34544,n34233,n33967 );
   nand U35530 ( n33967,n34545,n34546 );
   nor U35531 ( n34546,n34547,n34548 );
   nand U35532 ( n34548,n34549,n34550 );
   nor U35533 ( n34550,n34551,n34552 );
   nor U35534 ( n34552,n33802,n34306 );
   nor U35535 ( n34551,n33799,n34307 );
   nor U35536 ( n34549,n34553,n34554 );
   nor U35537 ( n34554,n33812,n34310 );
   nor U35538 ( n34553,n33791,n34311 );
   nand U35539 ( n34547,n34555,n34556 );
   nor U35540 ( n34556,n34557,n34558 );
   nor U35541 ( n34558,n33790,n34316 );
   nor U35542 ( n34557,n33809,n34317 );
   nor U35543 ( n34555,n34559,n34560 );
   nor U35544 ( n34560,n33786,n34320 );
   nor U35545 ( n34559,n33781,n34321 );
   nor U35546 ( n34545,n34561,n34562 );
   nand U35547 ( n34562,n34563,n34564 );
   nor U35548 ( n34564,n34565,n34566 );
   nor U35549 ( n34566,n33808,n34328 );
   nor U35550 ( n34565,n33777,n34329 );
   nor U35551 ( n34563,n34567,n34568 );
   nor U35552 ( n34568,n33776,n34332 );
   nor U35553 ( n34567,n30662,n34333 );
   nand U35554 ( n34561,n34569,n34570 );
   nor U35555 ( n34570,n34571,n34572 );
   nor U35556 ( n34572,n33787,n34338 );
   nor U35557 ( n34571,n33780,n34339 );
   nor U35558 ( n34569,n34573,n34574 );
   nor U35559 ( n34574,n33803,n34342 );
   nor U35560 ( n34573,n33798,n34343 );
   nor U35561 ( n34543,n34575,n34576 );
   nor U35562 ( n34576,p3_ebx_reg_14_,n34577 );
   nand U35563 ( n34577,n34578,p3_ebx_reg_13_ );
   nor U35564 ( n34578,n28173,n34541 );
   nor U35565 ( n34575,n34579,n34580 );
   nor U35566 ( n34579,n34581,n34542 );
   nand U35567 ( n34542,n34236,n34582 );
   nand U35568 ( n34582,n34245,n34541 );
   nor U35569 ( n34581,p3_ebx_reg_13_,n28173 );
   nand U35570 ( n34584,n34233,n33978 );
   nand U35571 ( n33978,n34585,n34586 );
   nor U35572 ( n34586,n34587,n34588 );
   nand U35573 ( n34588,n34589,n34590 );
   nor U35574 ( n34590,n34591,n34592 );
   nor U35575 ( n34592,n33863,n34306 );
   nand U35576 ( n34306,n34593,n34594 );
   nor U35577 ( n34591,n33859,n34307 );
   nand U35578 ( n34307,n34593,n29294 );
   nor U35579 ( n34589,n34595,n34596 );
   nor U35580 ( n34596,n33876,n34310 );
   nand U35581 ( n34310,n34593,n34597 );
   nor U35582 ( n34595,n33851,n34311 );
   nand U35583 ( n34311,n34598,n34594 );
   nand U35584 ( n34587,n34599,n34600 );
   nor U35585 ( n34600,n34601,n34602 );
   nor U35586 ( n34602,n33849,n34316 );
   nand U35587 ( n34316,n34598,n29294 );
   nor U35588 ( n34601,n33872,n34317 );
   nand U35589 ( n34317,n34598,n34597 );
   nor U35590 ( n34599,n34603,n34604 );
   nor U35591 ( n34604,n33845,n34320 );
   nand U35592 ( n34320,n34605,n34594 );
   nor U35593 ( n34603,n33839,n34321 );
   nand U35594 ( n34321,n34605,n29294 );
   nor U35595 ( n34585,n34606,n34607 );
   nand U35596 ( n34607,n34608,n34609 );
   nor U35597 ( n34609,n34610,n34611 );
   nor U35598 ( n34611,n33869,n34328 );
   nand U35599 ( n34328,n34605,n34597 );
   nor U35600 ( n34610,n33833,n34329 );
   nand U35601 ( n34329,n34612,n34594 );
   nor U35602 ( n34608,n34613,n34614 );
   nor U35603 ( n34614,n33830,n34332 );
   nand U35604 ( n34332,n34612,n29294 );
   nor U35605 ( n34613,n30650,n34333 );
   nand U35606 ( n34333,n34612,n34597 );
   nand U35607 ( n34606,n34615,n34616 );
   nor U35608 ( n34616,n34617,n34618 );
   nor U35609 ( n34618,n33846,n34338 );
   nand U35610 ( n34338,n34605,n34619 );
   and U35611 ( n34605,n34620,n29261 );
   nor U35612 ( n34617,n33837,n34339 );
   nand U35613 ( n34339,n34612,n34619 );
   and U35614 ( n34612,n29261,n29312 );
   nor U35615 ( n34615,n34621,n34622 );
   nor U35616 ( n34622,n33864,n34342 );
   nand U35617 ( n34342,n34593,n34619 );
   nor U35618 ( n34593,n29261,n29312 );
   nor U35619 ( n34621,n33858,n34343 );
   nand U35620 ( n34343,n34598,n34619 );
   nor U35621 ( n34598,n29261,n34620 );
   not U35622 ( n34620,n29312 );
   nand U35623 ( n29312,n29267,n34623 );
   nand U35624 ( n34623,n29341,n29257 );
   nand U35625 ( n29261,n34624,n34625 );
   nand U35626 ( n34625,n34626,n29254 );
   nand U35627 ( n34626,n34627,p3_instqueuerd_addr_reg_1_ );
   or U35628 ( n34624,n29267,n34627 );
   nand U35629 ( n29267,p3_instqueuerd_addr_reg_2_,p3_instqueuerd_addr_reg_1_ );
   nor U35630 ( n34583,n34628,n34629 );
   nor U35631 ( n34629,p3_ebx_reg_15_,n34630 );
   or U35632 ( n34630,n34631,n28173 );
   and U35633 ( n34628,n34632,p3_ebx_reg_15_ );
   nand U35634 ( n34634,n34233,n33985 );
   nand U35635 ( n33985,n34635,n34636 );
   nor U35636 ( n34636,n34637,n34638 );
   nand U35637 ( n34638,n34639,n34640 );
   nor U35638 ( n34640,n34641,n34642 );
   nor U35639 ( n34642,n33441,n34643 );
   nor U35640 ( n34641,n33435,n34644 );
   nor U35641 ( n34639,n34645,n34646 );
   nor U35642 ( n34646,n33471,n34647 );
   nor U35643 ( n34645,n33429,n34648 );
   nand U35644 ( n34637,n34649,n34650 );
   nor U35645 ( n34650,n34651,n34652 );
   nor U35646 ( n34652,n33427,n34653 );
   nor U35647 ( n34651,n33479,n34654 );
   nor U35648 ( n34649,n34655,n34656 );
   nor U35649 ( n34656,n33463,n34657 );
   nor U35650 ( n34655,n33459,n34658 );
   nor U35651 ( n34635,n34659,n34660 );
   nand U35652 ( n34660,n34661,n34662 );
   nor U35653 ( n34662,n34663,n34664 );
   nor U35654 ( n34664,n33477,n34665 );
   nor U35655 ( n34663,n33449,n34666 );
   nor U35656 ( n34661,n34667,n34668 );
   nor U35657 ( n34668,n33447,n34669 );
   nor U35658 ( n34667,n33473,n34670 );
   nand U35659 ( n34659,n34671,n34672 );
   nor U35660 ( n34672,n34673,n34674 );
   nor U35661 ( n34674,n33443,n34675 );
   nor U35662 ( n34673,n33433,n34676 );
   nor U35663 ( n34671,n34677,n34678 );
   nor U35664 ( n34678,n33465,n34679 );
   nor U35665 ( n34677,n33457,n34680 );
   nor U35666 ( n34633,n34681,n34682 );
   nor U35667 ( n34682,p3_ebx_reg_16_,n34683 );
   nand U35668 ( n34683,n34684,p3_ebx_reg_15_ );
   nor U35669 ( n34684,n28171,n34631 );
   nor U35670 ( n34681,n34685,n34686 );
   nor U35671 ( n34685,n34687,n34632 );
   nand U35672 ( n34632,n34236,n34688 );
   nand U35673 ( n34688,n34245,n34631 );
   nor U35674 ( n34687,p3_ebx_reg_15_,n28172 );
   nand U35675 ( n34690,n28283,n34002 );
   nand U35676 ( n34002,n34691,n34692 );
   nor U35677 ( n34692,n34693,n34694 );
   nand U35678 ( n34694,n34695,n34696 );
   nor U35679 ( n34696,n34697,n34698 );
   nor U35680 ( n34698,n33508,n34643 );
   nor U35681 ( n34697,n33503,n34644 );
   nor U35682 ( n34695,n34699,n34700 );
   nor U35683 ( n34700,n33530,n34647 );
   nor U35684 ( n34699,n33499,n34648 );
   nand U35685 ( n34693,n34701,n34702 );
   nor U35686 ( n34702,n34703,n34704 );
   nor U35687 ( n34704,n33498,n34653 );
   nor U35688 ( n34703,n30716,n34654 );
   nor U35689 ( n34701,n34705,n34706 );
   nor U35690 ( n34706,n33524,n34657 );
   nor U35691 ( n34705,n33521,n34658 );
   nor U35692 ( n34691,n34707,n34708 );
   nand U35693 ( n34708,n34709,n34710 );
   nor U35694 ( n34710,n34711,n34712 );
   nor U35695 ( n34712,n33534,n34665 );
   nor U35696 ( n34711,n33513,n34666 );
   nor U35697 ( n34709,n34713,n34714 );
   nor U35698 ( n34714,n33512,n34669 );
   nor U35699 ( n34713,n33531,n34670 );
   nand U35700 ( n34707,n34715,n34716 );
   nor U35701 ( n34716,n34717,n34718 );
   nor U35702 ( n34718,n33509,n34675 );
   nor U35703 ( n34717,n33502,n34676 );
   nor U35704 ( n34715,n34719,n34720 );
   nor U35705 ( n34720,n33525,n34679 );
   nor U35706 ( n34719,n33520,n34680 );
   nor U35707 ( n34689,n34721,n34722 );
   nor U35708 ( n34722,p3_ebx_reg_17_,n34723 );
   or U35709 ( n34723,n34724,n28172 );
   and U35710 ( n34721,n34725,p3_ebx_reg_17_ );
   nand U35711 ( n34727,n28283,n34015 );
   nand U35712 ( n34015,n34728,n34729 );
   nor U35713 ( n34729,n34730,n34731 );
   nand U35714 ( n34731,n34732,n34733 );
   nor U35715 ( n34733,n34734,n34735 );
   nor U35716 ( n34735,n33575,n34643 );
   nor U35717 ( n34734,n33590,n34644 );
   nor U35718 ( n34732,n34736,n34737 );
   nor U35719 ( n34737,n33554,n34647 );
   nor U35720 ( n34736,n33586,n34648 );
   nand U35721 ( n34730,n34738,n34739 );
   nor U35722 ( n34739,n34740,n34741 );
   nor U35723 ( n34741,n33585,n34653 );
   nor U35724 ( n34740,n30705,n34654 );
   nor U35725 ( n34738,n34742,n34743 );
   nor U35726 ( n34743,n33567,n34657 );
   nor U35727 ( n34742,n33564,n34658 );
   nor U35728 ( n34728,n34744,n34745 );
   nand U35729 ( n34745,n34746,n34747 );
   nor U35730 ( n34747,n34748,n34749 );
   nor U35731 ( n34749,n33558,n34665 );
   nor U35732 ( n34748,n33580,n34666 );
   nor U35733 ( n34746,n34750,n34751 );
   nor U35734 ( n34751,n33579,n34669 );
   nor U35735 ( n34750,n33555,n34670 );
   nand U35736 ( n34744,n34752,n34753 );
   nor U35737 ( n34753,n34754,n34755 );
   nor U35738 ( n34755,n33576,n34675 );
   nor U35739 ( n34754,n33589,n34676 );
   nor U35740 ( n34752,n34756,n34757 );
   nor U35741 ( n34757,n33568,n34679 );
   nor U35742 ( n34756,n33563,n34680 );
   nor U35743 ( n34726,n34758,n34759 );
   nor U35744 ( n34759,p3_ebx_reg_18_,n34760 );
   nand U35745 ( n34760,n34761,p3_ebx_reg_17_ );
   nor U35746 ( n34761,n28171,n34724 );
   nor U35747 ( n34758,n34762,n34763 );
   nor U35748 ( n34762,n34764,n34725 );
   nand U35749 ( n34725,n34236,n34765 );
   nand U35750 ( n34765,n34245,n34724 );
   nor U35751 ( n34764,p3_ebx_reg_17_,n28173 );
   nand U35752 ( n34767,n28283,n34031 );
   nand U35753 ( n34031,n34768,n34769 );
   nor U35754 ( n34769,n34770,n34771 );
   nand U35755 ( n34771,n34772,n34773 );
   nor U35756 ( n34773,n34774,n34775 );
   nor U35757 ( n34775,n33618,n34643 );
   nor U35758 ( n34774,n33613,n34644 );
   nor U35759 ( n34772,n34776,n34777 );
   nor U35760 ( n34777,n33640,n34647 );
   nor U35761 ( n34776,n33609,n34648 );
   nand U35762 ( n34770,n34778,n34779 );
   nor U35763 ( n34779,n34780,n34781 );
   nor U35764 ( n34781,n33608,n34653 );
   nor U35765 ( n34780,n30694,n34654 );
   nor U35766 ( n34778,n34782,n34783 );
   nor U35767 ( n34783,n33634,n34657 );
   nor U35768 ( n34782,n33631,n34658 );
   nor U35769 ( n34768,n34784,n34785 );
   nand U35770 ( n34785,n34786,n34787 );
   nor U35771 ( n34787,n34788,n34789 );
   nor U35772 ( n34789,n33644,n34665 );
   nor U35773 ( n34788,n33623,n34666 );
   nor U35774 ( n34786,n34790,n34791 );
   nor U35775 ( n34791,n33622,n34669 );
   nor U35776 ( n34790,n33641,n34670 );
   nand U35777 ( n34784,n34792,n34793 );
   nor U35778 ( n34793,n34794,n34795 );
   nor U35779 ( n34795,n33619,n34675 );
   nor U35780 ( n34794,n33612,n34676 );
   nor U35781 ( n34792,n34796,n34797 );
   nor U35782 ( n34797,n33635,n34679 );
   nor U35783 ( n34796,n33630,n34680 );
   nor U35784 ( n34766,n34798,n34799 );
   nor U35785 ( n34799,p3_ebx_reg_19_,n34800 );
   or U35786 ( n34800,n34801,n28171 );
   and U35787 ( n34798,n34802,p3_ebx_reg_19_ );
   nand U35788 ( n34804,n28283,n34044 );
   nand U35789 ( n34044,n34805,n34806 );
   nor U35790 ( n34806,n34807,n34808 );
   nand U35791 ( n34808,n34809,n34810 );
   nor U35792 ( n34810,n34811,n34812 );
   nor U35793 ( n34812,n33686,n34643 );
   nor U35794 ( n34811,n33701,n34644 );
   nor U35795 ( n34809,n34813,n34814 );
   nor U35796 ( n34814,n33665,n34647 );
   nor U35797 ( n34813,n33697,n34648 );
   nand U35798 ( n34807,n34815,n34816 );
   nor U35799 ( n34816,n34817,n34818 );
   nor U35800 ( n34818,n33696,n34653 );
   nor U35801 ( n34817,n30683,n34654 );
   nor U35802 ( n34815,n34819,n34820 );
   nor U35803 ( n34820,n33678,n34657 );
   nor U35804 ( n34819,n33675,n34658 );
   nor U35805 ( n34805,n34821,n34822 );
   nand U35806 ( n34822,n34823,n34824 );
   nor U35807 ( n34824,n34825,n34826 );
   nor U35808 ( n34826,n33669,n34665 );
   nor U35809 ( n34825,n33691,n34666 );
   nor U35810 ( n34823,n34827,n34828 );
   nor U35811 ( n34828,n33690,n34669 );
   nor U35812 ( n34827,n33666,n34670 );
   nand U35813 ( n34821,n34829,n34830 );
   nor U35814 ( n34830,n34831,n34832 );
   nor U35815 ( n34832,n33687,n34675 );
   nor U35816 ( n34831,n33700,n34676 );
   nor U35817 ( n34829,n34833,n34834 );
   nor U35818 ( n34834,n33679,n34679 );
   nor U35819 ( n34833,n33674,n34680 );
   nor U35820 ( n34803,n34835,n34836 );
   nor U35821 ( n34836,p3_ebx_reg_20_,n34837 );
   nand U35822 ( n34837,n34838,p3_ebx_reg_19_ );
   nor U35823 ( n34838,n28172,n34801 );
   nor U35824 ( n34835,n34839,n34840 );
   nor U35825 ( n34839,n34841,n34802 );
   nand U35826 ( n34802,n34236,n34842 );
   nand U35827 ( n34842,n34245,n34801 );
   nor U35828 ( n34841,p3_ebx_reg_19_,n28171 );
   nand U35829 ( n34844,n28283,n34061 );
   nand U35830 ( n34061,n34845,n34846 );
   nor U35831 ( n34846,n34847,n34848 );
   nand U35832 ( n34848,n34849,n34850 );
   nor U35833 ( n34850,n34851,n34852 );
   nor U35834 ( n34852,n33740,n34643 );
   nor U35835 ( n34851,n33755,n34644 );
   nor U35836 ( n34849,n34853,n34854 );
   nor U35837 ( n34854,n33719,n34647 );
   nor U35838 ( n34853,n33751,n34648 );
   nand U35839 ( n34847,n34855,n34856 );
   nor U35840 ( n34856,n34857,n34858 );
   nor U35841 ( n34858,n33750,n34653 );
   nor U35842 ( n34857,n30673,n34654 );
   nor U35843 ( n34855,n34859,n34860 );
   nor U35844 ( n34860,n33732,n34657 );
   nor U35845 ( n34859,n33729,n34658 );
   nor U35846 ( n34845,n34861,n34862 );
   nand U35847 ( n34862,n34863,n34864 );
   nor U35848 ( n34864,n34865,n34866 );
   nor U35849 ( n34866,n33723,n34665 );
   nor U35850 ( n34865,n33745,n34666 );
   nor U35851 ( n34863,n34867,n34868 );
   nor U35852 ( n34868,n33744,n34669 );
   nor U35853 ( n34867,n33720,n34670 );
   nand U35854 ( n34861,n34869,n34870 );
   nor U35855 ( n34870,n34871,n34872 );
   nor U35856 ( n34872,n33741,n34675 );
   nor U35857 ( n34871,n33754,n34676 );
   nor U35858 ( n34869,n34873,n34874 );
   nor U35859 ( n34874,n33733,n34679 );
   nor U35860 ( n34873,n33728,n34680 );
   nor U35861 ( n34843,n34875,n34876 );
   nor U35862 ( n34876,p3_ebx_reg_21_,n34877 );
   or U35863 ( n34877,n34878,n28173 );
   and U35864 ( n34875,n34879,p3_ebx_reg_21_ );
   nand U35865 ( n34881,n28283,n34074 );
   nand U35866 ( n34074,n34882,n34883 );
   nor U35867 ( n34883,n34884,n34885 );
   nand U35868 ( n34885,n34886,n34887 );
   nor U35869 ( n34887,n34888,n34889 );
   nor U35870 ( n34889,n33786,n34643 );
   nor U35871 ( n34888,n33781,n34644 );
   nor U35872 ( n34886,n34890,n34891 );
   nor U35873 ( n34891,n33808,n34647 );
   nor U35874 ( n34890,n33777,n34648 );
   nand U35875 ( n34884,n34892,n34893 );
   nor U35876 ( n34893,n34894,n34895 );
   nor U35877 ( n34895,n33776,n34653 );
   nor U35878 ( n34894,n30662,n34654 );
   nor U35879 ( n34892,n34896,n34897 );
   nor U35880 ( n34897,n33802,n34657 );
   nor U35881 ( n34896,n33799,n34658 );
   nor U35882 ( n34882,n34898,n34899 );
   nand U35883 ( n34899,n34900,n34901 );
   nor U35884 ( n34901,n34902,n34903 );
   nor U35885 ( n34903,n33812,n34665 );
   nor U35886 ( n34902,n33791,n34666 );
   nor U35887 ( n34900,n34904,n34905 );
   nor U35888 ( n34905,n33790,n34669 );
   nor U35889 ( n34904,n33809,n34670 );
   nand U35890 ( n34898,n34906,n34907 );
   nor U35891 ( n34907,n34908,n34909 );
   nor U35892 ( n34909,n33787,n34675 );
   nor U35893 ( n34908,n33780,n34676 );
   nor U35894 ( n34906,n34910,n34911 );
   nor U35895 ( n34911,n33803,n34679 );
   nor U35896 ( n34910,n33798,n34680 );
   nor U35897 ( n34880,n34912,n34913 );
   nor U35898 ( n34913,p3_ebx_reg_22_,n34914 );
   nand U35899 ( n34914,n34915,p3_ebx_reg_21_ );
   nor U35900 ( n34915,n28171,n34878 );
   nor U35901 ( n34912,n34916,n34917 );
   nor U35902 ( n34916,n34918,n34879 );
   nand U35903 ( n34879,n34236,n34919 );
   nand U35904 ( n34919,n34245,n34878 );
   nor U35905 ( n34918,p3_ebx_reg_21_,n28171 );
   nand U35906 ( n34921,n28283,n34090 );
   xor U35907 ( n34090,n34922,n34923 );
   nor U35908 ( n34920,n34924,n34925 );
   nor U35909 ( n34925,p3_ebx_reg_23_,n34926 );
   or U35910 ( n34926,n34927,n28171 );
   and U35911 ( n34924,n34928,p3_ebx_reg_23_ );
   nand U35912 ( n34930,n28283,n34931 );
   not U35913 ( n34931,n34102 );
   nand U35914 ( n34102,n34932,n34933 );
   nand U35915 ( n34933,n34934,n34935 );
   nand U35916 ( n34935,n34923,n34922 );
   not U35917 ( n34934,n34936 );
   nor U35918 ( n34929,n34937,n34938 );
   nor U35919 ( n34938,p3_ebx_reg_24_,n34939 );
   nand U35920 ( n34939,n34940,p3_ebx_reg_23_ );
   nor U35921 ( n34940,n28173,n34927 );
   nor U35922 ( n34937,n34941,n34942 );
   nor U35923 ( n34941,n34943,n34928 );
   nand U35924 ( n34928,n34236,n34944 );
   nand U35925 ( n34944,n34245,n34927 );
   nor U35926 ( n34943,p3_ebx_reg_23_,n28171 );
   nand U35927 ( n34946,n34947,n28283 );
   nor U35928 ( n34947,n34120,n34119 );
   nor U35929 ( n34119,n34948,n34949 );
   nor U35930 ( n34945,n34950,n34951 );
   nor U35931 ( n34951,p3_ebx_reg_25_,n34952 );
   or U35932 ( n34952,n34953,n28172 );
   and U35933 ( n34950,n34954,p3_ebx_reg_25_ );
   nand U35934 ( n34956,n28283,n34957 );
   not U35935 ( n34957,n34132 );
   xor U35936 ( n34132,n34958,n34120 );
   nor U35937 ( n34955,n34959,n34960 );
   nor U35938 ( n34960,p3_ebx_reg_26_,n34961 );
   nand U35939 ( n34961,n34962,p3_ebx_reg_25_ );
   nor U35940 ( n34962,n28172,n34953 );
   nor U35941 ( n34959,n34963,n34964 );
   nor U35942 ( n34963,n34965,n34954 );
   nand U35943 ( n34954,n34236,n34966 );
   nand U35944 ( n34966,n34245,n34953 );
   nor U35945 ( n34965,p3_ebx_reg_25_,n28173 );
   nand U35946 ( n34968,n34969,n28283 );
   and U35947 ( n34969,n34149,n34148 );
   nand U35948 ( n34148,n34970,n34971 );
   nand U35949 ( n34971,n34120,n34972 );
   nor U35950 ( n34967,n34973,n34974 );
   nor U35951 ( n34974,p3_ebx_reg_27_,n34975 );
   or U35952 ( n34975,n34976,n28171 );
   and U35953 ( n34973,n34977,p3_ebx_reg_27_ );
   nand U35954 ( n34979,n28283,n34980 );
   not U35955 ( n34980,n34161 );
   xor U35956 ( n34161,n34981,n34149 );
   nor U35957 ( n34978,n34982,n34983 );
   nor U35958 ( n34983,p3_ebx_reg_28_,n34984 );
   nand U35959 ( n34984,n34985,p3_ebx_reg_27_ );
   nor U35960 ( n34985,n28173,n34976 );
   nor U35961 ( n34982,n34986,n34987 );
   nor U35962 ( n34986,n34988,n34977 );
   nand U35963 ( n34977,n34236,n34989 );
   nand U35964 ( n34989,n34245,n34976 );
   nor U35965 ( n34988,p3_ebx_reg_27_,n28171 );
   nand U35966 ( n34991,n34233,n34183 );
   xor U35967 ( n34183,n34992,n34993 );
   nor U35968 ( n34990,n34994,n34995 );
   and U35969 ( n34995,n34996,n34997 );
   nor U35970 ( n34994,n34998,n34996 );
   nand U35971 ( n35000,n34233,n34192 );
   xor U35972 ( n34192,n35001,n35002 );
   nand U35973 ( n35002,n35003,n35004 );
   nor U35974 ( n35004,n35005,n35006 );
   nand U35975 ( n35006,n35007,n35008 );
   nor U35976 ( n35008,n35009,n35010 );
   nor U35977 ( n35010,n33839,n35011 );
   nor U35978 ( n35009,n33845,n35012 );
   nor U35979 ( n35007,n35013,n35014 );
   nor U35980 ( n35014,n33833,n35015 );
   nor U35981 ( n35013,n33869,n35016 );
   nand U35982 ( n35005,n35017,n35018 );
   nor U35983 ( n35018,n35019,n35020 );
   nor U35984 ( n35020,n30650,n35021 );
   nor U35985 ( n35019,n33830,n35022 );
   nor U35986 ( n35017,n35023,n35024 );
   nor U35987 ( n35024,n33859,n35025 );
   nor U35988 ( n35023,n33863,n35026 );
   nor U35989 ( n35003,n35027,n35028 );
   nand U35990 ( n35028,n35029,n35030 );
   nor U35991 ( n35030,n35031,n35032 );
   nor U35992 ( n35032,n33851,n35033 );
   nor U35993 ( n35031,n33876,n35034 );
   nor U35994 ( n35029,n35035,n35036 );
   nor U35995 ( n35036,n33872,n35037 );
   nor U35996 ( n35035,n33849,n35038 );
   nand U35997 ( n35027,n35039,n35040 );
   nor U35998 ( n35040,n35041,n35042 );
   nor U35999 ( n35042,n33837,n35043 );
   nor U36000 ( n35041,n33846,n35044 );
   nor U36001 ( n35039,n35045,n35046 );
   nor U36002 ( n35046,n33858,n35047 );
   nor U36003 ( n35045,n33864,n35048 );
   nor U36004 ( n35001,n34992,n34993 );
   nand U36005 ( n34993,n35049,n34981 );
   nand U36006 ( n34981,n35050,n35051 );
   nor U36007 ( n35051,n35052,n35053 );
   nand U36008 ( n35053,n35054,n35055 );
   nor U36009 ( n35055,n35056,n35057 );
   nor U36010 ( n35057,n33728,n35047 );
   nor U36011 ( n35056,n33733,n35048 );
   nor U36012 ( n35054,n35058,n35059 );
   nor U36013 ( n35059,n33754,n35043 );
   nor U36014 ( n35058,n33741,n35044 );
   nand U36015 ( n35052,n35060,n35061 );
   nor U36016 ( n35061,n35062,n35063 );
   nor U36017 ( n35063,n33720,n35037 );
   nor U36018 ( n35062,n33744,n35038 );
   nor U36019 ( n35060,n35064,n35065 );
   nor U36020 ( n35065,n33745,n35033 );
   nor U36021 ( n35064,n33723,n35034 );
   nor U36022 ( n35050,n35066,n35067 );
   nand U36023 ( n35067,n35068,n35069 );
   nor U36024 ( n35069,n35070,n35071 );
   nor U36025 ( n35071,n33729,n35025 );
   nor U36026 ( n35070,n33732,n35026 );
   nor U36027 ( n35068,n35072,n35073 );
   nor U36028 ( n35073,n30673,n35021 );
   nor U36029 ( n35072,n33750,n35022 );
   nand U36030 ( n35066,n35074,n35075 );
   nor U36031 ( n35075,n35076,n35077 );
   nor U36032 ( n35077,n33751,n35015 );
   nor U36033 ( n35076,n33719,n35016 );
   nor U36034 ( n35074,n35078,n35079 );
   nor U36035 ( n35079,n33755,n35011 );
   nor U36036 ( n35078,n33740,n35012 );
   not U36037 ( n35049,n34149 );
   nand U36038 ( n34149,n35080,n34120 );
   and U36039 ( n34120,n34949,n34948 );
   nand U36040 ( n34948,n35081,n35082 );
   nor U36041 ( n35082,n35083,n35084 );
   nand U36042 ( n35084,n35085,n35086 );
   nor U36043 ( n35086,n35087,n35088 );
   nor U36044 ( n35088,n33563,n35047 );
   nor U36045 ( n35087,n33568,n35048 );
   nor U36046 ( n35085,n35089,n35090 );
   nor U36047 ( n35090,n33589,n35043 );
   nor U36048 ( n35089,n33576,n35044 );
   nand U36049 ( n35083,n35091,n35092 );
   nor U36050 ( n35092,n35093,n35094 );
   nor U36051 ( n35094,n33555,n35037 );
   nor U36052 ( n35093,n33579,n35038 );
   nor U36053 ( n35091,n35095,n35096 );
   nor U36054 ( n35096,n33580,n35033 );
   nor U36055 ( n35095,n33558,n35034 );
   nor U36056 ( n35081,n35097,n35098 );
   nand U36057 ( n35098,n35099,n35100 );
   nor U36058 ( n35100,n35101,n35102 );
   nor U36059 ( n35102,n33564,n35025 );
   nor U36060 ( n35101,n33567,n35026 );
   nor U36061 ( n35099,n35103,n35104 );
   nor U36062 ( n35104,n30705,n35021 );
   nor U36063 ( n35103,n33585,n35022 );
   nand U36064 ( n35097,n35105,n35106 );
   nor U36065 ( n35106,n35107,n35108 );
   nor U36066 ( n35108,n33586,n35015 );
   nor U36067 ( n35107,n33554,n35016 );
   nor U36068 ( n35105,n35109,n35110 );
   nor U36069 ( n35110,n33590,n35011 );
   nor U36070 ( n35109,n33575,n35012 );
   not U36071 ( n34949,n34932 );
   nand U36072 ( n34932,n35111,n34936 );
   nand U36073 ( n34936,n35112,n35113 );
   nor U36074 ( n35113,n35114,n35115 );
   nand U36075 ( n35115,n35116,n35117 );
   nor U36076 ( n35117,n35118,n35119 );
   nor U36077 ( n35119,n33520,n35047 );
   nor U36078 ( n35118,n33525,n35048 );
   nor U36079 ( n35116,n35120,n35121 );
   nor U36080 ( n35121,n33502,n35043 );
   nor U36081 ( n35120,n33509,n35044 );
   nand U36082 ( n35114,n35122,n35123 );
   nor U36083 ( n35123,n35124,n35125 );
   nor U36084 ( n35125,n33531,n35037 );
   nor U36085 ( n35124,n33512,n35038 );
   nor U36086 ( n35122,n35126,n35127 );
   nor U36087 ( n35127,n33513,n35033 );
   nor U36088 ( n35126,n33534,n35034 );
   nor U36089 ( n35112,n35128,n35129 );
   nand U36090 ( n35129,n35130,n35131 );
   nor U36091 ( n35131,n35132,n35133 );
   nor U36092 ( n35133,n33521,n35025 );
   nor U36093 ( n35132,n33524,n35026 );
   nor U36094 ( n35130,n35134,n35135 );
   nor U36095 ( n35135,n30716,n35021 );
   nor U36096 ( n35134,n33498,n35022 );
   nand U36097 ( n35128,n35136,n35137 );
   nor U36098 ( n35137,n35138,n35139 );
   nor U36099 ( n35139,n33499,n35015 );
   nor U36100 ( n35138,n33530,n35016 );
   nor U36101 ( n35136,n35140,n35141 );
   nor U36102 ( n35141,n33503,n35011 );
   nor U36103 ( n35140,n33508,n35012 );
   and U36104 ( n35111,n34923,n34922 );
   nand U36105 ( n34922,n35142,n35143 );
   nor U36106 ( n35143,n35144,n35145 );
   nand U36107 ( n35145,n35146,n35147 );
   nor U36108 ( n35147,n35148,n35149 );
   nor U36109 ( n35149,n33846,n34675 );
   nand U36110 ( n34675,n35150,n33832 );
   nor U36111 ( n35148,n33837,n34676 );
   nand U36112 ( n34676,n35151,n33832 );
   nor U36113 ( n35146,n35152,n35153 );
   nor U36114 ( n35153,n33864,n34679 );
   nand U36115 ( n34679,n35154,n33832 );
   nor U36116 ( n35152,n33858,n34680 );
   nand U36117 ( n34680,n35155,n33832 );
   nor U36118 ( n33832,n28849,p3_instqueuerd_addr_reg_0_ );
   nand U36119 ( n35144,n35156,n35157 );
   nor U36120 ( n35157,n35158,n35159 );
   nor U36121 ( n35159,n33876,n34665 );
   nand U36122 ( n34665,n35154,n33834 );
   nor U36123 ( n35158,n33851,n34666 );
   nand U36124 ( n34666,n35155,n33870 );
   nor U36125 ( n35156,n35160,n35161 );
   nor U36126 ( n35161,n33849,n34669 );
   nand U36127 ( n34669,n35155,n33838 );
   nor U36128 ( n35160,n33872,n34670 );
   nand U36129 ( n34670,n35155,n33834 );
   nor U36130 ( n35155,n35162,n35163 );
   nor U36131 ( n35142,n35164,n35165 );
   nand U36132 ( n35165,n35166,n35167 );
   nor U36133 ( n35167,n35168,n35169 );
   nor U36134 ( n35169,n33830,n34653 );
   nand U36135 ( n34653,n35151,n33838 );
   nor U36136 ( n35168,n30650,n34654 );
   nand U36137 ( n34654,n35151,n33834 );
   nor U36138 ( n35166,n35170,n35171 );
   nor U36139 ( n35171,n33863,n34657 );
   nand U36140 ( n34657,n35154,n33870 );
   nor U36141 ( n35170,n33859,n34658 );
   nand U36142 ( n34658,n35154,n33838 );
   nor U36143 ( n35154,n35172,n35163 );
   not U36144 ( n35163,n35173 );
   nand U36145 ( n35164,n35174,n35175 );
   nor U36146 ( n35175,n35176,n35177 );
   nor U36147 ( n35177,n33845,n34643 );
   nand U36148 ( n34643,n35150,n33870 );
   nor U36149 ( n35176,n33839,n34644 );
   nand U36150 ( n34644,n35150,n33838 );
   nor U36151 ( n33838,n29368,p3_instqueuerd_addr_reg_0_ );
   nor U36152 ( n35174,n35178,n35179 );
   nor U36153 ( n35179,n33869,n34647 );
   nand U36154 ( n34647,n35150,n33834 );
   nor U36155 ( n33834,n29368,n29275 );
   not U36156 ( n29368,n28849 );
   nor U36157 ( n35150,n35172,n35173 );
   not U36158 ( n35172,n35162 );
   nor U36159 ( n35178,n33833,n34648 );
   nand U36160 ( n34648,n35151,n33870 );
   nor U36161 ( n33870,n29275,n28849 );
   nor U36162 ( n35151,n35173,n35162 );
   nor U36163 ( n35162,n35180,n35181 );
   nand U36164 ( n35173,n35182,n35183 );
   or U36165 ( n35183,n29254,n35180 );
   nor U36166 ( n35180,n29257,n34594 );
   nand U36167 ( n35182,n34627,n30802 );
   nand U36168 ( n34923,n35184,n35185 );
   nor U36169 ( n35185,n35186,n35187 );
   nand U36170 ( n35187,n35188,n35189 );
   nor U36171 ( n35189,n35190,n35191 );
   nor U36172 ( n35191,n33457,n35047 );
   nor U36173 ( n35190,n33465,n35048 );
   nor U36174 ( n35188,n35192,n35193 );
   nor U36175 ( n35193,n33433,n35043 );
   nor U36176 ( n35192,n33443,n35044 );
   nand U36177 ( n35186,n35194,n35195 );
   nor U36178 ( n35195,n35196,n35197 );
   nor U36179 ( n35197,n33473,n35037 );
   nor U36180 ( n35196,n33447,n35038 );
   nor U36181 ( n35194,n35198,n35199 );
   nor U36182 ( n35199,n33449,n35033 );
   nor U36183 ( n35198,n33477,n35034 );
   nor U36184 ( n35184,n35200,n35201 );
   nand U36185 ( n35201,n35202,n35203 );
   nor U36186 ( n35203,n35204,n35205 );
   nor U36187 ( n35205,n33459,n35025 );
   nor U36188 ( n35204,n33463,n35026 );
   nor U36189 ( n35202,n35206,n35207 );
   nor U36190 ( n35207,n33479,n35021 );
   nor U36191 ( n35206,n33427,n35022 );
   nand U36192 ( n35200,n35208,n35209 );
   nor U36193 ( n35209,n35210,n35211 );
   nor U36194 ( n35211,n33429,n35015 );
   nor U36195 ( n35210,n33471,n35016 );
   nor U36196 ( n35208,n35212,n35213 );
   nor U36197 ( n35213,n33435,n35011 );
   nor U36198 ( n35212,n33441,n35012 );
   nor U36199 ( n35080,n34970,n34958 );
   not U36200 ( n34958,n34972 );
   nand U36201 ( n34972,n35214,n35215 );
   nor U36202 ( n35215,n35216,n35217 );
   nand U36203 ( n35217,n35218,n35219 );
   nor U36204 ( n35219,n35220,n35221 );
   nor U36205 ( n35221,n33630,n35047 );
   nor U36206 ( n35220,n33635,n35048 );
   nor U36207 ( n35218,n35222,n35223 );
   nor U36208 ( n35223,n33612,n35043 );
   nor U36209 ( n35222,n33619,n35044 );
   nand U36210 ( n35216,n35224,n35225 );
   nor U36211 ( n35225,n35226,n35227 );
   nor U36212 ( n35227,n33641,n35037 );
   nor U36213 ( n35226,n33622,n35038 );
   nor U36214 ( n35224,n35228,n35229 );
   nor U36215 ( n35229,n33623,n35033 );
   nor U36216 ( n35228,n33644,n35034 );
   nor U36217 ( n35214,n35230,n35231 );
   nand U36218 ( n35231,n35232,n35233 );
   nor U36219 ( n35233,n35234,n35235 );
   nor U36220 ( n35235,n33631,n35025 );
   nor U36221 ( n35234,n33634,n35026 );
   nor U36222 ( n35232,n35236,n35237 );
   nor U36223 ( n35237,n30694,n35021 );
   nor U36224 ( n35236,n33608,n35022 );
   nand U36225 ( n35230,n35238,n35239 );
   nor U36226 ( n35239,n35240,n35241 );
   nor U36227 ( n35241,n33609,n35015 );
   nor U36228 ( n35240,n33640,n35016 );
   nor U36229 ( n35238,n35242,n35243 );
   nor U36230 ( n35243,n33613,n35011 );
   nor U36231 ( n35242,n33618,n35012 );
   and U36232 ( n34970,n35244,n35245 );
   nor U36233 ( n35245,n35246,n35247 );
   nand U36234 ( n35247,n35248,n35249 );
   nor U36235 ( n35249,n35250,n35251 );
   nor U36236 ( n35251,n33674,n35047 );
   nor U36237 ( n35250,n33679,n35048 );
   nor U36238 ( n35248,n35252,n35253 );
   nor U36239 ( n35253,n33700,n35043 );
   nor U36240 ( n35252,n33687,n35044 );
   nand U36241 ( n35246,n35254,n35255 );
   nor U36242 ( n35255,n35256,n35257 );
   nor U36243 ( n35257,n33666,n35037 );
   nor U36244 ( n35256,n33690,n35038 );
   nor U36245 ( n35254,n35258,n35259 );
   nor U36246 ( n35259,n33691,n35033 );
   nor U36247 ( n35258,n33669,n35034 );
   nor U36248 ( n35244,n35260,n35261 );
   nand U36249 ( n35261,n35262,n35263 );
   nor U36250 ( n35263,n35264,n35265 );
   nor U36251 ( n35265,n33675,n35025 );
   nor U36252 ( n35264,n33678,n35026 );
   nor U36253 ( n35262,n35266,n35267 );
   nor U36254 ( n35267,n30683,n35021 );
   nor U36255 ( n35266,n33696,n35022 );
   nand U36256 ( n35260,n35268,n35269 );
   nor U36257 ( n35269,n35270,n35271 );
   nor U36258 ( n35271,n33697,n35015 );
   nor U36259 ( n35270,n33665,n35016 );
   nor U36260 ( n35268,n35272,n35273 );
   nor U36261 ( n35273,n33701,n35011 );
   nor U36262 ( n35272,n33686,n35012 );
   and U36263 ( n34992,n35274,n35275 );
   nor U36264 ( n35275,n35276,n35277 );
   nand U36265 ( n35277,n35278,n35279 );
   nor U36266 ( n35279,n35280,n35281 );
   nor U36267 ( n35281,n33798,n35047 );
   nand U36268 ( n35047,n35282,n35283 );
   nor U36269 ( n35280,n33803,n35048 );
   nand U36270 ( n35048,n35284,n35283 );
   nor U36271 ( n35278,n35285,n35286 );
   nor U36272 ( n35286,n33780,n35043 );
   nand U36273 ( n35043,n35287,n35282 );
   nor U36274 ( n35285,n33787,n35044 );
   nand U36275 ( n35044,n35287,n35284 );
   nand U36276 ( n35276,n35288,n35289 );
   nor U36277 ( n35289,n35290,n35291 );
   nor U36278 ( n35291,n33809,n35037 );
   nand U36279 ( n35037,n35292,n34594 );
   nor U36280 ( n35290,n33790,n35038 );
   nand U36281 ( n35038,n35292,n34619 );
   nor U36282 ( n35288,n35293,n35294 );
   nor U36283 ( n35294,n33791,n35033 );
   nand U36284 ( n35033,n35292,n34597 );
   nor U36285 ( n35292,n29257,n35287 );
   nor U36286 ( n35293,n33812,n35034 );
   nand U36287 ( n35034,n35181,n35283 );
   nor U36288 ( n35274,n35295,n35296 );
   nand U36289 ( n35296,n35297,n35298 );
   nor U36290 ( n35298,n35299,n35300 );
   nor U36291 ( n35300,n33799,n35025 );
   nand U36292 ( n35025,n35301,n35283 );
   nor U36293 ( n35299,n33802,n35026 );
   nand U36294 ( n35026,n35302,n35283 );
   nor U36295 ( n35297,n35303,n35304 );
   nor U36296 ( n35304,n30662,n35021 );
   nand U36297 ( n35021,n35305,n34594 );
   nor U36298 ( n35303,n33776,n35022 );
   nand U36299 ( n35022,n35305,n34619 );
   nand U36300 ( n35295,n35306,n35307 );
   nor U36301 ( n35307,n35308,n35309 );
   nor U36302 ( n35309,n33777,n35015 );
   nand U36303 ( n35015,n35305,n34597 );
   nor U36304 ( n35305,n35283,n29257 );
   nor U36305 ( n35308,n33808,n35016 );
   nand U36306 ( n35016,n35287,n35181 );
   nor U36307 ( n35306,n35310,n35311 );
   nor U36308 ( n35311,n33781,n35011 );
   nand U36309 ( n35011,n35287,n35301 );
   nor U36310 ( n35310,n33786,n35012 );
   nand U36311 ( n35012,n35287,n35302 );
   not U36312 ( n35287,n35283 );
   nand U36313 ( n35283,n29245,n35312 );
   nand U36314 ( n35312,p3_instqueuerd_addr_reg_3_,n29257 );
   not U36315 ( n29245,n34627 );
   nor U36316 ( n34233,n34241,n31809 );
   nor U36317 ( n34999,n35313,n35314 );
   nor U36318 ( n35314,p3_ebx_reg_30_,n35315 );
   nor U36319 ( n35313,n35316,n35317 );
   nand U36320 ( n35319,p3_ebx_reg_31_,n35320 );
   nand U36321 ( n35320,n35316,n35321 );
   nand U36322 ( n35321,n34245,n35317 );
   and U36323 ( n35316,n34998,n35322 );
   nand U36324 ( n35322,n34245,n34996 );
   and U36325 ( n34998,n34236,n35323 );
   nand U36326 ( n35323,n34245,n35324 );
   not U36327 ( n34236,n34241 );
   nand U36328 ( n35318,n35325,n35326 );
   nor U36329 ( n35325,n35317,n35315 );
   nand U36330 ( n35315,p3_ebx_reg_29_,n34997 );
   nor U36331 ( n34997,n35324,n28173 );
   not U36332 ( n34238,n34245 );
   nor U36333 ( n34245,n34241,n30646 );
   nand U36334 ( n34241,n31747,n35327 );
   nand U36335 ( n35327,n35328,n31874 );
   not U36336 ( n31874,n29359 );
   nor U36337 ( n29359,n29301,n35329 );
   nand U36338 ( n29301,n35330,n31809 );
   nor U36339 ( n35330,n29309,n31808 );
   nand U36340 ( n31808,n35331,n31779 );
   nor U36341 ( n31779,n30670,n34202 );
   nor U36342 ( n35331,n30691,n30702 );
   nand U36343 ( n35328,n31759,n29208 );
   nor U36344 ( n29208,n29247,n35329 );
   nand U36345 ( n29247,n35332,n35333 );
   nor U36346 ( n35333,n31778,n35334 );
   nand U36347 ( n35334,n29309,n30646 );
   nor U36348 ( n35332,n30702,n31886 );
   nand U36349 ( n31886,n34202,n30670 );
   nand U36350 ( n35324,n35335,p3_ebx_reg_28_ );
   nor U36351 ( n35335,n34976,n35336 );
   nand U36352 ( n34976,n35337,p3_ebx_reg_26_ );
   nor U36353 ( n35337,n34953,n35338 );
   nand U36354 ( n34953,n35339,p3_ebx_reg_24_ );
   nor U36355 ( n35339,n34927,n35340 );
   nand U36356 ( n34927,n35341,p3_ebx_reg_22_ );
   nor U36357 ( n35341,n34878,n35342 );
   nand U36358 ( n34878,n35343,p3_ebx_reg_20_ );
   nor U36359 ( n35343,n34801,n35344 );
   nand U36360 ( n34801,n35345,p3_ebx_reg_18_ );
   nor U36361 ( n35345,n34724,n35346 );
   nand U36362 ( n34724,n35347,p3_ebx_reg_16_ );
   nor U36363 ( n35347,n34631,n35348 );
   nand U36364 ( n34631,n35349,p3_ebx_reg_14_ );
   nor U36365 ( n35349,n34541,n35350 );
   nand U36366 ( n34541,n35351,p3_ebx_reg_12_ );
   nor U36367 ( n35351,n34464,n35352 );
   nand U36368 ( n34464,n35353,p3_ebx_reg_10_ );
   nor U36369 ( n35353,n34387,n35354 );
   nand U36370 ( n34387,n35355,p3_ebx_reg_8_ );
   nor U36371 ( n35355,n34294,n35356 );
   nand U36372 ( n34294,n35357,p3_ebx_reg_6_ );
   nor U36373 ( n35357,n34277,n35358 );
   nand U36374 ( n34277,n35359,p3_ebx_reg_4_ );
   nor U36375 ( n35359,n34260,n35360 );
   nand U36376 ( n34260,p3_ebx_reg_2_,n34251 );
   nor U36377 ( n34251,n35361,n34237 );
   nor U36378 ( n35363,n35364,n35365 );
   nor U36379 ( n35365,n35366,n28823 );
   not U36380 ( n28823,p3_reip_reg_0_ );
   nor U36381 ( n35366,n35367,n35368 );
   nor U36382 ( n35364,n35369,n34237 );
   nor U36383 ( n35369,n35370,n35371 );
   nor U36384 ( n35362,n35372,n35373 );
   and U36385 ( n35373,n29275,n35374 );
   nor U36386 ( n35372,n35375,n31931 );
   nor U36387 ( n35375,n35376,n35377 );
   nand U36388 ( n35377,n35378,n35379 );
   nor U36389 ( n35381,n35382,n35383 );
   nand U36390 ( n35383,n35384,n35385 );
   nand U36391 ( n35385,n35370,n34244 );
   xor U36392 ( n34244,p3_ebx_reg_1_,p3_ebx_reg_0_ );
   nand U36393 ( n35384,n35374,n28849 );
   nor U36394 ( n28849,n29294,n34594 );
   nor U36395 ( n35382,n35361,n35386 );
   not U36396 ( n35361,p3_ebx_reg_1_ );
   nor U36397 ( n35380,n35387,n35388 );
   nand U36398 ( n35388,n35389,n35390 );
   nand U36399 ( n35389,n35367,p3_reip_reg_1_ );
   nand U36400 ( n35387,n35391,n35392 );
   nand U36401 ( n35392,p3_phyaddrpointer_reg_1_,n35393 );
   nand U36402 ( n35393,n35379,n35394 );
   nand U36403 ( n35394,n35395,p3_phyaddrpointer_reg_0_ );
   nand U36404 ( n35391,n35396,n31947 );
   nand U36405 ( n35396,n28242,n35398 );
   nand U36406 ( n35398,n35395,n31931 );
   not U36407 ( n31931,p3_phyaddrpointer_reg_0_ );
   nor U36408 ( n35400,n35401,n35402 );
   nand U36409 ( n35402,n35403,n35404 );
   nand U36410 ( n35404,n35374,n28862 );
   not U36411 ( n28862,n33871 );
   nor U36412 ( n33871,n35405,n35284 );
   nor U36413 ( n35405,n29257,n29294 );
   or U36414 ( n35403,n35397,n31966 );
   nand U36415 ( n35401,n35406,n35407 );
   nand U36416 ( n35407,n35408,n28333 );
   nor U36417 ( n35408,n35409,n35410 );
   nor U36418 ( n35410,n35411,n31966 );
   nand U36419 ( n35406,n35412,n28090 );
   nor U36420 ( n35412,n35413,n35414 );
   nor U36421 ( n35414,n35415,n34253 );
   not U36422 ( n34253,p3_ebx_reg_2_ );
   nor U36423 ( n35415,p3_ebx_reg_1_,p3_ebx_reg_0_ );
   nor U36424 ( n35399,n35416,n35417 );
   nand U36425 ( n35417,n35418,n35419 );
   nand U36426 ( n35419,n35420,p3_phyaddrpointer_reg_2_ );
   nand U36427 ( n35418,n28339,p3_ebx_reg_2_ );
   nand U36428 ( n35416,n35421,n35422 );
   nand U36429 ( n35422,p3_reip_reg_2_,n35423 );
   nand U36430 ( n35421,n35424,n29059 );
   nor U36431 ( n35424,n28264,n29064 );
   nor U36432 ( n35427,n35428,n35429 );
   nand U36433 ( n35429,n35430,n35431 );
   nand U36434 ( n35431,n35432,n35374 );
   nor U36435 ( n35432,n35433,n35434 );
   nor U36436 ( n35434,n35282,p3_instqueuerd_addr_reg_3_ );
   nand U36437 ( n35430,n35435,n28333 );
   xor U36438 ( n35435,n35436,n32005 );
   nor U36439 ( n35428,n35437,n28242 );
   not U36440 ( n35437,n32005 );
   nor U36441 ( n35426,n35438,n35439 );
   nand U36442 ( n35439,n35440,n35441 );
   nand U36443 ( n35441,n35420,p3_phyaddrpointer_reg_3_ );
   nor U36444 ( n35440,n35442,n35443 );
   nor U36445 ( n35443,p3_ebx_reg_3_,n35444 );
   nand U36446 ( n35444,n35370,n35445 );
   nor U36447 ( n35442,n35446,n35360 );
   not U36448 ( n35360,p3_ebx_reg_3_ );
   nor U36449 ( n35446,n35447,n35371 );
   nor U36450 ( n35447,n35448,n35445 );
   nand U36451 ( n35438,n35449,n35450 );
   nand U36452 ( n35450,p3_reip_reg_3_,n35451 );
   nand U36453 ( n35451,n35452,n35453 );
   nand U36454 ( n35453,n28380,n29059 );
   not U36455 ( n35452,n35423 );
   nand U36456 ( n35423,n35454,n35390 );
   nand U36457 ( n35390,n28379,n29064 );
   nand U36458 ( n35449,n35455,n29054 );
   nor U36459 ( n35455,n29059,n35456 );
   nand U36460 ( n35456,p3_reip_reg_1_,n28380 );
   not U36461 ( n29059,p3_reip_reg_2_ );
   nor U36462 ( n35458,n35459,n35460 );
   nand U36463 ( n35460,n35461,n35462 );
   nand U36464 ( n35462,n35463,n28090 );
   nor U36465 ( n35463,n35464,n35465 );
   nor U36466 ( n35465,n35466,n34269 );
   not U36467 ( n34269,p3_ebx_reg_4_ );
   nor U36468 ( n35466,p3_ebx_reg_3_,n35445 );
   nand U36469 ( n35461,n35374,n35467 );
   nand U36470 ( n35467,n29197,n35468 );
   nor U36471 ( n35374,n35469,n35470 );
   nand U36472 ( n35459,n35471,n35472 );
   nand U36473 ( n35471,n35473,n35395 );
   nor U36474 ( n35473,n35474,n35475 );
   nor U36475 ( n35475,n35476,n35477 );
   nor U36476 ( n35476,n32005,n35436 );
   nor U36477 ( n35457,n35478,n35479 );
   nand U36478 ( n35479,n35480,n35481 );
   nand U36479 ( n35481,n28339,p3_ebx_reg_4_ );
   nor U36480 ( n35480,n35482,n35483 );
   nor U36481 ( n35483,p3_reip_reg_4_,n35484 );
   nand U36482 ( n35484,n35485,n35368 );
   nor U36483 ( n35482,n35486,n29049 );
   nand U36484 ( n35478,n35487,n35488 );
   nand U36485 ( n35488,n35376,n32036 );
   nand U36486 ( n35487,n28277,p3_phyaddrpointer_reg_4_ );
   nor U36487 ( n35490,n35491,n35492 );
   nand U36488 ( n35492,n35493,n35472 );
   nand U36489 ( n35493,n35494,n35395 );
   xor U36490 ( n35494,n35495,n32080 );
   nor U36491 ( n35491,n35496,n35397 );
   not U36492 ( n35496,n32080 );
   nor U36493 ( n35489,n35497,n35498 );
   nand U36494 ( n35498,n35499,n35500 );
   nand U36495 ( n35500,n35420,p3_phyaddrpointer_reg_5_ );
   nor U36496 ( n35499,n35501,n35502 );
   nor U36497 ( n35502,p3_ebx_reg_5_,n35503 );
   nand U36498 ( n35503,n35370,n35504 );
   nor U36499 ( n35501,n35505,n35358 );
   not U36500 ( n35358,p3_ebx_reg_5_ );
   nor U36501 ( n35505,n35506,n35371 );
   nor U36502 ( n35506,n35448,n35504 );
   nand U36503 ( n35497,n35507,n35508 );
   nand U36504 ( n35508,p3_reip_reg_5_,n35509 );
   nand U36505 ( n35509,n35486,n35510 );
   nand U36506 ( n35510,n28380,n29049 );
   and U36507 ( n35486,n35454,n35511 );
   nand U36508 ( n35511,n35512,n35368 );
   nand U36509 ( n35507,n35513,n29044 );
   nor U36510 ( n35513,n35512,n35514 );
   nand U36511 ( n35514,p3_reip_reg_4_,n28379 );
   nor U36512 ( n35516,n35517,n35518 );
   nand U36513 ( n35518,n35519,n35520 );
   nand U36514 ( n35520,n35521,n35370 );
   nor U36515 ( n35521,n35522,n35523 );
   nor U36516 ( n35523,n35524,n34286 );
   not U36517 ( n34286,p3_ebx_reg_6_ );
   nor U36518 ( n35524,p3_ebx_reg_5_,n35504 );
   nand U36519 ( n35519,n35376,n32105 );
   nand U36520 ( n35517,n35525,n35472 );
   nand U36521 ( n35525,n35526,n35395 );
   nor U36522 ( n35526,n35527,n35528 );
   nor U36523 ( n35528,n35529,n35530 );
   nor U36524 ( n35529,n32080,n35495 );
   nor U36525 ( n35515,n35531,n35532 );
   nand U36526 ( n35532,n35533,n35534 );
   nand U36527 ( n35534,n28277,p3_phyaddrpointer_reg_6_ );
   nand U36528 ( n35533,n28339,p3_ebx_reg_6_ );
   nand U36529 ( n35531,n35535,n35536 );
   nand U36530 ( n35536,p3_reip_reg_6_,n35537 );
   nand U36531 ( n35535,n35538,n29039 );
   nor U36532 ( n35538,n28264,n35539 );
   nor U36533 ( n35541,n35542,n35543 );
   nand U36534 ( n35543,n35544,n35472 );
   nand U36535 ( n35544,n35545,n35395 );
   xor U36536 ( n35545,n35546,n32136 );
   nor U36537 ( n35542,n35547,n35397 );
   not U36538 ( n35547,n32136 );
   nor U36539 ( n35540,n35548,n35549 );
   nand U36540 ( n35549,n35550,n35551 );
   nand U36541 ( n35551,n28277,p3_phyaddrpointer_reg_7_ );
   nor U36542 ( n35550,n35552,n35553 );
   nor U36543 ( n35553,p3_ebx_reg_7_,n35554 );
   nand U36544 ( n35554,n35370,n35555 );
   nor U36545 ( n35552,n35556,n35356 );
   not U36546 ( n35356,p3_ebx_reg_7_ );
   nor U36547 ( n35556,n35557,n35371 );
   nor U36548 ( n35557,n35448,n35555 );
   nand U36549 ( n35548,n35558,n35559 );
   nand U36550 ( n35559,p3_reip_reg_7_,n35560 );
   nand U36551 ( n35560,n35561,n35562 );
   nand U36552 ( n35562,n35368,n29039 );
   not U36553 ( n29039,p3_reip_reg_6_ );
   not U36554 ( n35561,n35537 );
   nand U36555 ( n35537,n35454,n35563 );
   nand U36556 ( n35563,n35539,n28380 );
   nand U36557 ( n35558,n35564,n29034 );
   not U36558 ( n29034,p3_reip_reg_7_ );
   nor U36559 ( n35564,n35539,n35565 );
   nand U36560 ( n35565,p3_reip_reg_6_,n35368 );
   nor U36561 ( n35567,n35568,n35569 );
   nand U36562 ( n35569,n35570,n35571 );
   nand U36563 ( n35571,n35572,n28090 );
   nor U36564 ( n35572,n35573,n35574 );
   nor U36565 ( n35574,n35575,n34349 );
   not U36566 ( n34349,p3_ebx_reg_8_ );
   nor U36567 ( n35575,p3_ebx_reg_7_,n35555 );
   nand U36568 ( n35570,n35376,n32161 );
   nand U36569 ( n35568,n35576,n35472 );
   nand U36570 ( n35576,n35577,n35395 );
   nor U36571 ( n35577,n35578,n35579 );
   nor U36572 ( n35579,n35580,n35581 );
   nor U36573 ( n35580,n32136,n35546 );
   nor U36574 ( n35566,n35582,n35583 );
   nand U36575 ( n35583,n35584,n35585 );
   nand U36576 ( n35585,n28277,p3_phyaddrpointer_reg_8_ );
   nand U36577 ( n35584,n28339,p3_ebx_reg_8_ );
   nand U36578 ( n35582,n35586,n35587 );
   nand U36579 ( n35587,p3_reip_reg_8_,n35588 );
   nand U36580 ( n35586,n35589,n29029 );
   nor U36581 ( n35589,n28264,n35590 );
   nor U36582 ( n35592,n35593,n35594 );
   nand U36583 ( n35594,n35595,n35472 );
   nand U36584 ( n35595,n35596,n35395 );
   xor U36585 ( n35596,n35597,n32185 );
   nor U36586 ( n35593,n35598,n28242 );
   not U36587 ( n35598,n32185 );
   nor U36588 ( n35591,n35599,n35600 );
   nand U36589 ( n35600,n35601,n35602 );
   nand U36590 ( n35602,n35420,p3_phyaddrpointer_reg_9_ );
   nor U36591 ( n35601,n35603,n35604 );
   nor U36592 ( n35604,p3_ebx_reg_9_,n35605 );
   nand U36593 ( n35605,n35370,n35606 );
   nor U36594 ( n35603,n35607,n35354 );
   not U36595 ( n35354,p3_ebx_reg_9_ );
   nor U36596 ( n35607,n35608,n35371 );
   nor U36597 ( n35608,n35448,n35606 );
   nand U36598 ( n35599,n35609,n35610 );
   nand U36599 ( n35610,p3_reip_reg_9_,n35611 );
   nand U36600 ( n35611,n35612,n35613 );
   nand U36601 ( n35613,n28380,n29029 );
   not U36602 ( n35612,n35588 );
   nand U36603 ( n35588,n35454,n35614 );
   nand U36604 ( n35614,n35590,n28379 );
   nand U36605 ( n35609,n35615,n29024 );
   nor U36606 ( n35615,n35590,n35616 );
   nand U36607 ( n35616,p3_reip_reg_8_,n28379 );
   not U36608 ( n35590,n35617 );
   nor U36609 ( n35619,n35620,n35621 );
   nand U36610 ( n35621,n35622,n35623 );
   nand U36611 ( n35623,n35624,n28090 );
   nor U36612 ( n35624,n35625,n35626 );
   nor U36613 ( n35626,n35627,n34426 );
   not U36614 ( n34426,p3_ebx_reg_10_ );
   nor U36615 ( n35627,p3_ebx_reg_9_,n35606 );
   nand U36616 ( n35622,n35376,n32212 );
   nand U36617 ( n35620,n35628,n35472 );
   nand U36618 ( n35628,n35629,n35395 );
   nor U36619 ( n35629,n35630,n35631 );
   nor U36620 ( n35631,n35632,n35633 );
   nor U36621 ( n35632,n32185,n35597 );
   nor U36622 ( n35618,n35634,n35635 );
   nand U36623 ( n35635,n35636,n35637 );
   nand U36624 ( n35637,n35420,p3_phyaddrpointer_reg_10_ );
   nand U36625 ( n35636,n28339,p3_ebx_reg_10_ );
   nand U36626 ( n35634,n35638,n35639 );
   nand U36627 ( n35639,p3_reip_reg_10_,n35640 );
   nand U36628 ( n35638,n35641,n29019 );
   nor U36629 ( n35641,n35425,n35642 );
   nor U36630 ( n35644,n35645,n35646 );
   nand U36631 ( n35646,n35647,n35472 );
   nand U36632 ( n35647,n35648,n35395 );
   xor U36633 ( n35648,n35649,n32241 );
   nor U36634 ( n35645,n35650,n28242 );
   not U36635 ( n35650,n32241 );
   nor U36636 ( n35643,n35651,n35652 );
   nand U36637 ( n35652,n35653,n35654 );
   nand U36638 ( n35654,n35420,p3_phyaddrpointer_reg_11_ );
   nor U36639 ( n35653,n35655,n35656 );
   nor U36640 ( n35656,p3_ebx_reg_11_,n35657 );
   nand U36641 ( n35657,n35370,n35658 );
   nor U36642 ( n35655,n35659,n35352 );
   not U36643 ( n35352,p3_ebx_reg_11_ );
   nor U36644 ( n35659,n35660,n35371 );
   nor U36645 ( n35660,n35448,n35658 );
   nand U36646 ( n35651,n35661,n35662 );
   nand U36647 ( n35662,p3_reip_reg_11_,n35663 );
   nand U36648 ( n35663,n35664,n35665 );
   nand U36649 ( n35665,n35368,n29019 );
   not U36650 ( n29019,p3_reip_reg_10_ );
   not U36651 ( n35664,n35640 );
   nand U36652 ( n35640,n35454,n35666 );
   nand U36653 ( n35666,n35642,n35368 );
   nand U36654 ( n35661,n35667,n29014 );
   not U36655 ( n29014,p3_reip_reg_11_ );
   nor U36656 ( n35667,n35642,n35668 );
   nand U36657 ( n35668,p3_reip_reg_10_,n35368 );
   nor U36658 ( n35670,n35671,n35672 );
   nand U36659 ( n35672,n35673,n35674 );
   nand U36660 ( n35674,n35675,n35370 );
   nor U36661 ( n35675,n35676,n35677 );
   nor U36662 ( n35677,n35678,n34503 );
   not U36663 ( n34503,p3_ebx_reg_12_ );
   nor U36664 ( n35678,p3_ebx_reg_11_,n35658 );
   nand U36665 ( n35673,n35376,n32268 );
   nand U36666 ( n35671,n35679,n35472 );
   nand U36667 ( n35679,n35680,n35395 );
   nor U36668 ( n35680,n35681,n35682 );
   nor U36669 ( n35682,n35683,n35684 );
   nor U36670 ( n35683,n32241,n35649 );
   nor U36671 ( n35669,n35685,n35686 );
   nand U36672 ( n35686,n35687,n35688 );
   nand U36673 ( n35688,n35420,p3_phyaddrpointer_reg_12_ );
   nand U36674 ( n35687,n28339,p3_ebx_reg_12_ );
   nand U36675 ( n35685,n35689,n35690 );
   nand U36676 ( n35690,p3_reip_reg_12_,n35691 );
   nand U36677 ( n35689,n35692,n29009 );
   nor U36678 ( n35692,n35425,n35693 );
   nor U36679 ( n35695,n35696,n35697 );
   nand U36680 ( n35697,n35698,n35472 );
   nand U36681 ( n35698,n35699,n35395 );
   xor U36682 ( n35699,n35700,n32293 );
   nor U36683 ( n35696,n35701,n35397 );
   not U36684 ( n35701,n32293 );
   nor U36685 ( n35694,n35702,n35703 );
   nand U36686 ( n35703,n35704,n35705 );
   nand U36687 ( n35705,n35420,p3_phyaddrpointer_reg_13_ );
   nor U36688 ( n35704,n35706,n35707 );
   nor U36689 ( n35707,p3_ebx_reg_13_,n35708 );
   nand U36690 ( n35708,n35370,n35709 );
   nor U36691 ( n35706,n35710,n35350 );
   not U36692 ( n35350,p3_ebx_reg_13_ );
   nor U36693 ( n35710,n35711,n35371 );
   nor U36694 ( n35711,n35448,n35709 );
   nand U36695 ( n35702,n35712,n35713 );
   or U36696 ( n35713,n29004,n35714 );
   nand U36697 ( n35712,n35715,n29004 );
   nor U36698 ( n35715,n35693,n35716 );
   nand U36699 ( n35716,p3_reip_reg_12_,n28380 );
   nor U36700 ( n35718,n35719,n35720 );
   nand U36701 ( n35720,n35721,n35722 );
   nand U36702 ( n35722,n35723,n35370 );
   nor U36703 ( n35723,n35724,n35725 );
   nor U36704 ( n35725,n35726,n34580 );
   not U36705 ( n34580,p3_ebx_reg_14_ );
   nor U36706 ( n35726,p3_ebx_reg_13_,n35709 );
   nand U36707 ( n35721,n35376,n35727 );
   nand U36708 ( n35719,n35728,n35472 );
   nand U36709 ( n35728,n35729,n35395 );
   nor U36710 ( n35729,n35730,n35731 );
   nor U36711 ( n35731,n35732,n32331 );
   nor U36712 ( n35732,n32293,n35700 );
   nor U36713 ( n35717,n35733,n35734 );
   nand U36714 ( n35734,n35735,n35736 );
   nand U36715 ( n35736,n35420,p3_phyaddrpointer_reg_14_ );
   nand U36716 ( n35735,n28339,p3_ebx_reg_14_ );
   nand U36717 ( n35733,n35737,n35738 );
   nand U36718 ( n35738,p3_reip_reg_14_,n35739 );
   nand U36719 ( n35737,n35740,n28999 );
   nor U36720 ( n35740,n35425,n35741 );
   nor U36721 ( n35743,n35744,n35745 );
   nand U36722 ( n35745,n35746,n35472 );
   nand U36723 ( n35746,n35747,n35395 );
   xor U36724 ( n35747,n35748,n35749 );
   nor U36725 ( n35744,n32369,n35397 );
   not U36726 ( n32369,n35749 );
   nor U36727 ( n35742,n35750,n35751 );
   nand U36728 ( n35751,n35752,n35753 );
   nand U36729 ( n35753,n35420,p3_phyaddrpointer_reg_15_ );
   nor U36730 ( n35752,n35754,n35755 );
   nor U36731 ( n35755,p3_ebx_reg_15_,n35756 );
   nand U36732 ( n35756,n35370,n35757 );
   nor U36733 ( n35754,n35758,n35348 );
   not U36734 ( n35348,p3_ebx_reg_15_ );
   nor U36735 ( n35758,n35759,n35371 );
   nor U36736 ( n35759,n35448,n35757 );
   nand U36737 ( n35750,n35760,n35761 );
   nand U36738 ( n35761,p3_reip_reg_15_,n35762 );
   nand U36739 ( n35762,n35763,n35764 );
   nand U36740 ( n35764,n28380,n28999 );
   not U36741 ( n28999,p3_reip_reg_14_ );
   not U36742 ( n35763,n35739 );
   nand U36743 ( n35739,n35714,n35765 );
   nand U36744 ( n35765,n28380,n29004 );
   nor U36745 ( n35714,n35691,n35766 );
   nor U36746 ( n35766,n35425,p3_reip_reg_12_ );
   nand U36747 ( n35691,n35454,n35767 );
   nand U36748 ( n35767,n35693,n28380 );
   not U36749 ( n35693,n35768 );
   nand U36750 ( n35760,n35769,n28994 );
   not U36751 ( n28994,p3_reip_reg_15_ );
   nor U36752 ( n35769,n35741,n35770 );
   nand U36753 ( n35770,p3_reip_reg_14_,n35368 );
   nor U36754 ( n35772,n35773,n35774 );
   nand U36755 ( n35774,n35775,n35776 );
   nand U36756 ( n35776,n35777,n28090 );
   nor U36757 ( n35777,n35778,n35779 );
   nor U36758 ( n35779,n35780,n34686 );
   not U36759 ( n34686,p3_ebx_reg_16_ );
   nor U36760 ( n35780,p3_ebx_reg_15_,n35757 );
   nand U36761 ( n35775,n35376,n35781 );
   nand U36762 ( n35773,n35782,n35472 );
   nand U36763 ( n35782,n35783,n35395 );
   nor U36764 ( n35783,n35784,n35785 );
   nor U36765 ( n35785,n35786,n32394 );
   nor U36766 ( n35786,n35749,n35748 );
   nor U36767 ( n35771,n35787,n35788 );
   nand U36768 ( n35788,n35789,n35790 );
   nand U36769 ( n35790,n35420,p3_phyaddrpointer_reg_16_ );
   nand U36770 ( n35789,n35371,p3_ebx_reg_16_ );
   nand U36771 ( n35787,n35791,n35792 );
   nand U36772 ( n35792,p3_reip_reg_16_,n35793 );
   nand U36773 ( n35791,n35794,n28989 );
   nor U36774 ( n35794,n35425,n35795 );
   nor U36775 ( n35797,n35798,n35799 );
   nand U36776 ( n35799,n35800,n35472 );
   nand U36777 ( n35800,n35801,n35395 );
   xor U36778 ( n35801,n32427,n35802 );
   and U36779 ( n35798,n32427,n35376 );
   nor U36780 ( n35796,n35803,n35804 );
   nand U36781 ( n35804,n35805,n35806 );
   nand U36782 ( n35806,n28277,p3_phyaddrpointer_reg_17_ );
   nor U36783 ( n35805,n35807,n35808 );
   nor U36784 ( n35808,p3_ebx_reg_17_,n35809 );
   nand U36785 ( n35809,n35370,n35810 );
   nor U36786 ( n35807,n35811,n35346 );
   not U36787 ( n35346,p3_ebx_reg_17_ );
   nor U36788 ( n35811,n35812,n35371 );
   nor U36789 ( n35812,n35448,n35810 );
   nand U36790 ( n35803,n35813,n35814 );
   nand U36791 ( n35814,p3_reip_reg_17_,n35815 );
   nand U36792 ( n35815,n35816,n35817 );
   nand U36793 ( n35817,n35368,n28989 );
   not U36794 ( n35816,n35793 );
   nand U36795 ( n35793,n35454,n35818 );
   nand U36796 ( n35818,n28379,n35795 );
   nand U36797 ( n35813,n35819,n28984 );
   nor U36798 ( n35819,n35795,n35820 );
   nand U36799 ( n35820,p3_reip_reg_16_,n28379 );
   not U36800 ( n35795,n35821 );
   nor U36801 ( n35823,n35824,n35825 );
   nand U36802 ( n35825,n35826,n35827 );
   nand U36803 ( n35827,n35828,n28090 );
   nor U36804 ( n35828,n35829,n35830 );
   nor U36805 ( n35830,n35831,n34763 );
   not U36806 ( n34763,p3_ebx_reg_18_ );
   nor U36807 ( n35831,p3_ebx_reg_17_,n35810 );
   nand U36808 ( n35826,n35376,n35832 );
   nand U36809 ( n35824,n35833,n35472 );
   nand U36810 ( n35833,n35834,n35395 );
   nor U36811 ( n35834,n35835,n35836 );
   nor U36812 ( n35836,n35837,n32462 );
   nor U36813 ( n35837,n32427,n35802 );
   nor U36814 ( n35822,n35838,n35839 );
   nand U36815 ( n35839,n35840,n35841 );
   nand U36816 ( n35841,n35420,p3_phyaddrpointer_reg_18_ );
   nand U36817 ( n35840,n28339,p3_ebx_reg_18_ );
   nand U36818 ( n35838,n35842,n35843 );
   nand U36819 ( n35843,p3_reip_reg_18_,n35844 );
   nand U36820 ( n35842,n35845,n28979 );
   nor U36821 ( n35845,n35425,n35846 );
   nor U36822 ( n35848,n35849,n35850 );
   nand U36823 ( n35850,n35851,n35472 );
   nand U36824 ( n35472,n28775,n35454 );
   nand U36825 ( n35851,n35852,n35395 );
   xor U36826 ( n35852,n35835,n32500 );
   nor U36827 ( n35849,n32500,n35397 );
   nor U36828 ( n35847,n35853,n35854 );
   nand U36829 ( n35854,n35855,n35856 );
   nand U36830 ( n35856,n35420,p3_phyaddrpointer_reg_19_ );
   nor U36831 ( n35855,n35857,n35858 );
   nor U36832 ( n35858,p3_ebx_reg_19_,n35859 );
   nand U36833 ( n35859,n35370,n35860 );
   nor U36834 ( n35857,n35861,n35344 );
   not U36835 ( n35344,p3_ebx_reg_19_ );
   nor U36836 ( n35861,n35862,n35371 );
   nor U36837 ( n35862,n35448,n35860 );
   nand U36838 ( n35853,n35863,n35864 );
   nand U36839 ( n35864,p3_reip_reg_19_,n35865 );
   nand U36840 ( n35865,n35866,n35867 );
   nand U36841 ( n35867,n28379,n28979 );
   not U36842 ( n28979,p3_reip_reg_18_ );
   not U36843 ( n35866,n35844 );
   nand U36844 ( n35844,n35454,n35868 );
   nand U36845 ( n35868,n35846,n28379 );
   nand U36846 ( n35863,n35869,n28974 );
   not U36847 ( n28974,p3_reip_reg_19_ );
   nor U36848 ( n35869,n35846,n35870 );
   nand U36849 ( n35870,p3_reip_reg_18_,n28380 );
   nor U36850 ( n35872,n35873,n35874 );
   nand U36851 ( n35874,n35875,n35876 );
   nand U36852 ( n35876,n35877,n35395 );
   nor U36853 ( n35877,n35878,n35879 );
   nor U36854 ( n35879,n35880,n32534 );
   and U36855 ( n35880,n32500,n35835 );
   nand U36856 ( n35875,n35881,n28090 );
   nor U36857 ( n35881,n35882,n35883 );
   nor U36858 ( n35883,n35884,n34840 );
   not U36859 ( n34840,p3_ebx_reg_20_ );
   nor U36860 ( n35884,p3_ebx_reg_19_,n35860 );
   nor U36861 ( n35873,n32534,n35397 );
   nor U36862 ( n35871,n35885,n35886 );
   nand U36863 ( n35886,n35887,n35888 );
   nand U36864 ( n35888,n35420,p3_phyaddrpointer_reg_20_ );
   nand U36865 ( n35887,n28339,p3_ebx_reg_20_ );
   nand U36866 ( n35885,n35889,n35890 );
   or U36867 ( n35890,n35891,p3_reip_reg_20_ );
   nand U36868 ( n35889,p3_reip_reg_20_,n35892 );
   nor U36869 ( n35894,n35895,n35896 );
   nand U36870 ( n35896,n35897,n35898 );
   nand U36871 ( n35898,n35899,n35395 );
   xor U36872 ( n35899,n35900,n32567 );
   nand U36873 ( n35897,n35376,n32567 );
   nor U36874 ( n35895,n32588,n35379 );
   nor U36875 ( n35893,n35901,n35902 );
   nand U36876 ( n35902,n35903,n35904 );
   nand U36877 ( n35904,p3_ebx_reg_21_,n35905 );
   nand U36878 ( n35905,n35386,n35906 );
   nand U36879 ( n35906,n35882,n35370 );
   nand U36880 ( n35903,n35907,n35342 );
   not U36881 ( n35342,p3_ebx_reg_21_ );
   nor U36882 ( n35907,n35882,n28260 );
   nand U36883 ( n35901,n35908,n35909 );
   nand U36884 ( n35909,p3_reip_reg_21_,n35910 );
   nand U36885 ( n35910,n35911,n35912 );
   nand U36886 ( n35912,n28379,n28969 );
   not U36887 ( n35911,n35892 );
   nand U36888 ( n35892,n35454,n35913 );
   or U36889 ( n35913,n35425,n35914 );
   nand U36890 ( n35908,n35915,n28964 );
   nor U36891 ( n35915,n28969,n35891 );
   nand U36892 ( n35891,n35914,n28380 );
   nor U36893 ( n35917,n35918,n35919 );
   nand U36894 ( n35919,n35920,n35921 );
   nand U36895 ( n35921,n35922,n35395 );
   nor U36896 ( n35922,n35923,n35924 );
   nor U36897 ( n35924,n35925,n32602 );
   nor U36898 ( n35925,n32567,n35900 );
   nand U36899 ( n35920,n35926,n28090 );
   nor U36900 ( n35926,n35927,n35928 );
   nor U36901 ( n35928,n35929,n34917 );
   not U36902 ( n34917,p3_ebx_reg_22_ );
   nor U36903 ( n35929,p3_ebx_reg_21_,n35930 );
   nor U36904 ( n35918,n32602,n35397 );
   nor U36905 ( n35916,n35931,n35932 );
   nand U36906 ( n35932,n35933,n35934 );
   nand U36907 ( n35934,n35420,p3_phyaddrpointer_reg_22_ );
   nand U36908 ( n35933,n28339,p3_ebx_reg_22_ );
   nand U36909 ( n35931,n35935,n35936 );
   nand U36910 ( n35936,n35937,n28959 );
   nand U36911 ( n35935,p3_reip_reg_22_,n35938 );
   nor U36912 ( n35940,n35941,n35942 );
   nand U36913 ( n35942,n35943,n35944 );
   nand U36914 ( n35944,n35945,n35395 );
   xor U36915 ( n35945,n35946,n32635 );
   nand U36916 ( n35943,n35376,n32635 );
   nor U36917 ( n35941,n32660,n35379 );
   nor U36918 ( n35939,n35947,n35948 );
   nand U36919 ( n35948,n35949,n35950 );
   nand U36920 ( n35950,p3_ebx_reg_23_,n35951 );
   nand U36921 ( n35951,n35386,n35952 );
   nand U36922 ( n35952,n35927,n35370 );
   nand U36923 ( n35949,n35953,n35340 );
   not U36924 ( n35340,p3_ebx_reg_23_ );
   nor U36925 ( n35953,n35927,n28260 );
   nand U36926 ( n35947,n35954,n35955 );
   nand U36927 ( n35955,p3_reip_reg_23_,n35956 );
   nand U36928 ( n35956,n35957,n35958 );
   nand U36929 ( n35958,n28379,n28959 );
   not U36930 ( n28959,p3_reip_reg_22_ );
   not U36931 ( n35957,n35938 );
   nand U36932 ( n35938,n35454,n35959 );
   nand U36933 ( n35959,n35960,n28380 );
   nand U36934 ( n35954,n35961,n28954 );
   not U36935 ( n28954,p3_reip_reg_23_ );
   and U36936 ( n35961,p3_reip_reg_22_,n35937 );
   nor U36937 ( n35937,n35960,n28264 );
   nor U36938 ( n35963,n35964,n35965 );
   nand U36939 ( n35965,n35966,n35967 );
   nand U36940 ( n35967,n35968,n28333 );
   nor U36941 ( n35968,n35969,n35970 );
   nor U36942 ( n35970,n35971,n32673 );
   nor U36943 ( n35971,n32635,n35946 );
   nand U36944 ( n35966,n35972,n28090 );
   nor U36945 ( n35972,n35973,n35974 );
   nor U36946 ( n35974,n35975,n34942 );
   not U36947 ( n34942,p3_ebx_reg_24_ );
   nor U36948 ( n35975,p3_ebx_reg_23_,n35976 );
   nor U36949 ( n35964,n32673,n35397 );
   nor U36950 ( n35962,n35977,n35978 );
   nand U36951 ( n35978,n35979,n35980 );
   nand U36952 ( n35980,n35420,p3_phyaddrpointer_reg_24_ );
   nand U36953 ( n35979,n28339,p3_ebx_reg_24_ );
   nand U36954 ( n35977,n35981,n35982 );
   or U36955 ( n35982,n35983,p3_reip_reg_24_ );
   nand U36956 ( n35981,p3_reip_reg_24_,n35984 );
   nor U36957 ( n35986,n35987,n35988 );
   nand U36958 ( n35988,n35989,n35990 );
   nand U36959 ( n35990,n35991,n28333 );
   xor U36960 ( n35991,n35992,n32711 );
   nand U36961 ( n35989,n35376,n32711 );
   nor U36962 ( n35987,n32724,n35379 );
   nor U36963 ( n35985,n35993,n35994 );
   nand U36964 ( n35994,n35995,n35996 );
   nand U36965 ( n35996,p3_ebx_reg_25_,n35997 );
   nand U36966 ( n35997,n35386,n35998 );
   nand U36967 ( n35998,n35973,n35370 );
   nand U36968 ( n35995,n35999,n35338 );
   not U36969 ( n35338,p3_ebx_reg_25_ );
   nor U36970 ( n35999,n35973,n28260 );
   nand U36971 ( n35993,n36000,n36001 );
   nand U36972 ( n36001,p3_reip_reg_25_,n36002 );
   nand U36973 ( n36002,n36003,n36004 );
   nand U36974 ( n36004,n35368,n28949 );
   not U36975 ( n36003,n35984 );
   nand U36976 ( n35984,n35454,n36005 );
   or U36977 ( n36005,n35425,n36006 );
   nand U36978 ( n36000,n36007,n28944 );
   nor U36979 ( n36007,n28949,n35983 );
   nand U36980 ( n35983,n36006,n35368 );
   nor U36981 ( n36009,n36010,n36011 );
   nand U36982 ( n36011,n36012,n36013 );
   nand U36983 ( n36013,n36014,n28333 );
   nor U36984 ( n36014,n36015,n36016 );
   nor U36985 ( n36016,n36017,n36018 );
   nor U36986 ( n36017,n32711,n35992 );
   nand U36987 ( n36012,n36019,n28090 );
   nor U36988 ( n36019,n36020,n36021 );
   nor U36989 ( n36021,n36022,n34964 );
   not U36990 ( n34964,p3_ebx_reg_26_ );
   nor U36991 ( n36022,p3_ebx_reg_25_,n36023 );
   nor U36992 ( n36010,n36018,n35397 );
   nor U36993 ( n36008,n36024,n36025 );
   nand U36994 ( n36025,n36026,n36027 );
   nand U36995 ( n36027,n28277,p3_phyaddrpointer_reg_26_ );
   nand U36996 ( n36026,n28339,p3_ebx_reg_26_ );
   nand U36997 ( n36024,n36028,n36029 );
   nand U36998 ( n36029,n36030,n28939 );
   nand U36999 ( n36028,p3_reip_reg_26_,n36031 );
   nor U37000 ( n36033,n36034,n36035 );
   nand U37001 ( n36035,n36036,n36037 );
   nand U37002 ( n36037,n36038,n28333 );
   xor U37003 ( n36038,n36039,n32774 );
   nand U37004 ( n36036,n35376,n32774 );
   nor U37005 ( n36034,n32795,n35379 );
   nor U37006 ( n36032,n36040,n36041 );
   nand U37007 ( n36041,n36042,n36043 );
   nand U37008 ( n36043,p3_ebx_reg_27_,n36044 );
   nand U37009 ( n36044,n35386,n36045 );
   nand U37010 ( n36045,n36020,n35370 );
   nand U37011 ( n36042,n36046,n35336 );
   not U37012 ( n35336,p3_ebx_reg_27_ );
   nor U37013 ( n36046,n36020,n28260 );
   nand U37014 ( n36040,n36047,n36048 );
   nand U37015 ( n36048,p3_reip_reg_27_,n36049 );
   nand U37016 ( n36049,n36050,n36051 );
   nand U37017 ( n36051,n28380,n28939 );
   not U37018 ( n28939,p3_reip_reg_26_ );
   not U37019 ( n36050,n36031 );
   nand U37020 ( n36031,n35454,n36052 );
   nand U37021 ( n36052,n36053,n28380 );
   nand U37022 ( n36047,n36054,n28934 );
   not U37023 ( n28934,p3_reip_reg_27_ );
   and U37024 ( n36054,p3_reip_reg_26_,n36030 );
   nor U37025 ( n36030,n36053,n28264 );
   nor U37026 ( n36056,n36057,n36058 );
   nand U37027 ( n36058,n36059,n36060 );
   nand U37028 ( n36060,n36061,n28090 );
   nor U37029 ( n36061,n36062,n36063 );
   nor U37030 ( n36063,n36064,n34987 );
   not U37031 ( n34987,p3_ebx_reg_28_ );
   nor U37032 ( n36064,p3_ebx_reg_27_,n36065 );
   nand U37033 ( n36059,n36066,n28333 );
   nor U37034 ( n36066,n36067,n36068 );
   nor U37035 ( n36068,n36069,n36070 );
   nor U37036 ( n36069,n32774,n36039 );
   nor U37037 ( n36057,n36070,n35397 );
   nor U37038 ( n36055,n36071,n36072 );
   nand U37039 ( n36072,n36073,n36074 );
   nand U37040 ( n36074,n28277,p3_phyaddrpointer_reg_28_ );
   nand U37041 ( n36073,n35371,p3_ebx_reg_28_ );
   nand U37042 ( n36071,n36075,n36076 );
   or U37043 ( n36076,n36077,p3_reip_reg_28_ );
   nand U37044 ( n36075,p3_reip_reg_28_,n36078 );
   nor U37045 ( n36080,n36081,n36082 );
   nand U37046 ( n36082,n36083,n36084 );
   nand U37047 ( n36084,n36085,n28333 );
   nor U37048 ( n36085,n36086,n36087 );
   nor U37049 ( n36087,n36067,n32846 );
   nand U37050 ( n36083,n36088,n35370 );
   nor U37051 ( n36088,n36089,n36090 );
   nor U37052 ( n36090,n36062,n34996 );
   nor U37053 ( n36081,n32846,n35397 );
   nor U37054 ( n36079,n36091,n36092 );
   nand U37055 ( n36092,n36093,n36094 );
   nand U37056 ( n36094,n28277,p3_phyaddrpointer_reg_29_ );
   nand U37057 ( n36093,n35371,p3_ebx_reg_29_ );
   not U37058 ( n35371,n35386 );
   nand U37059 ( n36091,n36095,n36096 );
   nand U37060 ( n36096,p3_reip_reg_29_,n36097 );
   nand U37061 ( n36097,n36098,n36099 );
   nand U37062 ( n36099,n28379,n28929 );
   not U37063 ( n36098,n36078 );
   nand U37064 ( n36078,n35454,n36100 );
   or U37065 ( n36100,n35425,n36101 );
   nand U37066 ( n36095,n36102,n28924 );
   nor U37067 ( n36102,n28929,n36077 );
   nand U37068 ( n36077,n36101,n28379 );
   nor U37069 ( n36104,n36105,n36106 );
   nand U37070 ( n36106,n36107,n36108 );
   nand U37071 ( n36108,n36109,n28333 );
   not U37072 ( n35395,n35378 );
   xor U37073 ( n36109,n32873,n36086 );
   nand U37074 ( n36107,n35376,n36110 );
   not U37075 ( n35376,n35397 );
   nand U37076 ( n35397,n36111,n33055 );
   nor U37077 ( n36111,n35367,n28856 );
   nor U37078 ( n36105,n32879,n35379 );
   nor U37079 ( n36103,n36112,n36113 );
   nand U37080 ( n36113,n36114,n36115 );
   nand U37081 ( n36115,p3_ebx_reg_30_,n36116 );
   nand U37082 ( n36116,n35386,n36117 );
   nand U37083 ( n36117,n36089,n28090 );
   not U37084 ( n35370,n35448 );
   nand U37085 ( n36114,n36118,n35317 );
   not U37086 ( n35317,p3_ebx_reg_30_ );
   nor U37087 ( n36118,n36089,n28260 );
   nand U37088 ( n36112,n36119,n36120 );
   nand U37089 ( n36120,p3_reip_reg_30_,n36121 );
   nand U37090 ( n36119,n36122,n28919 );
   nor U37091 ( n36122,n35425,n36123 );
   not U37092 ( n35425,n28379 );
   nor U37093 ( n36125,n36126,n36127 );
   nand U37094 ( n36127,n36128,n36129 );
   nand U37095 ( n36129,n36130,n36086 );
   and U37096 ( n36086,n36067,n32846 );
   nand U37097 ( n32846,n36131,n36132 );
   nand U37098 ( n36132,n33064,n32862 );
   and U37099 ( n36067,n36133,n36015 );
   not U37100 ( n36015,n36039 );
   nand U37101 ( n36039,n36134,n35969 );
   not U37102 ( n35969,n35992 );
   nand U37103 ( n35992,n36135,n35923 );
   not U37104 ( n35923,n35946 );
   nand U37105 ( n35946,n36136,n35878 );
   not U37106 ( n35878,n35900 );
   nand U37107 ( n35900,n36137,n35835 );
   and U37108 ( n35835,n36138,n35784 );
   not U37109 ( n35784,n35802 );
   nand U37110 ( n35802,n36139,n35730 );
   not U37111 ( n35730,n35748 );
   nand U37112 ( n35748,n36140,n35681 );
   not U37113 ( n35681,n35700 );
   nand U37114 ( n35700,n36141,n35630 );
   not U37115 ( n35630,n35649 );
   nand U37116 ( n35649,n36142,n35578 );
   not U37117 ( n35578,n35597 );
   nand U37118 ( n35597,n36143,n35527 );
   not U37119 ( n35527,n35546 );
   nand U37120 ( n35546,n36144,n35474 );
   not U37121 ( n35474,n35495 );
   nand U37122 ( n35495,n36145,n35409 );
   not U37123 ( n35409,n35436 );
   nand U37124 ( n35436,n35411,n31966 );
   xor U37125 ( n31966,n31947,p3_phyaddrpointer_reg_2_ );
   nor U37126 ( n35411,p3_phyaddrpointer_reg_0_,n31947 );
   nor U37127 ( n36145,n32036,n32005 );
   xor U37128 ( n32005,n32011,n36146 );
   nand U37129 ( n36146,p3_phyaddrpointer_reg_2_,p3_phyaddrpointer_reg_1_ );
   not U37130 ( n32036,n35477 );
   nand U37131 ( n35477,n36147,n36148 );
   nand U37132 ( n36147,n32039,n36149 );
   nand U37133 ( n36149,n32043,p3_phyaddrpointer_reg_1_ );
   not U37134 ( n32039,p3_phyaddrpointer_reg_4_ );
   nor U37135 ( n36144,n32105,n32080 );
   xor U37136 ( n32080,p3_phyaddrpointer_reg_5_,n36150 );
   not U37137 ( n32105,n35530 );
   nand U37138 ( n35530,n36151,n36152 );
   nand U37139 ( n36151,n32115,n36153 );
   nand U37140 ( n36153,n36150,p3_phyaddrpointer_reg_5_ );
   not U37141 ( n32115,p3_phyaddrpointer_reg_6_ );
   nor U37142 ( n36143,n32161,n32136 );
   xor U37143 ( n32136,n32141,n36152 );
   not U37144 ( n32161,n35581 );
   nand U37145 ( n35581,n36154,n36155 );
   nand U37146 ( n36154,n32165,n36156 );
   or U37147 ( n36156,n36152,n32141 );
   not U37148 ( n32165,p3_phyaddrpointer_reg_8_ );
   nor U37149 ( n36142,n32212,n32185 );
   xor U37150 ( n32185,n32190,n36155 );
   not U37151 ( n32212,n35633 );
   nand U37152 ( n35633,n36157,n32278 );
   nand U37153 ( n36157,n32222,n36158 );
   or U37154 ( n36158,n36155,n32190 );
   not U37155 ( n32222,p3_phyaddrpointer_reg_10_ );
   nor U37156 ( n36141,n32268,n32241 );
   xor U37157 ( n32241,n32246,n32278 );
   not U37158 ( n32268,n35684 );
   nand U37159 ( n35684,n32356,n36159 );
   nand U37160 ( n36159,n36160,n32282 );
   not U37161 ( n32356,n32351 );
   nor U37162 ( n36140,n35727,n32293 );
   xor U37163 ( n32293,p3_phyaddrpointer_reg_13_,n32351 );
   not U37164 ( n35727,n32331 );
   nand U37165 ( n32331,n32419,n36161 );
   nand U37166 ( n36161,n36162,n32353 );
   nor U37167 ( n36139,n35781,n35749 );
   xor U37168 ( n35749,p3_phyaddrpointer_reg_15_,n32414 );
   not U37169 ( n35781,n32394 );
   nand U37170 ( n32394,n36163,n36164 );
   nand U37171 ( n36163,n32416,n36165 );
   nand U37172 ( n36165,n32414,p3_phyaddrpointer_reg_15_ );
   not U37173 ( n32416,p3_phyaddrpointer_reg_16_ );
   nor U37174 ( n36138,n35832,n32427 );
   xor U37175 ( n32427,n32450,n36164 );
   not U37176 ( n35832,n32462 );
   nand U37177 ( n32462,n36166,n36167 );
   or U37178 ( n36166,p3_phyaddrpointer_reg_18_,n32473 );
   and U37179 ( n36137,n32534,n32500 );
   xor U37180 ( n32500,p3_phyaddrpointer_reg_19_,n36167 );
   nand U37181 ( n32534,n36168,n36169 );
   or U37182 ( n36169,n32545,p3_phyaddrpointer_reg_20_ );
   nor U37183 ( n36136,n36170,n32567 );
   xor U37184 ( n32567,n32588,n36168 );
   not U37185 ( n36170,n32602 );
   nand U37186 ( n32602,n36171,n36172 );
   or U37187 ( n36172,n32613,p3_phyaddrpointer_reg_22_ );
   nor U37188 ( n36135,n36173,n32635 );
   xor U37189 ( n32635,n32660,n36171 );
   not U37190 ( n36173,n32673 );
   nand U37191 ( n32673,n36174,n36175 );
   or U37192 ( n36175,n32684,p3_phyaddrpointer_reg_24_ );
   nor U37193 ( n36134,n32752,n32711 );
   xor U37194 ( n32711,n32724,n36174 );
   not U37195 ( n32752,n36018 );
   nand U37196 ( n36018,n36176,n36177 );
   or U37197 ( n36177,n32761,p3_phyaddrpointer_reg_26_ );
   nor U37198 ( n36133,n32823,n32774 );
   xor U37199 ( n32774,n32795,n36176 );
   not U37200 ( n32823,n36070 );
   nand U37201 ( n36070,n33064,n36178 );
   or U37202 ( n36178,n32832,p3_phyaddrpointer_reg_28_ );
   nor U37203 ( n36130,n36110,n35378 );
   nand U37204 ( n35378,n36179,p3_state2_reg_1_ );
   nor U37205 ( n36179,n35367,n33055 );
   xor U37206 ( n33055,p3_phyaddrpointer_reg_31_,n36180 );
   not U37207 ( n36110,n32873 );
   nand U37208 ( n32873,n36180,n36181 );
   nand U37209 ( n36181,n36131,n32879 );
   not U37210 ( n32879,p3_phyaddrpointer_reg_30_ );
   not U37211 ( n36131,n33087 );
   nand U37212 ( n36180,p3_phyaddrpointer_reg_30_,n33087 );
   nor U37213 ( n33087,n32862,n33064 );
   nand U37214 ( n33064,p3_phyaddrpointer_reg_28_,n32832 );
   nor U37215 ( n32832,n36176,n32795 );
   not U37216 ( n32795,p3_phyaddrpointer_reg_27_ );
   nand U37217 ( n36176,p3_phyaddrpointer_reg_26_,n32761 );
   nor U37218 ( n32761,n36174,n32724 );
   not U37219 ( n32724,p3_phyaddrpointer_reg_25_ );
   nand U37220 ( n36174,p3_phyaddrpointer_reg_24_,n32684 );
   nor U37221 ( n32684,n36171,n32660 );
   not U37222 ( n32660,p3_phyaddrpointer_reg_23_ );
   nand U37223 ( n36171,p3_phyaddrpointer_reg_22_,n32613 );
   nor U37224 ( n32613,n36168,n32588 );
   not U37225 ( n32588,p3_phyaddrpointer_reg_21_ );
   nand U37226 ( n36168,p3_phyaddrpointer_reg_20_,n32545 );
   nor U37227 ( n32545,n36167,n32511 );
   not U37228 ( n32511,p3_phyaddrpointer_reg_19_ );
   nand U37229 ( n36167,p3_phyaddrpointer_reg_18_,n32473 );
   nor U37230 ( n32473,n36164,n32450 );
   not U37231 ( n32450,p3_phyaddrpointer_reg_17_ );
   nand U37232 ( n36164,n36182,p3_phyaddrpointer_reg_16_ );
   nor U37233 ( n36182,n32380,n32419 );
   not U37234 ( n32419,n32414 );
   nor U37235 ( n32414,n32353,n36162 );
   nand U37236 ( n36162,n32351,p3_phyaddrpointer_reg_13_ );
   nor U37237 ( n32351,n32282,n36160 );
   or U37238 ( n36160,n32278,n32246 );
   not U37239 ( n32246,p3_phyaddrpointer_reg_11_ );
   nand U37240 ( n32278,n36183,p3_phyaddrpointer_reg_10_ );
   nor U37241 ( n36183,n32190,n36155 );
   nand U37242 ( n36155,n36184,p3_phyaddrpointer_reg_8_ );
   nor U37243 ( n36184,n32141,n36152 );
   nand U37244 ( n36152,n36185,p3_phyaddrpointer_reg_6_ );
   nor U37245 ( n36185,n32085,n36148 );
   not U37246 ( n36148,n36150 );
   nor U37247 ( n36150,n32086,n31947 );
   not U37248 ( n31947,p3_phyaddrpointer_reg_1_ );
   nand U37249 ( n32086,p3_phyaddrpointer_reg_4_,n32043 );
   nor U37250 ( n32043,n32011,n32012 );
   not U37251 ( n32012,p3_phyaddrpointer_reg_2_ );
   not U37252 ( n32011,p3_phyaddrpointer_reg_3_ );
   not U37253 ( n32085,p3_phyaddrpointer_reg_5_ );
   not U37254 ( n32141,p3_phyaddrpointer_reg_7_ );
   not U37255 ( n32190,p3_phyaddrpointer_reg_9_ );
   not U37256 ( n32282,p3_phyaddrpointer_reg_12_ );
   not U37257 ( n32353,p3_phyaddrpointer_reg_14_ );
   not U37258 ( n32380,p3_phyaddrpointer_reg_15_ );
   not U37259 ( n32862,p3_phyaddrpointer_reg_29_ );
   nand U37260 ( n36128,n36186,n36089 );
   and U37261 ( n36089,n36062,n34996 );
   not U37262 ( n34996,p3_ebx_reg_29_ );
   and U37263 ( n36062,n36187,n36020 );
   not U37264 ( n36020,n36065 );
   nand U37265 ( n36065,n36188,n35973 );
   not U37266 ( n35973,n36023 );
   nand U37267 ( n36023,n36189,n35927 );
   not U37268 ( n35927,n35976 );
   nand U37269 ( n35976,n36190,n35882 );
   not U37270 ( n35882,n35930 );
   nand U37271 ( n35930,n36191,n35829 );
   not U37272 ( n35829,n35860 );
   nand U37273 ( n35860,n36192,n35778 );
   not U37274 ( n35778,n35810 );
   nand U37275 ( n35810,n36193,n35724 );
   not U37276 ( n35724,n35757 );
   nand U37277 ( n35757,n36194,n35676 );
   not U37278 ( n35676,n35709 );
   nand U37279 ( n35709,n36195,n35625 );
   not U37280 ( n35625,n35658 );
   nand U37281 ( n35658,n36196,n35573 );
   not U37282 ( n35573,n35606 );
   nand U37283 ( n35606,n36197,n35522 );
   not U37284 ( n35522,n35555 );
   nand U37285 ( n35555,n36198,n35464 );
   not U37286 ( n35464,n35504 );
   nand U37287 ( n35504,n36199,n35413 );
   not U37288 ( n35413,n35445 );
   nand U37289 ( n35445,n36200,n34237 );
   not U37290 ( n34237,p3_ebx_reg_0_ );
   nor U37291 ( n36200,p3_ebx_reg_2_,p3_ebx_reg_1_ );
   nor U37292 ( n36199,p3_ebx_reg_4_,p3_ebx_reg_3_ );
   nor U37293 ( n36198,p3_ebx_reg_6_,p3_ebx_reg_5_ );
   nor U37294 ( n36197,p3_ebx_reg_8_,p3_ebx_reg_7_ );
   nor U37295 ( n36196,p3_ebx_reg_9_,p3_ebx_reg_10_ );
   nor U37296 ( n36195,p3_ebx_reg_12_,p3_ebx_reg_11_ );
   nor U37297 ( n36194,p3_ebx_reg_14_,p3_ebx_reg_13_ );
   nor U37298 ( n36193,p3_ebx_reg_16_,p3_ebx_reg_15_ );
   nor U37299 ( n36192,p3_ebx_reg_18_,p3_ebx_reg_17_ );
   nor U37300 ( n36191,p3_ebx_reg_20_,p3_ebx_reg_19_ );
   nor U37301 ( n36190,p3_ebx_reg_22_,p3_ebx_reg_21_ );
   nor U37302 ( n36189,p3_ebx_reg_24_,p3_ebx_reg_23_ );
   nor U37303 ( n36188,p3_ebx_reg_26_,p3_ebx_reg_25_ );
   nor U37304 ( n36187,p3_ebx_reg_28_,p3_ebx_reg_27_ );
   nor U37305 ( n36186,p3_ebx_reg_30_,n28260 );
   nand U37306 ( n35448,n36201,n36202 );
   nor U37307 ( n36202,n36203,n35329 );
   not U37308 ( n35329,n29314 );
   nor U37309 ( n36201,n35326,n35469 );
   not U37310 ( n35469,n36204 );
   nor U37311 ( n36126,n33069,n35379 );
   not U37312 ( n35379,n35420 );
   nor U37313 ( n35420,n30726,n35367 );
   not U37314 ( n30726,p3_state2_reg_3_ );
   not U37315 ( n33069,p3_phyaddrpointer_reg_31_ );
   nor U37316 ( n36124,n36205,n36206 );
   nand U37317 ( n36206,n36207,n36208 );
   nand U37318 ( n36208,p3_reip_reg_31_,n36209 );
   nand U37319 ( n36209,n36210,n36211 );
   nand U37320 ( n36211,n35368,n28919 );
   not U37321 ( n28919,p3_reip_reg_30_ );
   not U37322 ( n36210,n36121 );
   nand U37323 ( n36121,n35454,n36212 );
   nand U37324 ( n36212,n36123,n35368 );
   nand U37325 ( n36207,n36213,n28917 );
   not U37326 ( n28917,p3_reip_reg_31_ );
   nor U37327 ( n36213,n36123,n36214 );
   nand U37328 ( n36214,p3_reip_reg_30_,n28379 );
   nand U37329 ( n35368,n36215,n36216 );
   nand U37330 ( n36216,n36217,n36204 );
   nor U37331 ( n36217,n28804,n29186 );
   not U37332 ( n28804,n31857 );
   nand U37333 ( n36215,n36218,n36204 );
   and U37334 ( n36218,n29314,n36203 );
   nand U37335 ( n36123,n36219,n36101 );
   nor U37336 ( n36101,n36220,n36053 );
   nand U37337 ( n36053,n36221,n36006 );
   nor U37338 ( n36006,n36222,n35960 );
   nand U37339 ( n35960,n36223,n35914 );
   nor U37340 ( n35914,n36224,n35846 );
   nand U37341 ( n35846,n36225,n35821 );
   nor U37342 ( n35821,n36226,n35741 );
   nand U37343 ( n35741,n36227,n35768 );
   nor U37344 ( n35768,n36228,n35642 );
   nand U37345 ( n35642,n36229,n35617 );
   nor U37346 ( n35617,n36230,n35539 );
   nand U37347 ( n35539,n36231,n35485 );
   not U37348 ( n35485,n35512 );
   nand U37349 ( n35512,n36232,p3_reip_reg_2_ );
   nor U37350 ( n36232,n29064,n29054 );
   not U37351 ( n29054,p3_reip_reg_3_ );
   nor U37352 ( n36231,n29044,n29049 );
   not U37353 ( n29049,p3_reip_reg_4_ );
   not U37354 ( n29044,p3_reip_reg_5_ );
   nand U37355 ( n36230,p3_reip_reg_7_,p3_reip_reg_6_ );
   nor U37356 ( n36229,n29024,n29029 );
   not U37357 ( n29029,p3_reip_reg_8_ );
   not U37358 ( n29024,p3_reip_reg_9_ );
   nand U37359 ( n36228,p3_reip_reg_11_,p3_reip_reg_10_ );
   nor U37360 ( n36227,n29004,n29009 );
   not U37361 ( n29009,p3_reip_reg_12_ );
   not U37362 ( n29004,p3_reip_reg_13_ );
   nand U37363 ( n36226,p3_reip_reg_15_,p3_reip_reg_14_ );
   nor U37364 ( n36225,n28984,n28989 );
   not U37365 ( n28989,p3_reip_reg_16_ );
   not U37366 ( n28984,p3_reip_reg_17_ );
   nand U37367 ( n36224,p3_reip_reg_19_,p3_reip_reg_18_ );
   nor U37368 ( n36223,n28964,n28969 );
   not U37369 ( n28969,p3_reip_reg_20_ );
   not U37370 ( n28964,p3_reip_reg_21_ );
   nand U37371 ( n36222,p3_reip_reg_23_,p3_reip_reg_22_ );
   nor U37372 ( n36221,n28944,n28949 );
   not U37373 ( n28949,p3_reip_reg_24_ );
   not U37374 ( n28944,p3_reip_reg_25_ );
   nand U37375 ( n36220,p3_reip_reg_27_,p3_reip_reg_26_ );
   nor U37376 ( n36219,n28924,n28929 );
   not U37377 ( n28929,p3_reip_reg_28_ );
   not U37378 ( n28924,p3_reip_reg_29_ );
   nor U37379 ( n36205,n35326,n35386 );
   nand U37380 ( n35386,n36204,n36233 );
   nand U37381 ( n36233,n36234,n36235 );
   nand U37382 ( n36235,n36236,n29314 );
   nor U37383 ( n36236,p3_ebx_reg_31_,n36203 );
   nand U37384 ( n36234,n31857,n29186 );
   nand U37385 ( n29186,n36203,n28809 );
   not U37386 ( n28809,n28805 );
   nor U37387 ( n36203,n28801,p3_statebs16_reg );
   nor U37388 ( n36204,n28808,n35367 );
   not U37389 ( n35367,n35454 );
   nand U37390 ( n35454,n36237,n36238 );
   nor U37391 ( n36238,n29153,n29167 );
   nor U37392 ( n29167,n36239,n28796 );
   nand U37393 ( n28796,n28856,n28808 );
   nand U37394 ( n36239,p3_state2_reg_0_,p3_state2_reg_3_ );
   and U37395 ( n29153,n36240,n29149 );
   nor U37396 ( n29149,n28856,p3_state2_reg_2_ );
   nor U37397 ( n36240,p3_statebs16_reg,p3_state2_reg_0_ );
   nor U37398 ( n36237,n28776,n36241 );
   and U37399 ( n36241,n28790,n28775 );
   not U37400 ( n28790,p3_state2_reg_0_ );
   and U37401 ( n28776,n31747,n36242 );
   nand U37402 ( n36242,n36243,n29374 );
   nand U37403 ( n29374,n29224,n36244 );
   nand U37404 ( n36244,n29187,n29352 );
   nand U37405 ( n29352,n36245,n31847 );
   nand U37406 ( n29187,n31857,n29349 );
   or U37407 ( n36243,n29211,n34230 );
   nor U37408 ( n34230,n28878,n29222 );
   not U37409 ( n29222,n33245 );
   nand U37410 ( n33245,n29314,n29349 );
   nor U37411 ( n29349,n36246,n30702 );
   not U37412 ( n28878,n29260 );
   nand U37413 ( n29260,n36245,n29315 );
   nor U37414 ( n36245,n29308,n31771 );
   not U37415 ( n28808,p3_state2_reg_2_ );
   not U37416 ( n35326,p3_ebx_reg_31_ );
   nor U37417 ( n36247,n36249,n36250 );
   nor U37418 ( n36250,n28822,n36251 );
   or U37419 ( n36251,p3_datawidth_reg_1_,p3_reip_reg_1_ );
   and U37420 ( n36249,n28822,p3_byteenable_reg_3_ );
   nand U37421 ( n36253,p3_byteenable_reg_1_,n28822 );
   and U37422 ( n36252,n36248,n28819 );
   not U37423 ( n28819,n28826 );
   nor U37424 ( n28826,n29064,n28822 );
   not U37425 ( n29064,p3_reip_reg_1_ );
   nand U37426 ( n36248,n36254,n36255 );
   nor U37427 ( n36255,p3_reip_reg_0_,p3_datawidth_reg_1_ );
   nor U37428 ( n36254,p3_datawidth_reg_0_,n28822 );
   nand U37429 ( n28822,n36256,n36257 );
   nor U37430 ( n36257,n36258,n36259 );
   nand U37431 ( n36259,n36260,n36261 );
   nor U37432 ( n36261,n36262,n36263 );
   nand U37433 ( n36263,n29139,n29140 );
   not U37434 ( n29140,p3_datawidth_reg_29_ );
   not U37435 ( n29139,p3_datawidth_reg_28_ );
   nand U37436 ( n36262,n29113,n29141 );
   not U37437 ( n29141,p3_datawidth_reg_30_ );
   not U37438 ( n29113,p3_datawidth_reg_2_ );
   nor U37439 ( n36260,n36264,n36265 );
   nand U37440 ( n36265,n29135,n29136 );
   not U37441 ( n29136,p3_datawidth_reg_25_ );
   not U37442 ( n29135,p3_datawidth_reg_24_ );
   nand U37443 ( n36264,n29137,n29138 );
   not U37444 ( n29138,p3_datawidth_reg_27_ );
   not U37445 ( n29137,p3_datawidth_reg_26_ );
   nand U37446 ( n36258,n36266,n36267 );
   nor U37447 ( n36267,n36268,n36269 );
   nand U37448 ( n36269,n29117,n29118 );
   not U37449 ( n29118,p3_datawidth_reg_7_ );
   not U37450 ( n29117,p3_datawidth_reg_6_ );
   nand U37451 ( n36268,n29119,n29120 );
   not U37452 ( n29120,p3_datawidth_reg_9_ );
   not U37453 ( n29119,p3_datawidth_reg_8_ );
   nor U37454 ( n36266,n36270,n36271 );
   nand U37455 ( n36271,n29142,n29114 );
   not U37456 ( n29114,p3_datawidth_reg_3_ );
   not U37457 ( n29142,p3_datawidth_reg_31_ );
   nand U37458 ( n36270,n29115,n29116 );
   not U37459 ( n29116,p3_datawidth_reg_5_ );
   not U37460 ( n29115,p3_datawidth_reg_4_ );
   nor U37461 ( n36256,n36272,n36273 );
   nand U37462 ( n36273,n36274,n36275 );
   nor U37463 ( n36275,n36276,n36277 );
   nand U37464 ( n36277,n29123,n29124 );
   not U37465 ( n29124,p3_datawidth_reg_13_ );
   not U37466 ( n29123,p3_datawidth_reg_12_ );
   nand U37467 ( n36276,n29125,n29126 );
   not U37468 ( n29126,p3_datawidth_reg_15_ );
   not U37469 ( n29125,p3_datawidth_reg_14_ );
   nor U37470 ( n36274,n36278,n36279 );
   nand U37471 ( n36279,n29121,n29122 );
   not U37472 ( n29122,p3_datawidth_reg_11_ );
   not U37473 ( n29121,p3_datawidth_reg_10_ );
   and U37474 ( n36278,p3_datawidth_reg_0_,p3_datawidth_reg_1_ );
   nand U37475 ( n36272,n36280,n36281 );
   nor U37476 ( n36281,n36282,n36283 );
   nand U37477 ( n36283,n29131,n29132 );
   not U37478 ( n29132,p3_datawidth_reg_21_ );
   not U37479 ( n29131,p3_datawidth_reg_20_ );
   nand U37480 ( n36282,n29133,n29134 );
   not U37481 ( n29134,p3_datawidth_reg_23_ );
   not U37482 ( n29133,p3_datawidth_reg_22_ );
   nor U37483 ( n36280,n36284,n36285 );
   nand U37484 ( n36285,n29127,n29128 );
   not U37485 ( n29128,p3_datawidth_reg_17_ );
   not U37486 ( n29127,p3_datawidth_reg_16_ );
   nand U37487 ( n36284,n29129,n29130 );
   not U37488 ( n29130,p3_datawidth_reg_19_ );
   not U37489 ( n29129,p3_datawidth_reg_18_ );
   nand U37490 ( n36286,p3_flush_reg,n28813 );
   nand U37491 ( n28813,n31747,n29200 );
   nand U37492 ( n29200,n36287,n36288 );
   nor U37493 ( n36287,n31763,n36289 );
   nor U37494 ( n36289,n30702,n31764 );
   nand U37495 ( n31764,n28794,n36290 );
   nand U37496 ( n36290,n29304,n28805 );
   and U37497 ( n31763,n36291,n36292 );
   nand U37498 ( n36292,n29366,n28805 );
   nand U37499 ( n28805,n36293,n36294 );
   nand U37500 ( n36294,p3_state_reg_2_,p3_state_reg_1_ );
   nor U37501 ( n36293,p3_state_reg_0_,n28903 );
   nor U37502 ( n36291,n29308,n28801 );
   not U37503 ( n28801,n28794 );
   nand U37504 ( n28794,ready22_reg,ready2 );
   nand U37505 ( n33089,n31747,n29227 );
   nand U37506 ( n29227,n36295,n36296 );
   nand U37507 ( n36296,n31759,n29214 );
   and U37508 ( n29214,n29365,n31857 );
   nor U37509 ( n31857,n29366,n28771 );
   not U37510 ( n31759,n29209 );
   nand U37511 ( n29209,n36297,n36298 );
   nand U37512 ( n36298,n36299,n36300 );
   nand U37513 ( n36300,n36301,n36302 );
   nand U37514 ( n36302,n36303,n36304 );
   not U37515 ( n36299,n36305 );
   nand U37516 ( n36295,n31757,n29215 );
   not U37517 ( n29215,n31695 );
   nand U37518 ( n31695,n29365,n29314 );
   nor U37519 ( n29314,n29304,n28771 );
   and U37520 ( n29365,n36306,n36307 );
   nor U37521 ( n36307,n29309,n36308 );
   nand U37522 ( n36308,n30691,n30646 );
   nor U37523 ( n36306,n31848,n30702 );
   not U37524 ( n31848,n31760 );
   not U37525 ( n31757,n29216 );
   nand U37526 ( n29216,n29224,n36309 );
   nand U37527 ( n36309,n36310,n36303 );
   nor U37528 ( n36303,n36311,n36312 );
   nor U37529 ( n36312,n30775,p3_instqueuerd_addr_reg_0_ );
   not U37530 ( n30775,p3_instqueuewr_addr_reg_0_ );
   nor U37531 ( n36313,n36315,n36316 );
   nor U37532 ( n36316,n28806,n28157 );
   not U37533 ( n28897,n28895 );
   not U37534 ( n28806,p3_statebs16_reg );
   nor U37535 ( n36315,n28895,n28898 );
   nand U37536 ( n36314,n28903,n29077 );
   not U37537 ( n29077,p3_state_reg_0_ );
   nor U37538 ( n28903,p3_state_reg_1_,p3_state_reg_2_ );
   nor U37539 ( n36317,n36318,n36319 );
   and U37540 ( n36319,n28780,p3_d_c_n_reg );
   nor U37541 ( n36318,p3_codefetch_reg,n28780 );
   not U37542 ( n28780,n28781 );
   nor U37543 ( n28781,n29074,p3_state_reg_0_ );
   nand U37544 ( n36321,p3_codefetch_reg,n36322 );
   nand U37545 ( n36322,n36288,n31747 );
   nor U37546 ( n31747,n29181,p3_state2_reg_1_ );
   nand U37547 ( n29181,p3_state2_reg_2_,p3_state2_reg_0_ );
   and U37548 ( n36288,n36323,n36324 );
   nand U37549 ( n36324,n29308,n36325 );
   nand U37550 ( n36325,n36326,n29224 );
   nor U37551 ( n36326,n28771,n36246 );
   nand U37552 ( n36246,n36327,n31862 );
   nor U37553 ( n31862,n31809,n31778 );
   not U37554 ( n31778,n30691 );
   nor U37555 ( n36327,n31841,n30670 );
   nand U37556 ( n31841,n34202,n31777 );
   not U37557 ( n31777,n29309 );
   not U37558 ( n28771,n29350 );
   not U37559 ( n29308,n30702 );
   nand U37560 ( n36323,n36328,n30702 );
   nand U37561 ( n30702,n36329,n36330 );
   nor U37562 ( n36330,n36331,n36332 );
   nand U37563 ( n36332,n36333,n36334 );
   nor U37564 ( n36334,n36335,n36336 );
   nor U37565 ( n36336,n36337,n33567 );
   not U37566 ( n33567,p3_instqueue_reg_14__2_ );
   nor U37567 ( n36335,n36338,n33564 );
   not U37568 ( n33564,p3_instqueue_reg_13__2_ );
   nor U37569 ( n36333,n36339,n36340 );
   nor U37570 ( n36340,n36341,n33558 );
   not U37571 ( n33558,p3_instqueue_reg_12__2_ );
   nor U37572 ( n36339,n36342,n33575 );
   not U37573 ( n33575,p3_instqueue_reg_6__2_ );
   nand U37574 ( n36331,n36343,n36344 );
   nor U37575 ( n36344,n36345,n36346 );
   nor U37576 ( n36346,n36347,n33590 );
   not U37577 ( n33590,p3_instqueue_reg_5__2_ );
   nor U37578 ( n36345,n36348,n33554 );
   not U37579 ( n33554,p3_instqueue_reg_4__2_ );
   nor U37580 ( n36343,n36349,n36350 );
   nor U37581 ( n36350,n36351,n33586 );
   not U37582 ( n33586,p3_instqueue_reg_2__2_ );
   nor U37583 ( n36349,n36352,n33585 );
   not U37584 ( n33585,p3_instqueue_reg_1__2_ );
   nor U37585 ( n36329,n36353,n36354 );
   nand U37586 ( n36354,n36355,n36356 );
   nor U37587 ( n36356,n36357,n36358 );
   nor U37588 ( n36358,n36359,n30705 );
   not U37589 ( n30705,p3_instqueue_reg_0__2_ );
   nor U37590 ( n36357,n36360,n33580 );
   not U37591 ( n33580,p3_instqueue_reg_10__2_ );
   nor U37592 ( n36355,n36361,n36362 );
   nor U37593 ( n36362,n36363,n33555 );
   not U37594 ( n33555,p3_instqueue_reg_8__2_ );
   nor U37595 ( n36361,n33877,n33576 );
   not U37596 ( n33576,p3_instqueue_reg_7__2_ );
   nand U37597 ( n36353,n36364,n36365 );
   nor U37598 ( n36365,n36366,n36367 );
   nor U37599 ( n36367,n36368,n33589 );
   not U37600 ( n33589,p3_instqueue_reg_3__2_ );
   nor U37601 ( n36366,n35468,n33568 );
   not U37602 ( n33568,p3_instqueue_reg_15__2_ );
   nor U37603 ( n36364,n36369,n36370 );
   nor U37604 ( n36370,n36371,n33563 );
   not U37605 ( n33563,p3_instqueue_reg_11__2_ );
   nor U37606 ( n36369,n36372,n33579 );
   not U37607 ( n33579,p3_instqueue_reg_9__2_ );
   nand U37608 ( n36328,n36373,n29224 );
   not U37609 ( n29224,n29211 );
   nand U37610 ( n29211,n36374,n36297 );
   nand U37611 ( n36297,n36375,n36376 );
   nand U37612 ( n36376,p3_instqueuewr_addr_reg_4_,n36377 );
   nand U37613 ( n36377,p3_instqueuerd_addr_reg_4_,n36378 );
   or U37614 ( n36375,n36378,p3_instqueuerd_addr_reg_4_ );
   nand U37615 ( n36374,n36310,n36379 );
   xor U37616 ( n36379,n36304,n36311 );
   xor U37617 ( n36304,p3_instqueuerd_addr_reg_1_,n29316 );
   nor U37618 ( n36310,n36301,n36305 );
   nand U37619 ( n36305,n36380,n36381 );
   xor U37620 ( n36381,n36382,n36378 );
   nand U37621 ( n36378,n36383,n36384 );
   nand U37622 ( n36384,n36385,n29235 );
   not U37623 ( n29235,p3_instqueuewr_addr_reg_3_ );
   or U37624 ( n36385,n36386,p3_instqueuerd_addr_reg_3_ );
   nand U37625 ( n36383,p3_instqueuerd_addr_reg_3_,n36386 );
   nand U37626 ( n36382,p3_instqueuewr_addr_reg_4_,n29197 );
   not U37627 ( n29197,p3_instqueuerd_addr_reg_4_ );
   xor U37628 ( n36380,n36387,n36386 );
   nand U37629 ( n36386,n36388,n36389 );
   nand U37630 ( n36389,n36390,n29278 );
   or U37631 ( n36390,n36391,p3_instqueuerd_addr_reg_2_ );
   nand U37632 ( n36388,p3_instqueuerd_addr_reg_2_,n36391 );
   xor U37633 ( n36387,n29254,p3_instqueuewr_addr_reg_3_ );
   xor U37634 ( n36301,n36392,n36391 );
   nand U37635 ( n36391,n36393,n36394 );
   nand U37636 ( n36394,n36395,n29316 );
   not U37637 ( n29316,p3_instqueuewr_addr_reg_1_ );
   or U37638 ( n36395,p3_instqueuerd_addr_reg_1_,n36311 );
   nand U37639 ( n36393,p3_instqueuerd_addr_reg_1_,n36311 );
   nor U37640 ( n36311,n29275,p3_instqueuewr_addr_reg_0_ );
   xor U37641 ( n36392,n29278,n29257 );
   not U37642 ( n29278,p3_instqueuewr_addr_reg_2_ );
   nor U37643 ( n36373,n35470,n31771 );
   or U37644 ( n31771,n31877,n31809 );
   not U37645 ( n31809,n30646 );
   nand U37646 ( n30646,n36396,n36397 );
   nor U37647 ( n36397,n36398,n36399 );
   nand U37648 ( n36399,n36400,n36401 );
   nor U37649 ( n36401,n36402,n36403 );
   nor U37650 ( n36403,n36337,n33863 );
   not U37651 ( n33863,p3_instqueue_reg_14__7_ );
   nor U37652 ( n36402,n36338,n33859 );
   not U37653 ( n33859,p3_instqueue_reg_13__7_ );
   nor U37654 ( n36400,n36404,n36405 );
   nor U37655 ( n36405,n36341,n33876 );
   not U37656 ( n33876,p3_instqueue_reg_12__7_ );
   nor U37657 ( n36404,n36342,n33845 );
   not U37658 ( n33845,p3_instqueue_reg_6__7_ );
   nand U37659 ( n36398,n36406,n36407 );
   nor U37660 ( n36407,n36408,n36409 );
   nor U37661 ( n36409,n36347,n33839 );
   not U37662 ( n33839,p3_instqueue_reg_5__7_ );
   nor U37663 ( n36408,n36348,n33869 );
   not U37664 ( n33869,p3_instqueue_reg_4__7_ );
   nor U37665 ( n36406,n36410,n36411 );
   nor U37666 ( n36411,n36351,n33833 );
   not U37667 ( n33833,p3_instqueue_reg_2__7_ );
   nor U37668 ( n36410,n36352,n33830 );
   not U37669 ( n33830,p3_instqueue_reg_1__7_ );
   nor U37670 ( n36396,n36412,n36413 );
   nand U37671 ( n36413,n36414,n36415 );
   nor U37672 ( n36415,n36416,n36417 );
   nor U37673 ( n36417,n36359,n30650 );
   not U37674 ( n30650,p3_instqueue_reg_0__7_ );
   nor U37675 ( n36416,n36360,n33851 );
   not U37676 ( n33851,p3_instqueue_reg_10__7_ );
   nor U37677 ( n36414,n36418,n36419 );
   nor U37678 ( n36419,n36363,n33872 );
   not U37679 ( n33872,p3_instqueue_reg_8__7_ );
   nor U37680 ( n36418,n33877,n33846 );
   not U37681 ( n33846,p3_instqueue_reg_7__7_ );
   nand U37682 ( n36412,n36420,n36421 );
   nor U37683 ( n36421,n36422,n36423 );
   nor U37684 ( n36423,n36368,n33837 );
   not U37685 ( n33837,p3_instqueue_reg_3__7_ );
   nor U37686 ( n36422,n35468,n33864 );
   not U37687 ( n33864,p3_instqueue_reg_15__7_ );
   nor U37688 ( n36420,n36424,n36425 );
   nor U37689 ( n36425,n36371,n33858 );
   not U37690 ( n33858,p3_instqueue_reg_11__7_ );
   nor U37691 ( n36424,n36372,n33849 );
   not U37692 ( n33849,p3_instqueue_reg_9__7_ );
   nand U37693 ( n31877,n36426,n31760 );
   nor U37694 ( n31760,n34202,n31837 );
   not U37695 ( n31837,n30670 );
   nand U37696 ( n30670,n36427,n36428 );
   nor U37697 ( n36428,n36429,n36430 );
   nand U37698 ( n36430,n36431,n36432 );
   nor U37699 ( n36432,n36433,n36434 );
   nor U37700 ( n36434,n36337,n33732 );
   not U37701 ( n33732,p3_instqueue_reg_14__5_ );
   nor U37702 ( n36433,n36338,n33729 );
   not U37703 ( n33729,p3_instqueue_reg_13__5_ );
   nor U37704 ( n36431,n36435,n36436 );
   nor U37705 ( n36436,n36341,n33723 );
   not U37706 ( n33723,p3_instqueue_reg_12__5_ );
   nor U37707 ( n36435,n36342,n33740 );
   not U37708 ( n33740,p3_instqueue_reg_6__5_ );
   nand U37709 ( n36429,n36437,n36438 );
   nor U37710 ( n36438,n36439,n36440 );
   nor U37711 ( n36440,n36347,n33755 );
   not U37712 ( n33755,p3_instqueue_reg_5__5_ );
   nor U37713 ( n36439,n36348,n33719 );
   not U37714 ( n33719,p3_instqueue_reg_4__5_ );
   nor U37715 ( n36437,n36441,n36442 );
   nor U37716 ( n36442,n36351,n33751 );
   not U37717 ( n33751,p3_instqueue_reg_2__5_ );
   nor U37718 ( n36441,n36352,n33750 );
   not U37719 ( n33750,p3_instqueue_reg_1__5_ );
   nor U37720 ( n36427,n36443,n36444 );
   nand U37721 ( n36444,n36445,n36446 );
   nor U37722 ( n36446,n36447,n36448 );
   nor U37723 ( n36448,n36359,n30673 );
   not U37724 ( n30673,p3_instqueue_reg_0__5_ );
   nor U37725 ( n36447,n36360,n33745 );
   not U37726 ( n33745,p3_instqueue_reg_10__5_ );
   nor U37727 ( n36445,n36449,n36450 );
   nor U37728 ( n36450,n36363,n33720 );
   not U37729 ( n33720,p3_instqueue_reg_8__5_ );
   nor U37730 ( n36449,n33877,n33741 );
   not U37731 ( n33741,p3_instqueue_reg_7__5_ );
   nand U37732 ( n36443,n36451,n36452 );
   nor U37733 ( n36452,n36453,n36454 );
   nor U37734 ( n36454,n36368,n33754 );
   not U37735 ( n33754,p3_instqueue_reg_3__5_ );
   nor U37736 ( n36453,n35468,n33733 );
   not U37737 ( n33733,p3_instqueue_reg_15__5_ );
   nor U37738 ( n36451,n36455,n36456 );
   nor U37739 ( n36456,n36371,n33728 );
   not U37740 ( n33728,p3_instqueue_reg_11__5_ );
   nor U37741 ( n36455,n36372,n33744 );
   not U37742 ( n33744,p3_instqueue_reg_9__5_ );
   not U37743 ( n34202,n30659 );
   nand U37744 ( n30659,n36457,n36458 );
   nor U37745 ( n36458,n36459,n36460 );
   nand U37746 ( n36460,n36461,n36462 );
   nor U37747 ( n36462,n36463,n36464 );
   nor U37748 ( n36464,n36337,n33802 );
   not U37749 ( n33802,p3_instqueue_reg_14__6_ );
   nor U37750 ( n36463,n36338,n33799 );
   not U37751 ( n33799,p3_instqueue_reg_13__6_ );
   nor U37752 ( n36461,n36465,n36466 );
   nor U37753 ( n36466,n36341,n33812 );
   not U37754 ( n33812,p3_instqueue_reg_12__6_ );
   nor U37755 ( n36465,n36342,n33786 );
   not U37756 ( n33786,p3_instqueue_reg_6__6_ );
   nand U37757 ( n36459,n36467,n36468 );
   nor U37758 ( n36468,n36469,n36470 );
   nor U37759 ( n36470,n36347,n33781 );
   not U37760 ( n33781,p3_instqueue_reg_5__6_ );
   nor U37761 ( n36469,n36348,n33808 );
   not U37762 ( n33808,p3_instqueue_reg_4__6_ );
   nor U37763 ( n36467,n36471,n36472 );
   nor U37764 ( n36472,n36351,n33777 );
   not U37765 ( n33777,p3_instqueue_reg_2__6_ );
   nor U37766 ( n36471,n36352,n33776 );
   not U37767 ( n33776,p3_instqueue_reg_1__6_ );
   nor U37768 ( n36457,n36473,n36474 );
   nand U37769 ( n36474,n36475,n36476 );
   nor U37770 ( n36476,n36477,n36478 );
   nor U37771 ( n36478,n36359,n30662 );
   not U37772 ( n30662,p3_instqueue_reg_0__6_ );
   nor U37773 ( n36477,n36360,n33791 );
   not U37774 ( n33791,p3_instqueue_reg_10__6_ );
   nor U37775 ( n36475,n36479,n36480 );
   nor U37776 ( n36480,n36363,n33809 );
   not U37777 ( n33809,p3_instqueue_reg_8__6_ );
   nor U37778 ( n36479,n33877,n33787 );
   not U37779 ( n33787,p3_instqueue_reg_7__6_ );
   nand U37780 ( n36473,n36481,n36482 );
   nor U37781 ( n36482,n36483,n36484 );
   nor U37782 ( n36484,n36368,n33780 );
   not U37783 ( n33780,p3_instqueue_reg_3__6_ );
   nor U37784 ( n36483,n35468,n33803 );
   not U37785 ( n33803,p3_instqueue_reg_15__6_ );
   nor U37786 ( n36481,n36485,n36486 );
   nor U37787 ( n36486,n36371,n33798 );
   not U37788 ( n33798,p3_instqueue_reg_11__6_ );
   nor U37789 ( n36485,n36372,n33790 );
   not U37790 ( n33790,p3_instqueue_reg_9__6_ );
   nor U37791 ( n36426,n30691,n29309 );
   nand U37792 ( n29309,n36487,n36488 );
   nor U37793 ( n36488,n36489,n36490 );
   nand U37794 ( n36490,n36491,n36492 );
   nor U37795 ( n36492,n36493,n36494 );
   nor U37796 ( n36494,n36337,n33678 );
   not U37797 ( n33678,p3_instqueue_reg_14__4_ );
   nor U37798 ( n36493,n36338,n33675 );
   not U37799 ( n33675,p3_instqueue_reg_13__4_ );
   nor U37800 ( n36491,n36495,n36496 );
   nor U37801 ( n36496,n36341,n33669 );
   not U37802 ( n33669,p3_instqueue_reg_12__4_ );
   nor U37803 ( n36495,n36342,n33686 );
   not U37804 ( n33686,p3_instqueue_reg_6__4_ );
   nand U37805 ( n36489,n36497,n36498 );
   nor U37806 ( n36498,n36499,n36500 );
   nor U37807 ( n36500,n36347,n33701 );
   not U37808 ( n33701,p3_instqueue_reg_5__4_ );
   nor U37809 ( n36499,n36348,n33665 );
   not U37810 ( n33665,p3_instqueue_reg_4__4_ );
   nor U37811 ( n36497,n36501,n36502 );
   nor U37812 ( n36502,n36351,n33697 );
   not U37813 ( n33697,p3_instqueue_reg_2__4_ );
   nor U37814 ( n36501,n36352,n33696 );
   not U37815 ( n33696,p3_instqueue_reg_1__4_ );
   nor U37816 ( n36487,n36503,n36504 );
   nand U37817 ( n36504,n36505,n36506 );
   nor U37818 ( n36506,n36507,n36508 );
   nor U37819 ( n36508,n36359,n30683 );
   not U37820 ( n30683,p3_instqueue_reg_0__4_ );
   nor U37821 ( n36507,n36360,n33691 );
   not U37822 ( n33691,p3_instqueue_reg_10__4_ );
   nor U37823 ( n36505,n36509,n36510 );
   nor U37824 ( n36510,n36363,n33666 );
   not U37825 ( n33666,p3_instqueue_reg_8__4_ );
   nor U37826 ( n36509,n33877,n33687 );
   not U37827 ( n33687,p3_instqueue_reg_7__4_ );
   nand U37828 ( n36503,n36511,n36512 );
   nor U37829 ( n36512,n36513,n36514 );
   nor U37830 ( n36514,n36368,n33700 );
   not U37831 ( n33700,p3_instqueue_reg_3__4_ );
   nor U37832 ( n36513,n35468,n33679 );
   not U37833 ( n33679,p3_instqueue_reg_15__4_ );
   nor U37834 ( n36511,n36515,n36516 );
   nor U37835 ( n36516,n36371,n33674 );
   not U37836 ( n33674,p3_instqueue_reg_11__4_ );
   nor U37837 ( n36515,n36372,n33690 );
   not U37838 ( n33690,p3_instqueue_reg_9__4_ );
   nand U37839 ( n30691,n36517,n36518 );
   nor U37840 ( n36518,n36519,n36520 );
   nand U37841 ( n36520,n36521,n36522 );
   nor U37842 ( n36522,n36523,n36524 );
   nor U37843 ( n36524,n36337,n33634 );
   not U37844 ( n33634,p3_instqueue_reg_14__3_ );
   nor U37845 ( n36523,n36338,n33631 );
   not U37846 ( n33631,p3_instqueue_reg_13__3_ );
   nor U37847 ( n36521,n36525,n36526 );
   nor U37848 ( n36526,n36341,n33644 );
   not U37849 ( n33644,p3_instqueue_reg_12__3_ );
   nor U37850 ( n36525,n36342,n33618 );
   not U37851 ( n33618,p3_instqueue_reg_6__3_ );
   nand U37852 ( n36519,n36527,n36528 );
   nor U37853 ( n36528,n36529,n36530 );
   nor U37854 ( n36530,n36347,n33613 );
   not U37855 ( n33613,p3_instqueue_reg_5__3_ );
   nor U37856 ( n36529,n36348,n33640 );
   not U37857 ( n33640,p3_instqueue_reg_4__3_ );
   nor U37858 ( n36527,n36531,n36532 );
   nor U37859 ( n36532,n36351,n33609 );
   not U37860 ( n33609,p3_instqueue_reg_2__3_ );
   nor U37861 ( n36531,n36352,n33608 );
   not U37862 ( n33608,p3_instqueue_reg_1__3_ );
   nor U37863 ( n36517,n36533,n36534 );
   nand U37864 ( n36534,n36535,n36536 );
   nor U37865 ( n36536,n36537,n36538 );
   nor U37866 ( n36538,n36359,n30694 );
   not U37867 ( n30694,p3_instqueue_reg_0__3_ );
   nor U37868 ( n36537,n36360,n33623 );
   not U37869 ( n33623,p3_instqueue_reg_10__3_ );
   nor U37870 ( n36535,n36539,n36540 );
   nor U37871 ( n36540,n36363,n33641 );
   not U37872 ( n33641,p3_instqueue_reg_8__3_ );
   nor U37873 ( n36539,n33877,n33619 );
   not U37874 ( n33619,p3_instqueue_reg_7__3_ );
   nand U37875 ( n36533,n36541,n36542 );
   nor U37876 ( n36542,n36543,n36544 );
   nor U37877 ( n36544,n36368,n33612 );
   not U37878 ( n33612,p3_instqueue_reg_3__3_ );
   nor U37879 ( n36543,n35468,n33635 );
   not U37880 ( n33635,p3_instqueue_reg_15__3_ );
   nor U37881 ( n36541,n36545,n36546 );
   nor U37882 ( n36546,n36371,n33630 );
   not U37883 ( n33630,p3_instqueue_reg_11__3_ );
   nor U37884 ( n36545,n36372,n33622 );
   not U37885 ( n33622,p3_instqueue_reg_9__3_ );
   nor U37886 ( n35470,n29315,n31847 );
   nor U37887 ( n31847,n29350,n29304 );
   not U37888 ( n29304,n29366 );
   nor U37889 ( n29315,n29366,n29350 );
   nand U37890 ( n29350,n36547,n36548 );
   nor U37891 ( n36548,n36549,n36550 );
   nand U37892 ( n36550,n36551,n36552 );
   nor U37893 ( n36552,n36553,n36554 );
   nor U37894 ( n36554,n36337,n33463 );
   not U37895 ( n33463,p3_instqueue_reg_14__0_ );
   nor U37896 ( n36553,n36338,n33459 );
   not U37897 ( n33459,p3_instqueue_reg_13__0_ );
   nor U37898 ( n36551,n36555,n36556 );
   nor U37899 ( n36556,n36341,n33477 );
   not U37900 ( n33477,p3_instqueue_reg_12__0_ );
   nor U37901 ( n36555,n36342,n33441 );
   not U37902 ( n33441,p3_instqueue_reg_6__0_ );
   nand U37903 ( n36549,n36557,n36558 );
   nor U37904 ( n36558,n36559,n36560 );
   nor U37905 ( n36560,n36347,n33435 );
   not U37906 ( n33435,p3_instqueue_reg_5__0_ );
   nor U37907 ( n36559,n36348,n33471 );
   not U37908 ( n33471,p3_instqueue_reg_4__0_ );
   nor U37909 ( n36557,n36561,n36562 );
   nor U37910 ( n36562,n36351,n33429 );
   not U37911 ( n33429,p3_instqueue_reg_2__0_ );
   nor U37912 ( n36561,n36352,n33427 );
   not U37913 ( n33427,p3_instqueue_reg_1__0_ );
   nor U37914 ( n36547,n36563,n36564 );
   nand U37915 ( n36564,n36565,n36566 );
   nor U37916 ( n36566,n36567,n36568 );
   nor U37917 ( n36568,n36359,n33479 );
   not U37918 ( n33479,p3_instqueue_reg_0__0_ );
   nor U37919 ( n36567,n36360,n33449 );
   not U37920 ( n33449,p3_instqueue_reg_10__0_ );
   nor U37921 ( n36565,n36569,n36570 );
   nor U37922 ( n36570,n36363,n33473 );
   not U37923 ( n33473,p3_instqueue_reg_8__0_ );
   nor U37924 ( n36569,n33877,n33443 );
   not U37925 ( n33443,p3_instqueue_reg_7__0_ );
   nand U37926 ( n36563,n36571,n36572 );
   nor U37927 ( n36572,n36573,n36574 );
   nor U37928 ( n36574,n36368,n33433 );
   not U37929 ( n33433,p3_instqueue_reg_3__0_ );
   nor U37930 ( n36573,n35468,n33465 );
   not U37931 ( n33465,p3_instqueue_reg_15__0_ );
   nor U37932 ( n36571,n36575,n36576 );
   nor U37933 ( n36576,n36371,n33457 );
   not U37934 ( n33457,p3_instqueue_reg_11__0_ );
   nor U37935 ( n36575,n36372,n33447 );
   not U37936 ( n33447,p3_instqueue_reg_9__0_ );
   nand U37937 ( n29366,n36577,n36578 );
   nor U37938 ( n36578,n36579,n36580 );
   nand U37939 ( n36580,n36581,n36582 );
   nor U37940 ( n36582,n36583,n36584 );
   nor U37941 ( n36584,n36337,n33524 );
   not U37942 ( n33524,p3_instqueue_reg_14__1_ );
   nand U37943 ( n36337,n28883,n34597 );
   nor U37944 ( n36583,n36338,n33521 );
   not U37945 ( n33521,p3_instqueue_reg_13__1_ );
   nand U37946 ( n36338,n28883,n34619 );
   nor U37947 ( n36581,n36585,n36586 );
   nor U37948 ( n36586,n36341,n33534 );
   not U37949 ( n33534,p3_instqueue_reg_12__1_ );
   nand U37950 ( n36341,n28883,n34594 );
   nor U37951 ( n28883,n29254,n29257 );
   nor U37952 ( n36585,n36342,n33508 );
   not U37953 ( n33508,p3_instqueue_reg_6__1_ );
   nand U37954 ( n36342,n34597,n34627 );
   nand U37955 ( n36579,n36587,n36588 );
   nor U37956 ( n36588,n36589,n36590 );
   nor U37957 ( n36590,n36347,n33503 );
   not U37958 ( n33503,p3_instqueue_reg_5__1_ );
   nand U37959 ( n36347,n34619,n34627 );
   nor U37960 ( n36589,n36348,n33530 );
   not U37961 ( n33530,p3_instqueue_reg_4__1_ );
   nand U37962 ( n36348,n34594,n34627 );
   nor U37963 ( n36587,n36591,n36592 );
   nor U37964 ( n36592,n36351,n33499 );
   not U37965 ( n33499,p3_instqueue_reg_2__1_ );
   nand U37966 ( n36351,n35302,n29254 );
   nor U37967 ( n36591,n36352,n33498 );
   not U37968 ( n33498,p3_instqueue_reg_1__1_ );
   nand U37969 ( n36352,n35301,n29254 );
   nor U37970 ( n36577,n36593,n36594 );
   nand U37971 ( n36594,n36595,n36596 );
   nor U37972 ( n36596,n36597,n36598 );
   nor U37973 ( n36598,n36359,n30716 );
   not U37974 ( n30716,p3_instqueue_reg_0__1_ );
   nand U37975 ( n36359,n35181,n29254 );
   nor U37976 ( n36597,n36360,n33513 );
   not U37977 ( n33513,p3_instqueue_reg_10__1_ );
   nand U37978 ( n36360,n35302,p3_instqueuerd_addr_reg_3_ );
   nor U37979 ( n35302,n29356,p3_instqueuerd_addr_reg_2_ );
   not U37980 ( n29356,n34597 );
   nor U37981 ( n34597,n29341,p3_instqueuerd_addr_reg_0_ );
   nor U37982 ( n36595,n36599,n36600 );
   nor U37983 ( n36600,n36363,n33531 );
   not U37984 ( n33531,p3_instqueue_reg_8__1_ );
   nand U37985 ( n36363,n35181,p3_instqueuerd_addr_reg_3_ );
   nor U37986 ( n35181,n30802,p3_instqueuerd_addr_reg_2_ );
   not U37987 ( n30802,n34594 );
   nor U37988 ( n34594,p3_instqueuerd_addr_reg_0_,p3_instqueuerd_addr_reg_1_ );
   nor U37989 ( n36599,n33877,n33509 );
   not U37990 ( n33509,p3_instqueue_reg_7__1_ );
   nand U37991 ( n33877,n29294,n34627 );
   nor U37992 ( n34627,n29257,p3_instqueuerd_addr_reg_3_ );
   nand U37993 ( n36593,n36601,n36602 );
   nor U37994 ( n36602,n36603,n36604 );
   nor U37995 ( n36604,n36368,n33502 );
   not U37996 ( n33502,p3_instqueue_reg_3__1_ );
   nand U37997 ( n36368,n35284,n29254 );
   nor U37998 ( n36603,n35468,n33525 );
   not U37999 ( n33525,p3_instqueue_reg_15__1_ );
   not U38000 ( n35468,n35433 );
   nor U38001 ( n35433,n29274,n29254 );
   not U38002 ( n29254,p3_instqueuerd_addr_reg_3_ );
   not U38003 ( n29274,n35282 );
   nor U38004 ( n35282,n29256,n29257 );
   nor U38005 ( n36601,n36605,n36606 );
   nor U38006 ( n36606,n36371,n33520 );
   not U38007 ( n33520,p3_instqueue_reg_11__1_ );
   nand U38008 ( n36371,n35284,p3_instqueuerd_addr_reg_3_ );
   nor U38009 ( n35284,n29256,p3_instqueuerd_addr_reg_2_ );
   not U38010 ( n29256,n29294 );
   nor U38011 ( n29294,n29341,n29275 );
   not U38012 ( n29341,p3_instqueuerd_addr_reg_1_ );
   nor U38013 ( n36605,n36372,n33512 );
   not U38014 ( n33512,p3_instqueue_reg_9__1_ );
   nand U38015 ( n36372,n35301,p3_instqueuerd_addr_reg_3_ );
   and U38016 ( n35301,n34619,n29257 );
   not U38017 ( n29257,p3_instqueuerd_addr_reg_2_ );
   nor U38018 ( n34619,n29275,p3_instqueuerd_addr_reg_1_ );
   not U38019 ( n29275,p3_instqueuerd_addr_reg_0_ );
   nand U38020 ( n36320,n28775,p3_state2_reg_0_ );
   and U38021 ( n28775,n28795,n28856 );
   not U38022 ( n28856,p3_state2_reg_1_ );
   nor U38023 ( n28795,p3_state2_reg_2_,p3_state2_reg_3_ );
   nand U38024 ( n36607,p3_ads_n_reg,p3_state_reg_0_ );
   nor U38025 ( n28895,n36608,n29101 );
   nor U38026 ( n29101,p3_state_reg_0_,p3_state_reg_1_ );
   and U38027 ( n36608,n36609,p3_state_reg_0_ );
   nor U38028 ( n36609,p3_state_reg_2_,n29074 );
   not U38029 ( n29074,p3_state_reg_1_ );
   nand U38030 ( n36611,p2_readrequest_reg,n36612 );
   nand U38031 ( n36610,n36613,n36614 );
   nand U38032 ( n36614,n36615,p2_state2_reg_2_ );
   nand U38033 ( n36613,n36612,n36616 );
   nand U38034 ( n36618,p2_m_io_n_reg,n28377 );
   nand U38035 ( n36617,p2_memoryfetch_reg,n36620 );
   nand U38036 ( n36622,n36623,p2_requestpending_reg );
   not U38037 ( n36623,n36624 );
   nand U38038 ( n36621,n36625,n36624 );
   nand U38039 ( n36624,n36626,n36627 );
   nor U38040 ( n36627,n36628,n36629 );
   nor U38041 ( n36626,n36630,n36631 );
   nor U38042 ( n36631,p2_state2_reg_0_,n36632 );
   nor U38043 ( n36630,n28178,n36633 );
   nand U38044 ( n36633,n36634,n36635 );
   nand U38045 ( n36625,n36636,n36637 );
   nor U38046 ( n36637,n36638,n36639 );
   nand U38047 ( n36639,n36640,n36641 );
   not U38048 ( n36641,n36642 );
   nand U38049 ( n36640,n36643,n36644 );
   nor U38050 ( n36643,n36645,n36646 );
   nor U38051 ( n36645,n36647,n36648 );
   nor U38052 ( n36638,n36649,n36635 );
   nor U38053 ( n36649,n36650,n36651 );
   nor U38054 ( n36636,n36652,n36653 );
   nor U38055 ( n36652,n36654,n36655 );
   nand U38056 ( n36657,n36658,n36659 );
   nand U38057 ( n36656,p2_more_reg,n36660 );
   or U38058 ( n36662,n36619,p2_readrequest_reg );
   nand U38059 ( n36661,p2_w_r_n_reg,n28377 );
   nand U38060 ( n36664,n36665,p2_instqueuewr_addr_reg_0_ );
   nand U38061 ( n36663,n36666,n36667 );
   nand U38062 ( n36666,n36668,n36669 );
   nand U38063 ( n36669,n36670,p2_state2_reg_3_ );
   nor U38064 ( n36668,n36671,n36672 );
   nor U38065 ( n36672,n36673,n36674 );
   nand U38066 ( n36676,n36665,p2_instqueuewr_addr_reg_1_ );
   nand U38067 ( n36675,n36677,n36667 );
   nand U38068 ( n36677,n36678,n36679 );
   nand U38069 ( n36679,p2_state2_reg_3_,n36680 );
   nor U38070 ( n36678,n36681,n36682 );
   nor U38071 ( n36682,n36683,n36684 );
   nor U38072 ( n36681,n36685,n36686 );
   nor U38073 ( n36685,n36687,n36688 );
   nand U38074 ( n36690,n36665,p2_instqueuewr_addr_reg_2_ );
   nand U38075 ( n36689,n36691,n36667 );
   nand U38076 ( n36691,n36692,n36693 );
   nand U38077 ( n36693,n36694,p2_state2_reg_3_ );
   nor U38078 ( n36692,n36695,n36696 );
   nor U38079 ( n36696,n36683,n36697 );
   nor U38080 ( n36695,n36686,n36698 );
   nand U38081 ( n36698,n36699,n36700 );
   or U38082 ( n36699,n36701,n36702 );
   nand U38083 ( n36704,n36665,p2_instqueuewr_addr_reg_3_ );
   nand U38084 ( n36703,n36705,n36667 );
   nand U38085 ( n36705,n36706,n36707 );
   nand U38086 ( n36707,p2_state2_reg_3_,n36708 );
   nor U38087 ( n36706,n36709,n36710 );
   nor U38088 ( n36710,n36683,n36711 );
   nor U38089 ( n36683,n36712,n36713 );
   nor U38090 ( n36709,n36714,n36686 );
   nor U38091 ( n36714,n36715,n36716 );
   nor U38092 ( n36715,n36717,n36718 );
   nand U38093 ( n36720,p2_instqueuerd_addr_reg_0_,n36721 );
   nand U38094 ( n36721,n36722,n36723 );
   nand U38095 ( n36723,n36713,n36724 );
   nand U38096 ( n36719,n36725,n36722 );
   nand U38097 ( n36725,n36726,n36727 );
   nand U38098 ( n36727,n36728,n36729 );
   nor U38099 ( n36726,n36730,n36731 );
   nor U38100 ( n36731,n36732,n36632 );
   nor U38101 ( n36730,n36733,n28181 );
   nand U38102 ( n36735,n36736,p2_instqueuerd_addr_reg_1_ );
   nand U38103 ( n36734,n36737,n36722 );
   nand U38104 ( n36737,n36738,n36739 );
   nand U38105 ( n36739,n36728,n36740 );
   nor U38106 ( n36738,n36741,n36742 );
   nor U38107 ( n36742,n36743,n36632 );
   nor U38108 ( n36741,n36744,n36745 );
   not U38109 ( n36744,n36746 );
   nand U38110 ( n36748,n36736,p2_instqueuerd_addr_reg_2_ );
   nand U38111 ( n36747,n36749,n36722 );
   nand U38112 ( n36749,n36750,n36751 );
   nand U38113 ( n36751,n36728,n36752 );
   nor U38114 ( n36750,n36753,n36754 );
   nor U38115 ( n36754,n36745,n36746 );
   nand U38116 ( n36746,n36755,n36756 );
   nand U38117 ( n36756,n36757,n36758 );
   or U38118 ( n36755,n36759,n36757 );
   nand U38119 ( n36745,n36733,p2_state2_reg_1_ );
   and U38120 ( n36733,n36760,n36761 );
   nand U38121 ( n36761,n36757,n36762 );
   nand U38122 ( n36760,n36763,n36764 );
   nor U38123 ( n36753,n36765,n36632 );
   nand U38124 ( n36767,n36736,p2_instqueuerd_addr_reg_3_ );
   nand U38125 ( n36766,n36768,n36722 );
   nand U38126 ( n36768,n36769,n36770 );
   nand U38127 ( n36770,n36713,n36771 );
   nand U38128 ( n36769,n36728,n36772 );
   nand U38129 ( n36774,n36775,n36776 );
   nor U38130 ( n36775,n36777,n36632 );
   nor U38131 ( n36777,n36778,p2_instqueuerd_addr_reg_4_ );
   nor U38132 ( n36778,n36779,n36780 );
   nand U38133 ( n36780,p2_instqueuerd_addr_reg_3_,n36722 );
   nand U38134 ( n36773,n36736,p2_instqueuerd_addr_reg_4_ );
   not U38135 ( n36736,n36722 );
   nand U38136 ( n36722,n36781,n36782 );
   nand U38137 ( n36782,p2_state2_reg_3_,n27895 );
   nor U38138 ( n36781,n36784,n36785 );
   nor U38139 ( n36785,n36786,n36787 );
   nand U38140 ( n36789,p2_state2_reg_3_,n36790 );
   nand U38141 ( n36790,p2_state2_reg_0_,n36791 );
   nand U38142 ( n36793,p2_datawidth_reg_1_,n28163 );
   nand U38143 ( n36792,n36794,n28166 );
   nand U38144 ( n36794,n28898,n36795 );
   nand U38145 ( n36797,n36798,n28165 );
   nor U38146 ( n36798,bs16,n36799 );
   nand U38147 ( n36796,p2_datawidth_reg_0_,n28163 );
   nand U38148 ( n36801,p2_be_n_reg_0_,n36619 );
   nand U38149 ( n36800,p2_byteenable_reg_0_,n36620 );
   nand U38150 ( n36803,p2_be_n_reg_1_,n36619 );
   nand U38151 ( n36802,p2_byteenable_reg_1_,n36620 );
   nand U38152 ( n36805,p2_be_n_reg_2_,n28377 );
   nand U38153 ( n36804,p2_byteenable_reg_2_,n36620 );
   nand U38154 ( n36807,p2_be_n_reg_3_,n28377 );
   nand U38155 ( n36806,p2_byteenable_reg_3_,n36620 );
   nand U38156 ( n36809,p2_address_reg_29_,n28377 );
   nor U38157 ( n36808,n36810,n36811 );
   nor U38158 ( n36811,n28388,n36813 );
   nor U38159 ( n36810,n28385,n36815 );
   nand U38160 ( n36817,p2_address_reg_28_,n28377 );
   nor U38161 ( n36816,n36818,n36819 );
   nor U38162 ( n36819,n36815,n28388 );
   nor U38163 ( n36818,n28386,n36820 );
   nand U38164 ( n36822,p2_address_reg_27_,n36619 );
   nor U38165 ( n36821,n36823,n36824 );
   nor U38166 ( n36824,n28387,n36820 );
   nor U38167 ( n36823,n28386,n36825 );
   nand U38168 ( n36827,p2_address_reg_26_,n28377 );
   nor U38169 ( n36826,n36828,n36829 );
   nor U38170 ( n36829,n36812,n36825 );
   nor U38171 ( n36828,n36814,n36830 );
   nand U38172 ( n36832,p2_address_reg_25_,n28377 );
   nor U38173 ( n36831,n36833,n36834 );
   nor U38174 ( n36834,n36812,n36830 );
   nor U38175 ( n36833,n36814,n36835 );
   nand U38176 ( n36837,p2_address_reg_24_,n28377 );
   nor U38177 ( n36836,n36838,n36839 );
   nor U38178 ( n36839,n28387,n36835 );
   nor U38179 ( n36838,n28385,n36840 );
   nand U38180 ( n36842,p2_address_reg_23_,n28377 );
   nor U38181 ( n36841,n36843,n36844 );
   nor U38182 ( n36844,n36812,n36840 );
   nor U38183 ( n36843,n28385,n36845 );
   nand U38184 ( n36847,p2_address_reg_22_,n28377 );
   nor U38185 ( n36846,n36848,n36849 );
   nor U38186 ( n36849,n28388,n36845 );
   nor U38187 ( n36848,n36814,n36850 );
   nand U38188 ( n36852,p2_address_reg_21_,n28377 );
   nor U38189 ( n36851,n36853,n36854 );
   nor U38190 ( n36854,n28387,n36850 );
   nor U38191 ( n36853,n28386,n36855 );
   nand U38192 ( n36857,p2_address_reg_20_,n36619 );
   nor U38193 ( n36856,n36858,n36859 );
   nor U38194 ( n36859,n36812,n36855 );
   nor U38195 ( n36858,n28385,n36860 );
   nand U38196 ( n36862,p2_address_reg_19_,n28377 );
   nor U38197 ( n36861,n36863,n36864 );
   nor U38198 ( n36864,n28388,n36860 );
   nor U38199 ( n36863,n36814,n36865 );
   nand U38200 ( n36867,p2_address_reg_18_,n36619 );
   nor U38201 ( n36866,n36868,n36869 );
   nor U38202 ( n36869,n28387,n36865 );
   nor U38203 ( n36868,n28386,n36870 );
   nand U38204 ( n36872,p2_address_reg_17_,n28377 );
   nor U38205 ( n36871,n36873,n36874 );
   nor U38206 ( n36874,n28387,n36870 );
   nor U38207 ( n36873,n28385,n36875 );
   nand U38208 ( n36877,p2_address_reg_16_,n28377 );
   nor U38209 ( n36876,n36878,n36879 );
   nor U38210 ( n36879,n28387,n36875 );
   nor U38211 ( n36878,n28386,n36880 );
   nand U38212 ( n36882,p2_address_reg_15_,n28377 );
   nor U38213 ( n36881,n36883,n36884 );
   nor U38214 ( n36884,n36812,n36880 );
   nor U38215 ( n36883,n36814,n36885 );
   nand U38216 ( n36887,p2_address_reg_14_,n28377 );
   nor U38217 ( n36886,n36888,n36889 );
   nor U38218 ( n36889,n28388,n36885 );
   nor U38219 ( n36888,n28385,n36890 );
   nand U38220 ( n36892,p2_address_reg_13_,n28377 );
   nor U38221 ( n36891,n36893,n36894 );
   nor U38222 ( n36894,n36812,n36890 );
   nor U38223 ( n36893,n36814,n36895 );
   nand U38224 ( n36897,p2_address_reg_12_,n36619 );
   nor U38225 ( n36896,n36898,n36899 );
   nor U38226 ( n36899,n28388,n36895 );
   nor U38227 ( n36898,n28386,n36900 );
   nand U38228 ( n36902,p2_address_reg_11_,n28377 );
   nor U38229 ( n36901,n36903,n36904 );
   nor U38230 ( n36904,n36812,n36900 );
   nor U38231 ( n36903,n36814,n36905 );
   nand U38232 ( n36907,p2_address_reg_10_,n28377 );
   nor U38233 ( n36906,n36908,n36909 );
   nor U38234 ( n36909,n28387,n36905 );
   nor U38235 ( n36908,n28385,n36910 );
   nand U38236 ( n36912,p2_address_reg_9_,n36619 );
   nor U38237 ( n36911,n36913,n36914 );
   nor U38238 ( n36914,n28388,n36910 );
   nor U38239 ( n36913,n28386,n36915 );
   nand U38240 ( n36917,p2_address_reg_8_,n36619 );
   nor U38241 ( n36916,n36918,n36919 );
   nor U38242 ( n36919,n28388,n36915 );
   nor U38243 ( n36918,n28385,n36920 );
   nand U38244 ( n36922,p2_address_reg_7_,n28377 );
   nor U38245 ( n36921,n36923,n36924 );
   nor U38246 ( n36924,n28387,n36920 );
   nor U38247 ( n36923,n36814,n36925 );
   nand U38248 ( n36927,p2_address_reg_6_,n36619 );
   nor U38249 ( n36926,n36928,n36929 );
   nor U38250 ( n36929,n36812,n36925 );
   nor U38251 ( n36928,n28386,n36930 );
   nand U38252 ( n36932,p2_address_reg_5_,n28377 );
   nor U38253 ( n36931,n36933,n36934 );
   nor U38254 ( n36934,n28388,n36930 );
   nor U38255 ( n36933,n28385,n36935 );
   nand U38256 ( n36937,p2_address_reg_4_,n36619 );
   nor U38257 ( n36936,n36938,n36939 );
   nor U38258 ( n36939,n28387,n36935 );
   nor U38259 ( n36938,n36814,n36940 );
   nand U38260 ( n36942,p2_address_reg_3_,n36619 );
   nor U38261 ( n36941,n36943,n36944 );
   nor U38262 ( n36944,n36812,n36940 );
   nor U38263 ( n36943,n28386,n36945 );
   nand U38264 ( n36947,p2_address_reg_2_,n36619 );
   nor U38265 ( n36946,n36948,n36949 );
   nor U38266 ( n36949,n28388,n36945 );
   nor U38267 ( n36948,n36950,n28386 );
   nand U38268 ( n36952,p2_address_reg_1_,n28377 );
   nor U38269 ( n36951,n36953,n36954 );
   nor U38270 ( n36954,n36950,n28387 );
   nor U38271 ( n36953,n36955,n28385 );
   nand U38272 ( n36957,p2_address_reg_0_,n36619 );
   nor U38273 ( n36956,n36958,n36959 );
   nor U38274 ( n36959,n36955,n36812 );
   not U38275 ( n36812,n36960 );
   nor U38276 ( n36958,n36961,n36814 );
   not U38277 ( n36814,n36962 );
   nand U38278 ( n36964,n36965,n36966 );
   nor U38279 ( n36966,n36967,n36968 );
   nor U38280 ( n36968,p2_requestpending_reg,hold );
   nor U38281 ( n36967,n36969,n36970 );
   nor U38282 ( n36970,p2_requestpending_reg,n36795 );
   nor U38283 ( n36965,n36971,n36972 );
   nor U38284 ( n36971,n29075,n36973 );
   nor U38285 ( n36963,n36962,n36974 );
   nor U38286 ( n36974,n36975,n36976 );
   nor U38287 ( n36975,n36969,n36977 );
   nand U38288 ( n36977,n36978,n36979 );
   nand U38289 ( n36979,n29075,n36972 );
   nand U38290 ( n36978,p2_state_reg_0_,hold );
   nor U38291 ( n36962,n36976,n36619 );
   nor U38292 ( n36981,n36960,n36969 );
   nor U38293 ( n36960,n36619,p2_state_reg_2_ );
   nor U38294 ( n36980,n36982,n36983 );
   nand U38295 ( n36983,n36984,n36985 );
   nand U38296 ( n36985,n36986,n36976 );
   nor U38297 ( n36986,n29093,n36973 );
   or U38298 ( n36984,n36987,n36976 );
   nor U38299 ( n36982,n36972,n36988 );
   nand U38300 ( n36988,p2_requestpending_reg,n36989 );
   nand U38301 ( n36989,hold,n36795 );
   nor U38302 ( n36991,n36992,n36993 );
   nor U38303 ( n36993,p2_state_reg_2_,n36994 );
   nor U38304 ( n36994,n36969,n36972 );
   nor U38305 ( n36969,n36635,n36973 );
   nor U38306 ( n36992,n29093,n36995 );
   nand U38307 ( n36995,n36996,n36997 );
   nand U38308 ( n36997,n36973,n36976 );
   not U38309 ( n36976,p2_state_reg_2_ );
   nand U38310 ( n36996,p2_state_reg_1_,n36972 );
   nor U38311 ( n36990,n36998,n36999 );
   nor U38312 ( n36999,p2_requestpending_reg,n36620 );
   nor U38313 ( n36998,n29075,n36987 );
   nand U38314 ( n37031,p2_state2_reg_1_,n37032 );
   nand U38315 ( n37032,n37033,n37034 );
   nand U38316 ( n37034,n36642,n36635 );
   nand U38317 ( n37033,p2_statebs16_reg,n27895 );
   nor U38318 ( n37030,n37035,n36634 );
   nand U38319 ( n37037,p2_state2_reg_1_,n37038 );
   nand U38320 ( n37038,n36791,n37039 );
   nor U38321 ( n37036,n37040,n37041 );
   nor U38322 ( n37041,n37042,n37043 );
   nor U38323 ( n37043,n37044,n37045 );
   nor U38324 ( n37044,n36632,n37046 );
   nand U38325 ( n37046,p2_state2_reg_0_,n36635 );
   not U38326 ( n36632,n36713 );
   nor U38327 ( n37048,n37049,n37050 );
   nand U38328 ( n37050,n37039,n37051 );
   nand U38329 ( n37039,n36642,n37052 );
   nor U38330 ( n37049,n37042,n37053 );
   nor U38331 ( n37053,n37054,n36634 );
   nor U38332 ( n37054,p2_state2_reg_0_,n37055 );
   and U38333 ( n37055,n28178,n36728 );
   nor U38334 ( n37047,n37056,n37057 );
   and U38335 ( n37057,n37058,n37045 );
   nor U38336 ( n37056,n37059,n36783 );
   nor U38337 ( n37059,n36671,n37042 );
   not U38338 ( n37042,n36791 );
   nand U38339 ( n36791,n37060,n37061 );
   nor U38340 ( n37061,n37062,n37063 );
   nor U38341 ( n37063,n37064,n36783 );
   nor U38342 ( n37064,n37058,n37065 );
   nand U38343 ( n37065,n37066,n28179 );
   nand U38344 ( n37066,n37067,n37068 );
   nand U38345 ( n37058,n37069,n37070 );
   nor U38346 ( n37070,n37071,n37072 );
   nand U38347 ( n37072,n37073,n37074 );
   nand U38348 ( n37074,n37075,n37076 );
   or U38349 ( n37076,p2_more_reg,p2_flush_reg );
   nand U38350 ( n37073,p2_instqueuerd_addr_reg_4_,n37077 );
   nand U38351 ( n37077,n37078,n37079 );
   nand U38352 ( n37071,n37080,n37081 );
   nand U38353 ( n37081,n37082,n37083 );
   nand U38354 ( n37083,p2_instqueuewr_addr_reg_3_,n37084 );
   nor U38355 ( n37082,p2_instqueuewr_addr_reg_4_,n37085 );
   nor U38356 ( n37085,n37086,n37087 );
   nand U38357 ( n37087,n37088,n37089 );
   nand U38358 ( n37089,n37090,n37091 );
   nand U38359 ( n37091,p2_instqueuewr_addr_reg_2_,n37092 );
   nor U38360 ( n37090,n37093,n37094 );
   nor U38361 ( n37094,n37095,n37096 );
   nor U38362 ( n37095,n37097,n37098 );
   nand U38363 ( n37098,n37099,n37100 );
   nand U38364 ( n37100,n36743,n37079 );
   nand U38365 ( n37099,n36786,n37101 );
   nand U38366 ( n37101,p2_instqueuerd_addr_reg_1_,n37102 );
   nor U38367 ( n37097,n37103,n37102 );
   nor U38368 ( n37093,n37102,n37104 );
   nand U38369 ( n37104,n37105,n37106 );
   nand U38370 ( n37106,n36786,p2_instqueuerd_addr_reg_1_ );
   nand U38371 ( n37105,n37107,n37079 );
   nand U38372 ( n37107,n36743,n37108 );
   not U38373 ( n37108,n37103 );
   nand U38374 ( n37103,n36732,n37109 );
   nand U38375 ( n37109,p2_instqueuerd_addr_reg_0_,n36724 );
   and U38376 ( n36732,n37110,n37111 );
   nand U38377 ( n37111,n37112,n37113 );
   and U38378 ( n37112,n37114,n37115 );
   nand U38379 ( n37110,n37116,n37117 );
   and U38380 ( n36743,n37118,n37119 );
   nand U38381 ( n37119,n36724,n37120 );
   not U38382 ( n36724,n37121 );
   nor U38383 ( n37118,n37122,n37123 );
   nor U38384 ( n37123,n37124,n37125 );
   nor U38385 ( n37122,n37126,n37127 );
   nand U38386 ( n37127,n37113,n37115 );
   nand U38387 ( n37115,n37128,n37129 );
   nand U38388 ( n37129,n37130,n37131 );
   nand U38389 ( n37131,n37132,n37133 );
   nand U38390 ( n37128,n37134,n37135 );
   nand U38391 ( n37135,n37132,n37136 );
   nand U38392 ( n37102,p2_instqueuewr_addr_reg_0_,n37137 );
   nand U38393 ( n37137,n36786,p2_instqueuerd_addr_reg_0_ );
   or U38394 ( n37088,n37084,p2_instqueuewr_addr_reg_3_ );
   nor U38395 ( n37086,p2_instqueuewr_addr_reg_2_,n37092 );
   nand U38396 ( n37080,n37138,n36776 );
   nor U38397 ( n37138,n37139,n36779 );
   nor U38398 ( n37069,n36659,n37140 );
   nand U38399 ( n37140,n37141,n37142 );
   or U38400 ( n37142,n37092,n37084 );
   nand U38401 ( n37084,n37143,n37144 );
   nand U38402 ( n37144,n36786,n37139 );
   or U38403 ( n37143,n36771,n36786 );
   nand U38404 ( n36771,n37145,n37146 );
   nor U38405 ( n37146,n37147,n37148 );
   nor U38406 ( n37148,n37149,n37150 );
   nor U38407 ( n37147,n37151,n37152 );
   xor U38408 ( n37152,n37153,n37139 );
   nand U38409 ( n37153,n37154,n37155 );
   nor U38410 ( n37145,n37156,n37157 );
   nor U38411 ( n37157,n37121,n37158 );
   nor U38412 ( n37156,n37124,n37159 );
   nand U38413 ( n37092,n37160,n37161 );
   nand U38414 ( n37161,n36786,n37154 );
   not U38415 ( n36786,n37079 );
   nand U38416 ( n37160,n36765,n37079 );
   nand U38417 ( n37079,n37162,n37163 );
   nor U38418 ( n37163,n37164,n37165 );
   nor U38419 ( n37165,n37166,n37167 );
   nor U38420 ( n37164,n37168,n37169 );
   nand U38421 ( n37169,n37170,n37171 );
   nor U38422 ( n37162,n37172,n37173 );
   and U38423 ( n36765,n37174,n37175 );
   nor U38424 ( n37175,n37176,n37177 );
   nor U38425 ( n37177,n37151,n37178 );
   nor U38426 ( n37151,n37179,n37180 );
   nor U38427 ( n37176,n37181,n37149 );
   nor U38428 ( n37149,n37182,n37183 );
   nor U38429 ( n37174,n37184,n37185 );
   nor U38430 ( n37185,n37121,n37186 );
   nor U38431 ( n37121,n37187,n37188 );
   nor U38432 ( n37184,n37124,n37189 );
   not U38433 ( n37124,n37117 );
   nand U38434 ( n37117,n37190,n37191 );
   nor U38435 ( n37191,n37192,n37193 );
   nor U38436 ( n37193,n37194,n37195 );
   not U38437 ( n37141,n37196 );
   nand U38438 ( n36659,n37197,n37198 );
   nor U38439 ( n37198,n37199,n37200 );
   and U38440 ( n37200,n37201,n37202 );
   nor U38441 ( n37199,n37203,n37204 );
   nand U38442 ( n37204,n37192,n37205 );
   nor U38443 ( n37197,n37206,n37207 );
   nand U38444 ( n37207,n37208,n37209 );
   nand U38445 ( n37209,n37180,n37166 );
   nand U38446 ( n37208,n37168,n37210 );
   nand U38447 ( n37210,n37211,n37212 );
   nor U38448 ( n37206,n37213,n37214 );
   not U38449 ( n37214,n37215 );
   nor U38450 ( n37062,p2_state2_reg_0_,n37052 );
   nor U38451 ( n37060,n37216,n37217 );
   and U38452 ( n36671,n37218,n37219 );
   nor U38453 ( n37218,n37217,n28181 );
   nor U38454 ( n37221,n37222,n37223 );
   nand U38455 ( n37223,n37224,n37225 );
   nand U38456 ( n37225,n37226,n37227 );
   nand U38457 ( n37224,p2_instqueue_reg_15__7_,n37228 );
   nor U38458 ( n37222,n28197,n37230 );
   nor U38459 ( n37220,n37231,n37232 );
   nor U38460 ( n37232,n37233,n37234 );
   nor U38461 ( n37231,n37235,n28193 );
   nor U38462 ( n37238,n37239,n37240 );
   nand U38463 ( n37240,n37241,n37242 );
   nand U38464 ( n37242,n37243,n37227 );
   nand U38465 ( n37241,p2_instqueue_reg_15__6_,n37228 );
   nor U38466 ( n37239,n28203,n37230 );
   nor U38467 ( n37237,n37245,n37246 );
   nor U38468 ( n37246,n37247,n37234 );
   nor U38469 ( n37245,n37235,n28199 );
   nor U38470 ( n37250,n37251,n37252 );
   nand U38471 ( n37252,n37253,n37254 );
   nand U38472 ( n37254,n37255,n37227 );
   nand U38473 ( n37253,p2_instqueue_reg_15__5_,n37228 );
   nor U38474 ( n37251,n28210,n37230 );
   nor U38475 ( n37249,n37257,n37258 );
   nor U38476 ( n37258,n37259,n37234 );
   nor U38477 ( n37257,n37235,n28206 );
   nor U38478 ( n37262,n37263,n37264 );
   nand U38479 ( n37264,n37265,n37266 );
   nand U38480 ( n37266,n37267,n37227 );
   nand U38481 ( n37265,p2_instqueue_reg_15__4_,n37228 );
   nor U38482 ( n37263,n28218,n37230 );
   nor U38483 ( n37261,n37269,n37270 );
   nor U38484 ( n37270,n37271,n37234 );
   nor U38485 ( n37269,n37235,n28214 );
   nor U38486 ( n37274,n37275,n37276 );
   nand U38487 ( n37276,n37277,n37278 );
   nand U38488 ( n37278,n37279,n37227 );
   nand U38489 ( n37277,p2_instqueue_reg_15__3_,n37228 );
   nor U38490 ( n37275,n28230,n37230 );
   nor U38491 ( n37273,n37281,n37282 );
   nor U38492 ( n37282,n37283,n37234 );
   nor U38493 ( n37281,n37235,n28226 );
   nor U38494 ( n37286,n37287,n37288 );
   nand U38495 ( n37288,n37289,n37290 );
   nand U38496 ( n37290,n37291,n37227 );
   nand U38497 ( n37289,p2_instqueue_reg_15__2_,n37228 );
   nor U38498 ( n37287,n28248,n37230 );
   nor U38499 ( n37285,n37293,n37294 );
   nor U38500 ( n37294,n37295,n37234 );
   nor U38501 ( n37293,n37235,n28267 );
   nor U38502 ( n37298,n37299,n37300 );
   nand U38503 ( n37300,n37301,n37302 );
   nand U38504 ( n37302,n37303,n37227 );
   nand U38505 ( n37301,p2_instqueue_reg_15__1_,n37228 );
   nor U38506 ( n37299,n28272,n37230 );
   nor U38507 ( n37297,n37305,n37306 );
   nor U38508 ( n37306,n37307,n37234 );
   nor U38509 ( n37305,n37235,n28244 );
   nor U38510 ( n37310,n37311,n37312 );
   nand U38511 ( n37312,n37313,n37314 );
   nand U38512 ( n37314,n37315,n37227 );
   nand U38513 ( n37227,n37316,n37317 );
   nand U38514 ( n37317,p2_state2_reg_2_,n37318 );
   nand U38515 ( n37316,n37319,n37320 );
   nand U38516 ( n37313,p2_instqueue_reg_15__0_,n37228 );
   nand U38517 ( n37228,n37321,n37322 );
   nand U38518 ( n37322,p2_state2_reg_3_,n37235 );
   nor U38519 ( n37321,n37323,n37324 );
   nor U38520 ( n37324,n37325,n37326 );
   and U38521 ( n37325,n37318,n37327 );
   nand U38522 ( n37318,n37328,n37235 );
   nor U38523 ( n37323,n37320,n37329 );
   nand U38524 ( n37329,n37330,n37331 );
   nand U38525 ( n37330,n37332,n37333 );
   nand U38526 ( n37333,n37230,n37234 );
   nand U38527 ( n37320,n37235,n37334 );
   nand U38528 ( n37334,n37335,n37336 );
   nor U38529 ( n37311,n28328,n37230 );
   nand U38530 ( n37230,n37338,n36772 );
   nor U38531 ( n37338,n37339,n36697 );
   nor U38532 ( n37309,n37340,n37341 );
   nor U38533 ( n37341,n37342,n37234 );
   nand U38534 ( n37234,n36717,n37343 );
   not U38535 ( n36717,n36700 );
   nor U38536 ( n37340,n37235,n28324 );
   nand U38537 ( n37235,n37345,n37346 );
   nor U38538 ( n37348,n37349,n37350 );
   nand U38539 ( n37350,n37351,n37352 );
   nand U38540 ( n37352,n37226,n37353 );
   nand U38541 ( n37351,p2_instqueue_reg_14__7_,n37354 );
   nor U38542 ( n37349,n37229,n37355 );
   nor U38543 ( n37347,n37356,n37357 );
   nor U38544 ( n37357,n28193,n37358 );
   nor U38545 ( n37356,n37233,n37359 );
   nor U38546 ( n37361,n37362,n37363 );
   nand U38547 ( n37363,n37364,n37365 );
   nand U38548 ( n37365,n37243,n37353 );
   nand U38549 ( n37364,p2_instqueue_reg_14__6_,n37354 );
   nor U38550 ( n37362,n37244,n37355 );
   nor U38551 ( n37360,n37366,n37367 );
   nor U38552 ( n37367,n28199,n37358 );
   nor U38553 ( n37366,n37247,n37359 );
   nor U38554 ( n37369,n37370,n37371 );
   nand U38555 ( n37371,n37372,n37373 );
   nand U38556 ( n37373,n37255,n37353 );
   nand U38557 ( n37372,p2_instqueue_reg_14__5_,n37354 );
   nor U38558 ( n37370,n37256,n37355 );
   nor U38559 ( n37368,n37374,n37375 );
   nor U38560 ( n37375,n28206,n37358 );
   nor U38561 ( n37374,n37259,n37359 );
   nor U38562 ( n37377,n37378,n37379 );
   nand U38563 ( n37379,n37380,n37381 );
   nand U38564 ( n37381,n37267,n37353 );
   nand U38565 ( n37380,p2_instqueue_reg_14__4_,n37354 );
   nor U38566 ( n37378,n37268,n37355 );
   nor U38567 ( n37376,n37382,n37383 );
   nor U38568 ( n37383,n28214,n37358 );
   nor U38569 ( n37382,n37271,n37359 );
   nor U38570 ( n37385,n37386,n37387 );
   nand U38571 ( n37387,n37388,n37389 );
   nand U38572 ( n37389,n37279,n37353 );
   nand U38573 ( n37388,p2_instqueue_reg_14__3_,n37354 );
   nor U38574 ( n37386,n37280,n37355 );
   nor U38575 ( n37384,n37390,n37391 );
   nor U38576 ( n37391,n28226,n37358 );
   nor U38577 ( n37390,n37283,n37359 );
   nor U38578 ( n37393,n37394,n37395 );
   nand U38579 ( n37395,n37396,n37397 );
   nand U38580 ( n37397,n37291,n37353 );
   nand U38581 ( n37396,p2_instqueue_reg_14__2_,n37354 );
   nor U38582 ( n37394,n37292,n37355 );
   nor U38583 ( n37392,n37398,n37399 );
   nor U38584 ( n37399,n28267,n37358 );
   nor U38585 ( n37398,n37295,n37359 );
   nor U38586 ( n37401,n37402,n37403 );
   nand U38587 ( n37403,n37404,n37405 );
   nand U38588 ( n37405,n37303,n37353 );
   nand U38589 ( n37404,p2_instqueue_reg_14__1_,n37354 );
   nor U38590 ( n37402,n37304,n37355 );
   nor U38591 ( n37400,n37406,n37407 );
   nor U38592 ( n37407,n28244,n37358 );
   nor U38593 ( n37406,n37307,n37359 );
   nor U38594 ( n37409,n37410,n37411 );
   nand U38595 ( n37411,n37412,n37413 );
   nand U38596 ( n37413,n37315,n37353 );
   nand U38597 ( n37353,n37414,n37415 );
   nand U38598 ( n37415,n37335,n37319 );
   not U38599 ( n37335,n37416 );
   nand U38600 ( n37414,p2_state2_reg_2_,n37417 );
   nand U38601 ( n37412,p2_instqueue_reg_14__0_,n37354 );
   nand U38602 ( n37354,n37418,n37419 );
   nand U38603 ( n37419,p2_state2_reg_3_,n37358 );
   nor U38604 ( n37418,n37420,n37421 );
   nor U38605 ( n37421,n37422,n37326 );
   and U38606 ( n37422,n37417,n37327 );
   nand U38607 ( n37417,n37423,n37358 );
   nor U38608 ( n37420,n37424,n37425 );
   nand U38609 ( n37425,n37331,n37416 );
   nand U38610 ( n37416,n37426,n37427 );
   nor U38611 ( n37424,n37428,n36712 );
   and U38612 ( n37428,n37355,n37359 );
   nor U38613 ( n37410,n37337,n37355 );
   nand U38614 ( n37355,n37429,n37430 );
   nor U38615 ( n37408,n37431,n37432 );
   nor U38616 ( n37432,n28324,n37358 );
   nand U38617 ( n37358,n37433,n37345 );
   nor U38618 ( n37431,n37342,n37359 );
   nand U38619 ( n37359,n36687,n37434 );
   nor U38620 ( n37436,n37437,n37438 );
   nand U38621 ( n37438,n37439,n37440 );
   nand U38622 ( n37440,n37226,n37441 );
   nand U38623 ( n37439,p2_instqueue_reg_13__7_,n37442 );
   nor U38624 ( n37437,n28197,n37443 );
   nor U38625 ( n37435,n37444,n37445 );
   nor U38626 ( n37445,n28308,n37446 );
   nor U38627 ( n37444,n28193,n37447 );
   nor U38628 ( n37449,n37450,n37451 );
   nand U38629 ( n37451,n37452,n37453 );
   nand U38630 ( n37453,n37243,n37441 );
   nand U38631 ( n37452,p2_instqueue_reg_13__6_,n37442 );
   nor U38632 ( n37450,n28203,n37443 );
   nor U38633 ( n37448,n37454,n37455 );
   nor U38634 ( n37455,n28309,n37446 );
   nor U38635 ( n37454,n28199,n37447 );
   nor U38636 ( n37457,n37458,n37459 );
   nand U38637 ( n37459,n37460,n37461 );
   nand U38638 ( n37461,n37255,n37441 );
   nand U38639 ( n37460,p2_instqueue_reg_13__5_,n37442 );
   nor U38640 ( n37458,n28210,n37443 );
   nor U38641 ( n37456,n37462,n37463 );
   nor U38642 ( n37463,n28310,n37446 );
   nor U38643 ( n37462,n28206,n37447 );
   nor U38644 ( n37465,n37466,n37467 );
   nand U38645 ( n37467,n37468,n37469 );
   nand U38646 ( n37469,n37267,n37441 );
   nand U38647 ( n37468,p2_instqueue_reg_13__4_,n37442 );
   nor U38648 ( n37466,n28218,n37443 );
   nor U38649 ( n37464,n37470,n37471 );
   nor U38650 ( n37471,n28311,n37446 );
   nor U38651 ( n37470,n28214,n37447 );
   nor U38652 ( n37473,n37474,n37475 );
   nand U38653 ( n37475,n37476,n37477 );
   nand U38654 ( n37477,n37279,n37441 );
   nand U38655 ( n37476,p2_instqueue_reg_13__3_,n37442 );
   nor U38656 ( n37474,n28230,n37443 );
   nor U38657 ( n37472,n37478,n37479 );
   nor U38658 ( n37479,n28312,n37446 );
   nor U38659 ( n37478,n28226,n37447 );
   nor U38660 ( n37481,n37482,n37483 );
   nand U38661 ( n37483,n37484,n37485 );
   nand U38662 ( n37485,n37291,n37441 );
   nand U38663 ( n37484,p2_instqueue_reg_13__2_,n37442 );
   nor U38664 ( n37482,n28248,n37443 );
   nor U38665 ( n37480,n37486,n37487 );
   nor U38666 ( n37487,n28313,n37446 );
   nor U38667 ( n37486,n28267,n37447 );
   nor U38668 ( n37489,n37490,n37491 );
   nand U38669 ( n37491,n37492,n37493 );
   nand U38670 ( n37493,n37303,n37441 );
   nand U38671 ( n37492,p2_instqueue_reg_13__1_,n37442 );
   nor U38672 ( n37490,n28272,n37443 );
   nor U38673 ( n37488,n37494,n37495 );
   nor U38674 ( n37495,n28314,n37446 );
   nor U38675 ( n37494,n28244,n37447 );
   nor U38676 ( n37497,n37498,n37499 );
   nand U38677 ( n37499,n37500,n37501 );
   nand U38678 ( n37501,n37315,n37441 );
   nand U38679 ( n37441,n37502,n37503 );
   nand U38680 ( n37503,p2_state2_reg_2_,n37504 );
   nand U38681 ( n37502,n37505,n37319 );
   nand U38682 ( n37500,p2_instqueue_reg_13__0_,n37442 );
   nand U38683 ( n37442,n37506,n37507 );
   nand U38684 ( n37507,p2_state2_reg_3_,n37447 );
   nor U38685 ( n37506,n37508,n37509 );
   nor U38686 ( n37509,n37510,n37326 );
   and U38687 ( n37510,n37504,n37327 );
   nand U38688 ( n37504,n37511,n37447 );
   nor U38689 ( n37508,n37505,n37512 );
   nand U38690 ( n37512,n37513,n37331 );
   nand U38691 ( n37513,n37332,n37514 );
   nand U38692 ( n37514,n37443,n37446 );
   nand U38693 ( n37505,n37447,n37515 );
   nand U38694 ( n37515,n37516,n37336 );
   nor U38695 ( n37498,n28328,n37443 );
   nand U38696 ( n37443,n37429,n37517 );
   nor U38697 ( n37429,n36697,n36711 );
   nor U38698 ( n37496,n37518,n37519 );
   nor U38699 ( n37519,n28315,n37446 );
   nand U38700 ( n37446,n36688,n37434 );
   nor U38701 ( n37518,n28324,n37447 );
   nand U38702 ( n37447,n37520,n37345 );
   nor U38703 ( n37522,n37523,n37524 );
   nand U38704 ( n37524,n37525,n37526 );
   nand U38705 ( n37526,n37226,n37527 );
   nand U38706 ( n37525,p2_instqueue_reg_12__7_,n37528 );
   nor U38707 ( n37523,n28197,n37529 );
   nor U38708 ( n37521,n37530,n37531 );
   nor U38709 ( n37531,n37236,n37532 );
   nor U38710 ( n37530,n28308,n37533 );
   nor U38711 ( n37535,n37536,n37537 );
   nand U38712 ( n37537,n37538,n37539 );
   nand U38713 ( n37539,n37243,n37527 );
   nand U38714 ( n37538,p2_instqueue_reg_12__6_,n37528 );
   nor U38715 ( n37536,n28203,n37529 );
   nor U38716 ( n37534,n37540,n37541 );
   nor U38717 ( n37541,n37248,n37532 );
   nor U38718 ( n37540,n28309,n37533 );
   nor U38719 ( n37543,n37544,n37545 );
   nand U38720 ( n37545,n37546,n37547 );
   nand U38721 ( n37547,n37255,n37527 );
   nand U38722 ( n37546,p2_instqueue_reg_12__5_,n37528 );
   nor U38723 ( n37544,n28210,n37529 );
   nor U38724 ( n37542,n37548,n37549 );
   nor U38725 ( n37549,n37260,n37532 );
   nor U38726 ( n37548,n28310,n37533 );
   nor U38727 ( n37551,n37552,n37553 );
   nand U38728 ( n37553,n37554,n37555 );
   nand U38729 ( n37555,n37267,n37527 );
   nand U38730 ( n37554,p2_instqueue_reg_12__4_,n37528 );
   nor U38731 ( n37552,n28218,n37529 );
   nor U38732 ( n37550,n37556,n37557 );
   nor U38733 ( n37557,n37272,n37532 );
   nor U38734 ( n37556,n28311,n37533 );
   nor U38735 ( n37559,n37560,n37561 );
   nand U38736 ( n37561,n37562,n37563 );
   nand U38737 ( n37563,n37279,n37527 );
   nand U38738 ( n37562,p2_instqueue_reg_12__3_,n37528 );
   nor U38739 ( n37560,n28230,n37529 );
   nor U38740 ( n37558,n37564,n37565 );
   nor U38741 ( n37565,n37284,n37532 );
   nor U38742 ( n37564,n28312,n37533 );
   nor U38743 ( n37567,n37568,n37569 );
   nand U38744 ( n37569,n37570,n37571 );
   nand U38745 ( n37571,n37291,n37527 );
   nand U38746 ( n37570,p2_instqueue_reg_12__2_,n37528 );
   nor U38747 ( n37568,n28248,n37529 );
   nor U38748 ( n37566,n37572,n37573 );
   nor U38749 ( n37573,n37296,n37532 );
   nor U38750 ( n37572,n28313,n37533 );
   nor U38751 ( n37575,n37576,n37577 );
   nand U38752 ( n37577,n37578,n37579 );
   nand U38753 ( n37579,n37303,n37527 );
   nand U38754 ( n37578,p2_instqueue_reg_12__1_,n37528 );
   nor U38755 ( n37576,n28272,n37529 );
   nor U38756 ( n37574,n37580,n37581 );
   nor U38757 ( n37581,n37308,n37532 );
   nor U38758 ( n37580,n28314,n37533 );
   nor U38759 ( n37583,n37584,n37585 );
   nand U38760 ( n37585,n37586,n37587 );
   nand U38761 ( n37587,n37315,n37527 );
   nand U38762 ( n37527,n37588,n37589 );
   nand U38763 ( n37589,n37516,n37319 );
   not U38764 ( n37516,n37590 );
   nand U38765 ( n37588,p2_state2_reg_2_,n37591 );
   nand U38766 ( n37586,p2_instqueue_reg_12__0_,n37528 );
   nand U38767 ( n37528,n37592,n37593 );
   nand U38768 ( n37593,p2_state2_reg_3_,n37532 );
   nor U38769 ( n37592,n37594,n37595 );
   nor U38770 ( n37595,n37596,n37326 );
   and U38771 ( n37596,n37591,n37327 );
   nand U38772 ( n37591,n37597,n37532 );
   nor U38773 ( n37594,n37598,n37599 );
   nand U38774 ( n37599,n37331,n37590 );
   nand U38775 ( n37590,n37600,n37427 );
   nor U38776 ( n37598,n37601,n36712 );
   and U38777 ( n37601,n37529,n37533 );
   nor U38778 ( n37584,n28328,n37529 );
   nand U38779 ( n37529,n37602,n36772 );
   nor U38780 ( n37582,n37603,n37604 );
   nor U38781 ( n37604,n37344,n37532 );
   nand U38782 ( n37532,n37605,n37345 );
   nor U38783 ( n37345,n37606,n37607 );
   nor U38784 ( n37603,n28315,n37533 );
   nand U38785 ( n37533,n37608,n37434 );
   nor U38786 ( n37434,n37609,n36718 );
   nor U38787 ( n37611,n37612,n37613 );
   nand U38788 ( n37613,n37614,n37615 );
   nand U38789 ( n37615,n37226,n37616 );
   nand U38790 ( n37614,p2_instqueue_reg_11__7_,n37617 );
   nor U38791 ( n37612,n28197,n37618 );
   nor U38792 ( n37610,n37619,n37620 );
   nor U38793 ( n37620,n28308,n37621 );
   nor U38794 ( n37619,n37236,n37622 );
   nor U38795 ( n37624,n37625,n37626 );
   nand U38796 ( n37626,n37627,n37628 );
   nand U38797 ( n37628,n37243,n37616 );
   nand U38798 ( n37627,p2_instqueue_reg_11__6_,n37617 );
   nor U38799 ( n37625,n28203,n37618 );
   nor U38800 ( n37623,n37629,n37630 );
   nor U38801 ( n37630,n28309,n37621 );
   nor U38802 ( n37629,n37248,n37622 );
   nor U38803 ( n37632,n37633,n37634 );
   nand U38804 ( n37634,n37635,n37636 );
   nand U38805 ( n37636,n37255,n37616 );
   nand U38806 ( n37635,p2_instqueue_reg_11__5_,n37617 );
   nor U38807 ( n37633,n28210,n37618 );
   nor U38808 ( n37631,n37637,n37638 );
   nor U38809 ( n37638,n28310,n37621 );
   nor U38810 ( n37637,n37260,n37622 );
   nor U38811 ( n37640,n37641,n37642 );
   nand U38812 ( n37642,n37643,n37644 );
   nand U38813 ( n37644,n37267,n37616 );
   nand U38814 ( n37643,p2_instqueue_reg_11__4_,n37617 );
   nor U38815 ( n37641,n28218,n37618 );
   nor U38816 ( n37639,n37645,n37646 );
   nor U38817 ( n37646,n28311,n37621 );
   nor U38818 ( n37645,n37272,n37622 );
   nor U38819 ( n37648,n37649,n37650 );
   nand U38820 ( n37650,n37651,n37652 );
   nand U38821 ( n37652,n37279,n37616 );
   nand U38822 ( n37651,p2_instqueue_reg_11__3_,n37617 );
   nor U38823 ( n37649,n28230,n37618 );
   nor U38824 ( n37647,n37653,n37654 );
   nor U38825 ( n37654,n28312,n37621 );
   nor U38826 ( n37653,n37284,n37622 );
   nor U38827 ( n37656,n37657,n37658 );
   nand U38828 ( n37658,n37659,n37660 );
   nand U38829 ( n37660,n37291,n37616 );
   nand U38830 ( n37659,p2_instqueue_reg_11__2_,n37617 );
   nor U38831 ( n37657,n28248,n37618 );
   nor U38832 ( n37655,n37661,n37662 );
   nor U38833 ( n37662,n28313,n37621 );
   nor U38834 ( n37661,n37296,n37622 );
   nor U38835 ( n37664,n37665,n37666 );
   nand U38836 ( n37666,n37667,n37668 );
   nand U38837 ( n37668,n37303,n37616 );
   nand U38838 ( n37667,p2_instqueue_reg_11__1_,n37617 );
   nor U38839 ( n37665,n28272,n37618 );
   nor U38840 ( n37663,n37669,n37670 );
   nor U38841 ( n37670,n28314,n37621 );
   nor U38842 ( n37669,n37308,n37622 );
   nor U38843 ( n37672,n37673,n37674 );
   nand U38844 ( n37674,n37675,n37676 );
   nand U38845 ( n37676,n37315,n37616 );
   nand U38846 ( n37616,n37677,n37678 );
   nand U38847 ( n37678,p2_state2_reg_2_,n37679 );
   nand U38848 ( n37677,n37680,n37319 );
   nand U38849 ( n37675,p2_instqueue_reg_11__0_,n37617 );
   nand U38850 ( n37617,n37681,n37682 );
   nand U38851 ( n37682,p2_state2_reg_3_,n37622 );
   nor U38852 ( n37681,n37683,n37684 );
   nor U38853 ( n37684,n37685,n28303 );
   and U38854 ( n37685,n37679,n37327 );
   nand U38855 ( n37679,n37686,n37622 );
   nor U38856 ( n37683,n37680,n37687 );
   nand U38857 ( n37687,n37688,n37331 );
   nand U38858 ( n37688,n37332,n37689 );
   nand U38859 ( n37689,n37618,n37621 );
   nand U38860 ( n37680,n37622,n37690 );
   nand U38861 ( n37690,n37691,n37336 );
   nor U38862 ( n37673,n28328,n37618 );
   nand U38863 ( n37618,n37692,n37693 );
   nor U38864 ( n37671,n37694,n37695 );
   nor U38865 ( n37695,n28315,n37621 );
   nand U38866 ( n37621,n37696,n36702 );
   nor U38867 ( n37694,n37344,n37622 );
   nand U38868 ( n37622,n37697,n37346 );
   nor U38869 ( n37699,n37700,n37701 );
   nand U38870 ( n37701,n37702,n37703 );
   nand U38871 ( n37703,n37226,n37704 );
   nand U38872 ( n37702,p2_instqueue_reg_10__7_,n37705 );
   nor U38873 ( n37700,n28197,n37706 );
   nor U38874 ( n37698,n37707,n37708 );
   nor U38875 ( n37708,n37236,n37709 );
   nor U38876 ( n37707,n28308,n37710 );
   nor U38877 ( n37712,n37713,n37714 );
   nand U38878 ( n37714,n37715,n37716 );
   nand U38879 ( n37716,n37243,n37704 );
   nand U38880 ( n37715,p2_instqueue_reg_10__6_,n37705 );
   nor U38881 ( n37713,n28203,n37706 );
   nor U38882 ( n37711,n37717,n37718 );
   nor U38883 ( n37718,n37248,n37709 );
   nor U38884 ( n37717,n28309,n37710 );
   nor U38885 ( n37720,n37721,n37722 );
   nand U38886 ( n37722,n37723,n37724 );
   nand U38887 ( n37724,n37255,n37704 );
   nand U38888 ( n37723,p2_instqueue_reg_10__5_,n37705 );
   nor U38889 ( n37721,n28210,n37706 );
   nor U38890 ( n37719,n37725,n37726 );
   nor U38891 ( n37726,n37260,n37709 );
   nor U38892 ( n37725,n28310,n37710 );
   nor U38893 ( n37728,n37729,n37730 );
   nand U38894 ( n37730,n37731,n37732 );
   nand U38895 ( n37732,n37267,n37704 );
   nand U38896 ( n37731,p2_instqueue_reg_10__4_,n37705 );
   nor U38897 ( n37729,n28218,n37706 );
   nor U38898 ( n37727,n37733,n37734 );
   nor U38899 ( n37734,n37272,n37709 );
   nor U38900 ( n37733,n28311,n37710 );
   nor U38901 ( n37736,n37737,n37738 );
   nand U38902 ( n37738,n37739,n37740 );
   nand U38903 ( n37740,n37279,n37704 );
   nand U38904 ( n37739,p2_instqueue_reg_10__3_,n37705 );
   nor U38905 ( n37737,n28230,n37706 );
   nor U38906 ( n37735,n37741,n37742 );
   nor U38907 ( n37742,n37284,n37709 );
   nor U38908 ( n37741,n28312,n37710 );
   nor U38909 ( n37744,n37745,n37746 );
   nand U38910 ( n37746,n37747,n37748 );
   nand U38911 ( n37748,n37291,n37704 );
   nand U38912 ( n37747,p2_instqueue_reg_10__2_,n37705 );
   nor U38913 ( n37745,n28248,n37706 );
   nor U38914 ( n37743,n37749,n37750 );
   nor U38915 ( n37750,n37296,n37709 );
   nor U38916 ( n37749,n28313,n37710 );
   nor U38917 ( n37752,n37753,n37754 );
   nand U38918 ( n37754,n37755,n37756 );
   nand U38919 ( n37756,n37303,n37704 );
   nand U38920 ( n37755,p2_instqueue_reg_10__1_,n37705 );
   nor U38921 ( n37753,n28272,n37706 );
   nor U38922 ( n37751,n37757,n37758 );
   nor U38923 ( n37758,n37308,n37709 );
   nor U38924 ( n37757,n28314,n37710 );
   nor U38925 ( n37760,n37761,n37762 );
   nand U38926 ( n37762,n37763,n37764 );
   nand U38927 ( n37764,n37315,n37704 );
   nand U38928 ( n37704,n37765,n37766 );
   nand U38929 ( n37766,n37691,n37319 );
   not U38930 ( n37691,n37767 );
   nand U38931 ( n37765,p2_state2_reg_2_,n37768 );
   nand U38932 ( n37763,p2_instqueue_reg_10__0_,n37705 );
   nand U38933 ( n37705,n37769,n37770 );
   nand U38934 ( n37770,p2_state2_reg_3_,n37709 );
   nor U38935 ( n37769,n37771,n37772 );
   nor U38936 ( n37772,n37773,n28303 );
   and U38937 ( n37773,n37768,n37327 );
   nand U38938 ( n37768,n37774,n37709 );
   nor U38939 ( n37771,n37775,n37776 );
   nand U38940 ( n37776,n37331,n37767 );
   nand U38941 ( n37767,n37777,n37427 );
   nor U38942 ( n37775,n37778,n36712 );
   and U38943 ( n37778,n37706,n37710 );
   nor U38944 ( n37761,n28328,n37706 );
   nand U38945 ( n37706,n37692,n37430 );
   nor U38946 ( n37759,n37779,n37780 );
   nor U38947 ( n37780,n37344,n37709 );
   nand U38948 ( n37709,n37697,n37433 );
   nor U38949 ( n37779,n28315,n37710 );
   nand U38950 ( n37710,n37696,n36687 );
   nor U38951 ( n37782,n37783,n37784 );
   nand U38952 ( n37784,n37785,n37786 );
   nand U38953 ( n37786,n37226,n37787 );
   nand U38954 ( n37785,p2_instqueue_reg_9__7_,n37788 );
   nor U38955 ( n37783,n28197,n37789 );
   nor U38956 ( n37781,n37790,n37791 );
   nor U38957 ( n37791,n28308,n37792 );
   nor U38958 ( n37790,n28193,n37793 );
   nor U38959 ( n37795,n37796,n37797 );
   nand U38960 ( n37797,n37798,n37799 );
   nand U38961 ( n37799,n37243,n37787 );
   nand U38962 ( n37798,p2_instqueue_reg_9__6_,n37788 );
   nor U38963 ( n37796,n28203,n37789 );
   nor U38964 ( n37794,n37800,n37801 );
   nor U38965 ( n37801,n28309,n37792 );
   nor U38966 ( n37800,n28199,n37793 );
   nor U38967 ( n37803,n37804,n37805 );
   nand U38968 ( n37805,n37806,n37807 );
   nand U38969 ( n37807,n37255,n37787 );
   nand U38970 ( n37806,p2_instqueue_reg_9__5_,n37788 );
   nor U38971 ( n37804,n28210,n37789 );
   nor U38972 ( n37802,n37808,n37809 );
   nor U38973 ( n37809,n28310,n37792 );
   nor U38974 ( n37808,n28206,n37793 );
   nor U38975 ( n37811,n37812,n37813 );
   nand U38976 ( n37813,n37814,n37815 );
   nand U38977 ( n37815,n37267,n37787 );
   nand U38978 ( n37814,p2_instqueue_reg_9__4_,n37788 );
   nor U38979 ( n37812,n28218,n37789 );
   nor U38980 ( n37810,n37816,n37817 );
   nor U38981 ( n37817,n28311,n37792 );
   nor U38982 ( n37816,n28214,n37793 );
   nor U38983 ( n37819,n37820,n37821 );
   nand U38984 ( n37821,n37822,n37823 );
   nand U38985 ( n37823,n37279,n37787 );
   nand U38986 ( n37822,p2_instqueue_reg_9__3_,n37788 );
   nor U38987 ( n37820,n28230,n37789 );
   nor U38988 ( n37818,n37824,n37825 );
   nor U38989 ( n37825,n28312,n37792 );
   nor U38990 ( n37824,n28226,n37793 );
   nor U38991 ( n37827,n37828,n37829 );
   nand U38992 ( n37829,n37830,n37831 );
   nand U38993 ( n37831,n37291,n37787 );
   nand U38994 ( n37830,p2_instqueue_reg_9__2_,n37788 );
   nor U38995 ( n37828,n28248,n37789 );
   nor U38996 ( n37826,n37832,n37833 );
   nor U38997 ( n37833,n28313,n37792 );
   nor U38998 ( n37832,n28267,n37793 );
   nor U38999 ( n37835,n37836,n37837 );
   nand U39000 ( n37837,n37838,n37839 );
   nand U39001 ( n37839,n37303,n37787 );
   nand U39002 ( n37838,p2_instqueue_reg_9__1_,n37788 );
   nor U39003 ( n37836,n28272,n37789 );
   nor U39004 ( n37834,n37840,n37841 );
   nor U39005 ( n37841,n28314,n37792 );
   nor U39006 ( n37840,n28244,n37793 );
   nor U39007 ( n37843,n37844,n37845 );
   nand U39008 ( n37845,n37846,n37847 );
   nand U39009 ( n37847,n37315,n37787 );
   nand U39010 ( n37787,n37848,n37849 );
   nand U39011 ( n37849,p2_state2_reg_2_,n37850 );
   nand U39012 ( n37848,n37851,n37319 );
   nand U39013 ( n37846,p2_instqueue_reg_9__0_,n37788 );
   nand U39014 ( n37788,n37852,n37853 );
   nand U39015 ( n37853,p2_state2_reg_3_,n37793 );
   nor U39016 ( n37852,n37854,n37855 );
   nor U39017 ( n37855,n37856,n37326 );
   and U39018 ( n37856,n37850,n37327 );
   nand U39019 ( n37850,n37857,n37793 );
   nor U39020 ( n37854,n37851,n37858 );
   nand U39021 ( n37858,n37859,n37331 );
   nand U39022 ( n37859,n37332,n37860 );
   nand U39023 ( n37860,n37789,n37792 );
   nand U39024 ( n37851,n37793,n37861 );
   nand U39025 ( n37861,n37862,n37336 );
   nor U39026 ( n37844,n28328,n37789 );
   nand U39027 ( n37789,n37692,n37517 );
   nor U39028 ( n37842,n37863,n37864 );
   nor U39029 ( n37864,n28315,n37792 );
   nand U39030 ( n37792,n37696,n36688 );
   nor U39031 ( n37863,n28324,n37793 );
   nand U39032 ( n37793,n37697,n37520 );
   nor U39033 ( n37866,n37867,n37868 );
   nand U39034 ( n37868,n37869,n37870 );
   nand U39035 ( n37870,n37226,n37871 );
   nand U39036 ( n37869,p2_instqueue_reg_8__7_,n37872 );
   nor U39037 ( n37867,n37229,n37873 );
   nor U39038 ( n37865,n37874,n37875 );
   nor U39039 ( n37875,n28193,n37876 );
   nor U39040 ( n37874,n37233,n37877 );
   nor U39041 ( n37879,n37880,n37881 );
   nand U39042 ( n37881,n37882,n37883 );
   nand U39043 ( n37883,n37243,n37871 );
   nand U39044 ( n37882,p2_instqueue_reg_8__6_,n37872 );
   nor U39045 ( n37880,n37244,n37873 );
   nor U39046 ( n37878,n37884,n37885 );
   nor U39047 ( n37885,n28199,n37876 );
   nor U39048 ( n37884,n37247,n37877 );
   nor U39049 ( n37887,n37888,n37889 );
   nand U39050 ( n37889,n37890,n37891 );
   nand U39051 ( n37891,n37255,n37871 );
   nand U39052 ( n37890,p2_instqueue_reg_8__5_,n37872 );
   nor U39053 ( n37888,n37256,n37873 );
   nor U39054 ( n37886,n37892,n37893 );
   nor U39055 ( n37893,n28206,n37876 );
   nor U39056 ( n37892,n37259,n37877 );
   nor U39057 ( n37895,n37896,n37897 );
   nand U39058 ( n37897,n37898,n37899 );
   nand U39059 ( n37899,n37267,n37871 );
   nand U39060 ( n37898,p2_instqueue_reg_8__4_,n37872 );
   nor U39061 ( n37896,n37268,n37873 );
   nor U39062 ( n37894,n37900,n37901 );
   nor U39063 ( n37901,n28214,n37876 );
   nor U39064 ( n37900,n37271,n37877 );
   nor U39065 ( n37903,n37904,n37905 );
   nand U39066 ( n37905,n37906,n37907 );
   nand U39067 ( n37907,n37279,n37871 );
   nand U39068 ( n37906,p2_instqueue_reg_8__3_,n37872 );
   nor U39069 ( n37904,n37280,n37873 );
   nor U39070 ( n37902,n37908,n37909 );
   nor U39071 ( n37909,n28226,n37876 );
   nor U39072 ( n37908,n37283,n37877 );
   nor U39073 ( n37911,n37912,n37913 );
   nand U39074 ( n37913,n37914,n37915 );
   nand U39075 ( n37915,n37291,n37871 );
   nand U39076 ( n37914,p2_instqueue_reg_8__2_,n37872 );
   nor U39077 ( n37912,n37292,n37873 );
   nor U39078 ( n37910,n37916,n37917 );
   nor U39079 ( n37917,n28267,n37876 );
   nor U39080 ( n37916,n37295,n37877 );
   nor U39081 ( n37919,n37920,n37921 );
   nand U39082 ( n37921,n37922,n37923 );
   nand U39083 ( n37923,n37303,n37871 );
   nand U39084 ( n37922,p2_instqueue_reg_8__1_,n37872 );
   nor U39085 ( n37920,n37304,n37873 );
   nor U39086 ( n37918,n37924,n37925 );
   nor U39087 ( n37925,n28244,n37876 );
   nor U39088 ( n37924,n37307,n37877 );
   nor U39089 ( n37927,n37928,n37929 );
   nand U39090 ( n37929,n37930,n37931 );
   nand U39091 ( n37931,n37315,n37871 );
   nand U39092 ( n37871,n37932,n37933 );
   nand U39093 ( n37933,n37862,n37319 );
   not U39094 ( n37862,n37934 );
   nand U39095 ( n37932,p2_state2_reg_2_,n37935 );
   nand U39096 ( n37930,p2_instqueue_reg_8__0_,n37872 );
   nand U39097 ( n37872,n37936,n37937 );
   nand U39098 ( n37937,p2_state2_reg_3_,n37876 );
   nor U39099 ( n37936,n37938,n37939 );
   nor U39100 ( n37939,n37940,n37326 );
   and U39101 ( n37940,n37935,n37327 );
   nand U39102 ( n37935,n37941,n37876 );
   nor U39103 ( n37938,n37942,n37943 );
   nand U39104 ( n37943,n37331,n37934 );
   nand U39105 ( n37934,n37944,n37427 );
   nor U39106 ( n37942,n37945,n36712 );
   and U39107 ( n37945,n37873,n37877 );
   nor U39108 ( n37928,n37337,n37873 );
   nand U39109 ( n37873,n37946,n37692 );
   nor U39110 ( n37926,n37947,n37948 );
   nor U39111 ( n37948,n28324,n37876 );
   nand U39112 ( n37876,n37697,n37605 );
   nor U39113 ( n37947,n37342,n37877 );
   nand U39114 ( n37877,n37696,n37608 );
   nor U39115 ( n37696,n36701,n36718 );
   not U39116 ( n36718,n37343 );
   nor U39117 ( n37950,n37951,n37952 );
   nand U39118 ( n37952,n37953,n37954 );
   nand U39119 ( n37954,n37226,n37955 );
   nand U39120 ( n37953,p2_instqueue_reg_7__7_,n37956 );
   nor U39121 ( n37951,n37233,n37957 );
   nor U39122 ( n37949,n37958,n37959 );
   nor U39123 ( n37959,n37229,n37960 );
   nor U39124 ( n37958,n37236,n37961 );
   nor U39125 ( n37963,n37964,n37965 );
   nand U39126 ( n37965,n37966,n37967 );
   nand U39127 ( n37967,n37243,n37955 );
   nand U39128 ( n37966,p2_instqueue_reg_7__6_,n37956 );
   nor U39129 ( n37964,n37247,n37957 );
   nor U39130 ( n37962,n37968,n37969 );
   nor U39131 ( n37969,n37244,n37960 );
   nor U39132 ( n37968,n37248,n37961 );
   nor U39133 ( n37971,n37972,n37973 );
   nand U39134 ( n37973,n37974,n37975 );
   nand U39135 ( n37975,n37255,n37955 );
   nand U39136 ( n37974,p2_instqueue_reg_7__5_,n37956 );
   nor U39137 ( n37972,n37259,n37957 );
   nor U39138 ( n37970,n37976,n37977 );
   nor U39139 ( n37977,n37256,n37960 );
   nor U39140 ( n37976,n37260,n37961 );
   nor U39141 ( n37979,n37980,n37981 );
   nand U39142 ( n37981,n37982,n37983 );
   nand U39143 ( n37983,n37267,n37955 );
   nand U39144 ( n37982,p2_instqueue_reg_7__4_,n37956 );
   nor U39145 ( n37980,n37271,n37957 );
   nor U39146 ( n37978,n37984,n37985 );
   nor U39147 ( n37985,n37268,n37960 );
   nor U39148 ( n37984,n37272,n37961 );
   nor U39149 ( n37987,n37988,n37989 );
   nand U39150 ( n37989,n37990,n37991 );
   nand U39151 ( n37991,n37279,n37955 );
   nand U39152 ( n37990,p2_instqueue_reg_7__3_,n37956 );
   nor U39153 ( n37988,n37283,n37957 );
   nor U39154 ( n37986,n37992,n37993 );
   nor U39155 ( n37993,n37280,n37960 );
   nor U39156 ( n37992,n37284,n37961 );
   nor U39157 ( n37995,n37996,n37997 );
   nand U39158 ( n37997,n37998,n37999 );
   nand U39159 ( n37999,n37291,n37955 );
   nand U39160 ( n37998,p2_instqueue_reg_7__2_,n37956 );
   nor U39161 ( n37996,n37295,n37957 );
   nor U39162 ( n37994,n38000,n38001 );
   nor U39163 ( n38001,n37292,n37960 );
   nor U39164 ( n38000,n37296,n37961 );
   nor U39165 ( n38003,n38004,n38005 );
   nand U39166 ( n38005,n38006,n38007 );
   nand U39167 ( n38007,n37303,n37955 );
   nand U39168 ( n38006,p2_instqueue_reg_7__1_,n37956 );
   nor U39169 ( n38004,n37307,n37957 );
   nor U39170 ( n38002,n38008,n38009 );
   nor U39171 ( n38009,n37304,n37960 );
   nor U39172 ( n38008,n37308,n37961 );
   nor U39173 ( n38011,n38012,n38013 );
   nand U39174 ( n38013,n38014,n38015 );
   nand U39175 ( n38015,n37315,n37955 );
   nand U39176 ( n37955,n38016,n38017 );
   nand U39177 ( n38017,p2_state2_reg_2_,n38018 );
   nand U39178 ( n38018,n37961,n38019 );
   nand U39179 ( n38016,n38020,n37319 );
   nand U39180 ( n38014,p2_instqueue_reg_7__0_,n37956 );
   nand U39181 ( n37956,n38021,n37327 );
   nor U39182 ( n38021,n38022,n38023 );
   nor U39183 ( n38023,n38024,n38025 );
   nor U39184 ( n38025,n38026,p2_state2_reg_3_ );
   nor U39185 ( n38026,n37326,n38027 );
   not U39186 ( n38027,n38019 );
   nor U39187 ( n38022,n38020,n38028 );
   nand U39188 ( n38028,n38029,n37331 );
   nand U39189 ( n38029,n37332,n38030 );
   nand U39190 ( n38030,n37960,n37957 );
   nand U39191 ( n38020,n37961,n38031 );
   nand U39192 ( n38031,n38032,n37426 );
   nor U39193 ( n38012,n37342,n37957 );
   not U39194 ( n37957,n36716 );
   nor U39195 ( n36716,n36700,n37343 );
   nand U39196 ( n36700,n36702,n36701 );
   nor U39197 ( n38010,n38033,n38034 );
   nor U39198 ( n38034,n37337,n37960 );
   nor U39199 ( n38033,n37344,n37961 );
   nor U39200 ( n38036,n38037,n38038 );
   nand U39201 ( n38038,n38039,n38040 );
   nand U39202 ( n38040,n37226,n38041 );
   nand U39203 ( n38039,p2_instqueue_reg_6__7_,n38042 );
   nor U39204 ( n38037,n37229,n38043 );
   nor U39205 ( n38035,n38044,n38045 );
   nor U39206 ( n38045,n28193,n38046 );
   nor U39207 ( n38044,n37233,n38047 );
   nor U39208 ( n38049,n38050,n38051 );
   nand U39209 ( n38051,n38052,n38053 );
   nand U39210 ( n38053,n37243,n38041 );
   nand U39211 ( n38052,p2_instqueue_reg_6__6_,n38042 );
   nor U39212 ( n38050,n37244,n38043 );
   nor U39213 ( n38048,n38054,n38055 );
   nor U39214 ( n38055,n28199,n38046 );
   nor U39215 ( n38054,n37247,n38047 );
   nor U39216 ( n38057,n38058,n38059 );
   nand U39217 ( n38059,n38060,n38061 );
   nand U39218 ( n38061,n37255,n38041 );
   nand U39219 ( n38060,p2_instqueue_reg_6__5_,n38042 );
   nor U39220 ( n38058,n37256,n38043 );
   nor U39221 ( n38056,n38062,n38063 );
   nor U39222 ( n38063,n28206,n38046 );
   nor U39223 ( n38062,n37259,n38047 );
   nor U39224 ( n38065,n38066,n38067 );
   nand U39225 ( n38067,n38068,n38069 );
   nand U39226 ( n38069,n37267,n38041 );
   nand U39227 ( n38068,p2_instqueue_reg_6__4_,n38042 );
   nor U39228 ( n38066,n37268,n38043 );
   nor U39229 ( n38064,n38070,n38071 );
   nor U39230 ( n38071,n28214,n38046 );
   nor U39231 ( n38070,n37271,n38047 );
   nor U39232 ( n38073,n38074,n38075 );
   nand U39233 ( n38075,n38076,n38077 );
   nand U39234 ( n38077,n37279,n38041 );
   nand U39235 ( n38076,p2_instqueue_reg_6__3_,n38042 );
   nor U39236 ( n38074,n37280,n38043 );
   nor U39237 ( n38072,n38078,n38079 );
   nor U39238 ( n38079,n28226,n38046 );
   nor U39239 ( n38078,n37283,n38047 );
   nor U39240 ( n38081,n38082,n38083 );
   nand U39241 ( n38083,n38084,n38085 );
   nand U39242 ( n38085,n37291,n38041 );
   nand U39243 ( n38084,p2_instqueue_reg_6__2_,n38042 );
   nor U39244 ( n38082,n37292,n38043 );
   nor U39245 ( n38080,n38086,n38087 );
   nor U39246 ( n38087,n28267,n38046 );
   nor U39247 ( n38086,n37295,n38047 );
   nor U39248 ( n38089,n38090,n38091 );
   nand U39249 ( n38091,n38092,n38093 );
   nand U39250 ( n38093,n37303,n38041 );
   nand U39251 ( n38092,p2_instqueue_reg_6__1_,n38042 );
   nor U39252 ( n38090,n37304,n38043 );
   nor U39253 ( n38088,n38094,n38095 );
   nor U39254 ( n38095,n28244,n38046 );
   nor U39255 ( n38094,n37307,n38047 );
   nor U39256 ( n38097,n38098,n38099 );
   nand U39257 ( n38099,n38100,n38101 );
   nand U39258 ( n38101,n37315,n38041 );
   nand U39259 ( n38041,n38102,n38103 );
   nand U39260 ( n38103,n38104,n37426 );
   nand U39261 ( n38102,p2_state2_reg_2_,n38105 );
   nand U39262 ( n38100,p2_instqueue_reg_6__0_,n38042 );
   nand U39263 ( n38042,n38106,n38107 );
   nand U39264 ( n38107,p2_state2_reg_3_,n38046 );
   nor U39265 ( n38106,n38108,n38109 );
   nor U39266 ( n38109,n38110,n37326 );
   and U39267 ( n38110,n37327,n38105 );
   nand U39268 ( n38105,n38111,n38046 );
   nor U39269 ( n38108,n38112,n38113 );
   nand U39270 ( n38113,n38114,n37331 );
   nand U39271 ( n38114,n38115,n37426 );
   nor U39272 ( n37426,n38116,n38117 );
   nor U39273 ( n38112,n38118,n36712 );
   and U39274 ( n38118,n38043,n38047 );
   nor U39275 ( n38098,n37337,n38043 );
   nand U39276 ( n38043,n38119,n37430 );
   nor U39277 ( n38096,n38120,n38121 );
   nor U39278 ( n38121,n28324,n38046 );
   nand U39279 ( n38046,n37433,n38122 );
   nor U39280 ( n38120,n37342,n38047 );
   nand U39281 ( n38047,n38123,n36687 );
   nor U39282 ( n38125,n38126,n38127 );
   nand U39283 ( n38127,n38128,n38129 );
   nand U39284 ( n38129,n37226,n38130 );
   nand U39285 ( n38128,p2_instqueue_reg_5__7_,n38131 );
   nor U39286 ( n38126,n37229,n38132 );
   nor U39287 ( n38124,n38133,n38134 );
   nor U39288 ( n38134,n37233,n38135 );
   nor U39289 ( n38133,n37236,n38136 );
   nor U39290 ( n38138,n38139,n38140 );
   nand U39291 ( n38140,n38141,n38142 );
   nand U39292 ( n38142,n37243,n38130 );
   nand U39293 ( n38141,p2_instqueue_reg_5__6_,n38131 );
   nor U39294 ( n38139,n37244,n38132 );
   nor U39295 ( n38137,n38143,n38144 );
   nor U39296 ( n38144,n37247,n38135 );
   nor U39297 ( n38143,n37248,n38136 );
   nor U39298 ( n38146,n38147,n38148 );
   nand U39299 ( n38148,n38149,n38150 );
   nand U39300 ( n38150,n37255,n38130 );
   nand U39301 ( n38149,p2_instqueue_reg_5__5_,n38131 );
   nor U39302 ( n38147,n37256,n38132 );
   nor U39303 ( n38145,n38151,n38152 );
   nor U39304 ( n38152,n37259,n38135 );
   nor U39305 ( n38151,n37260,n38136 );
   nor U39306 ( n38154,n38155,n38156 );
   nand U39307 ( n38156,n38157,n38158 );
   nand U39308 ( n38158,n37267,n38130 );
   nand U39309 ( n38157,p2_instqueue_reg_5__4_,n38131 );
   nor U39310 ( n38155,n37268,n38132 );
   nor U39311 ( n38153,n38159,n38160 );
   nor U39312 ( n38160,n37271,n38135 );
   nor U39313 ( n38159,n37272,n38136 );
   nor U39314 ( n38162,n38163,n38164 );
   nand U39315 ( n38164,n38165,n38166 );
   nand U39316 ( n38166,n37279,n38130 );
   nand U39317 ( n38165,p2_instqueue_reg_5__3_,n38131 );
   nor U39318 ( n38163,n37280,n38132 );
   nor U39319 ( n38161,n38167,n38168 );
   nor U39320 ( n38168,n37283,n38135 );
   nor U39321 ( n38167,n37284,n38136 );
   nor U39322 ( n38170,n38171,n38172 );
   nand U39323 ( n38172,n38173,n38174 );
   nand U39324 ( n38174,n37291,n38130 );
   nand U39325 ( n38173,p2_instqueue_reg_5__2_,n38131 );
   nor U39326 ( n38171,n37292,n38132 );
   nor U39327 ( n38169,n38175,n38176 );
   nor U39328 ( n38176,n37295,n38135 );
   nor U39329 ( n38175,n37296,n38136 );
   nor U39330 ( n38178,n38179,n38180 );
   nand U39331 ( n38180,n38181,n38182 );
   nand U39332 ( n38182,n37303,n38130 );
   nand U39333 ( n38181,p2_instqueue_reg_5__1_,n38131 );
   nor U39334 ( n38179,n37304,n38132 );
   nor U39335 ( n38177,n38183,n38184 );
   nor U39336 ( n38184,n37307,n38135 );
   nor U39337 ( n38183,n37308,n38136 );
   nor U39338 ( n38186,n38187,n38188 );
   nand U39339 ( n38188,n38189,n38190 );
   nand U39340 ( n38190,n37315,n38130 );
   nand U39341 ( n38130,n38191,n38192 );
   nand U39342 ( n38192,p2_state2_reg_2_,n38193 );
   nand U39343 ( n38191,n38194,n37319 );
   nand U39344 ( n38189,p2_instqueue_reg_5__0_,n38131 );
   nand U39345 ( n38131,n38195,n38196 );
   nand U39346 ( n38196,p2_state2_reg_3_,n38136 );
   nor U39347 ( n38195,n38197,n38198 );
   nor U39348 ( n38198,n38199,n37326 );
   and U39349 ( n38199,n37327,n38193 );
   nand U39350 ( n38193,n38200,n38136 );
   nor U39351 ( n38197,n38194,n38201 );
   nand U39352 ( n38201,n38202,n37331 );
   nand U39353 ( n38202,n37332,n38203 );
   nand U39354 ( n38203,n38132,n38135 );
   nand U39355 ( n38194,n38136,n38204 );
   nand U39356 ( n38204,n38032,n37600 );
   nor U39357 ( n38187,n37337,n38132 );
   nand U39358 ( n38132,n38119,n37517 );
   nor U39359 ( n38119,n36772,n36697 );
   nor U39360 ( n38185,n38205,n38206 );
   nor U39361 ( n38206,n37342,n38135 );
   nand U39362 ( n38135,n38123,n36688 );
   nor U39363 ( n38205,n37344,n38136 );
   nand U39364 ( n38136,n37520,n38122 );
   nor U39365 ( n38208,n38209,n38210 );
   nand U39366 ( n38210,n38211,n38212 );
   nand U39367 ( n38212,n37226,n38213 );
   nand U39368 ( n38211,p2_instqueue_reg_4__7_,n38214 );
   nor U39369 ( n38209,n37229,n38215 );
   nor U39370 ( n38207,n38216,n38217 );
   nor U39371 ( n38217,n37236,n38218 );
   nor U39372 ( n38216,n37233,n38219 );
   nor U39373 ( n38221,n38222,n38223 );
   nand U39374 ( n38223,n38224,n38225 );
   nand U39375 ( n38225,n37243,n38213 );
   nand U39376 ( n38224,p2_instqueue_reg_4__6_,n38214 );
   nor U39377 ( n38222,n37244,n38215 );
   nor U39378 ( n38220,n38226,n38227 );
   nor U39379 ( n38227,n37248,n38218 );
   nor U39380 ( n38226,n37247,n38219 );
   nor U39381 ( n38229,n38230,n38231 );
   nand U39382 ( n38231,n38232,n38233 );
   nand U39383 ( n38233,n37255,n38213 );
   nand U39384 ( n38232,p2_instqueue_reg_4__5_,n38214 );
   nor U39385 ( n38230,n37256,n38215 );
   nor U39386 ( n38228,n38234,n38235 );
   nor U39387 ( n38235,n37260,n38218 );
   nor U39388 ( n38234,n37259,n38219 );
   nor U39389 ( n38237,n38238,n38239 );
   nand U39390 ( n38239,n38240,n38241 );
   nand U39391 ( n38241,n37267,n38213 );
   nand U39392 ( n38240,p2_instqueue_reg_4__4_,n38214 );
   nor U39393 ( n38238,n37268,n38215 );
   nor U39394 ( n38236,n38242,n38243 );
   nor U39395 ( n38243,n37272,n38218 );
   nor U39396 ( n38242,n37271,n38219 );
   nor U39397 ( n38245,n38246,n38247 );
   nand U39398 ( n38247,n38248,n38249 );
   nand U39399 ( n38249,n37279,n38213 );
   nand U39400 ( n38248,p2_instqueue_reg_4__3_,n38214 );
   nor U39401 ( n38246,n37280,n38215 );
   nor U39402 ( n38244,n38250,n38251 );
   nor U39403 ( n38251,n37284,n38218 );
   nor U39404 ( n38250,n37283,n38219 );
   nor U39405 ( n38253,n38254,n38255 );
   nand U39406 ( n38255,n38256,n38257 );
   nand U39407 ( n38257,n37291,n38213 );
   nand U39408 ( n38256,p2_instqueue_reg_4__2_,n38214 );
   nor U39409 ( n38254,n37292,n38215 );
   nor U39410 ( n38252,n38258,n38259 );
   nor U39411 ( n38259,n37296,n38218 );
   nor U39412 ( n38258,n37295,n38219 );
   nor U39413 ( n38261,n38262,n38263 );
   nand U39414 ( n38263,n38264,n38265 );
   nand U39415 ( n38265,n37303,n38213 );
   nand U39416 ( n38264,p2_instqueue_reg_4__1_,n38214 );
   nor U39417 ( n38262,n37304,n38215 );
   nor U39418 ( n38260,n38266,n38267 );
   nor U39419 ( n38267,n37308,n38218 );
   nor U39420 ( n38266,n37307,n38219 );
   nor U39421 ( n38269,n38270,n38271 );
   nand U39422 ( n38271,n38272,n38273 );
   nand U39423 ( n38273,n37315,n38213 );
   nand U39424 ( n38213,n38274,n38275 );
   nand U39425 ( n38275,n38104,n37600 );
   nand U39426 ( n38274,p2_state2_reg_2_,n38276 );
   nand U39427 ( n38272,p2_instqueue_reg_4__0_,n38214 );
   nand U39428 ( n38214,n38277,n38278 );
   nand U39429 ( n38278,p2_state2_reg_3_,n38218 );
   nor U39430 ( n38277,n38279,n38280 );
   nor U39431 ( n38280,n38281,n37326 );
   and U39432 ( n38281,n37327,n38276 );
   nand U39433 ( n38276,n38282,n38218 );
   nor U39434 ( n38279,n38283,n38284 );
   nand U39435 ( n38284,n38285,n37331 );
   nand U39436 ( n38285,n38115,n37600 );
   nor U39437 ( n37600,n38286,n38116 );
   nor U39438 ( n38283,n38287,n36712 );
   and U39439 ( n38287,n38215,n38219 );
   nor U39440 ( n38270,n37337,n38215 );
   nand U39441 ( n38215,n37602,n36711 );
   and U39442 ( n37602,n37946,n36752 );
   nor U39443 ( n38268,n38288,n38289 );
   nor U39444 ( n38289,n37344,n38218 );
   nand U39445 ( n38218,n37605,n38122 );
   nor U39446 ( n38288,n37342,n38219 );
   nand U39447 ( n38219,n38123,n37608 );
   nor U39448 ( n38123,n37343,n37609 );
   not U39449 ( n37609,n36701 );
   nor U39450 ( n38291,n38292,n38293 );
   nand U39451 ( n38293,n38294,n38295 );
   nand U39452 ( n38295,n37226,n38296 );
   nand U39453 ( n38294,p2_instqueue_reg_3__7_,n38297 );
   nor U39454 ( n38292,n37229,n38298 );
   nor U39455 ( n38290,n38299,n38300 );
   nor U39456 ( n38300,n37233,n38301 );
   nor U39457 ( n38299,n37236,n38302 );
   nor U39458 ( n38304,n38305,n38306 );
   nand U39459 ( n38306,n38307,n38308 );
   nand U39460 ( n38308,n37243,n38296 );
   nand U39461 ( n38307,p2_instqueue_reg_3__6_,n38297 );
   nor U39462 ( n38305,n37244,n38298 );
   nor U39463 ( n38303,n38309,n38310 );
   nor U39464 ( n38310,n37247,n38301 );
   nor U39465 ( n38309,n37248,n38302 );
   nor U39466 ( n38312,n38313,n38314 );
   nand U39467 ( n38314,n38315,n38316 );
   nand U39468 ( n38316,n37255,n38296 );
   nand U39469 ( n38315,p2_instqueue_reg_3__5_,n38297 );
   nor U39470 ( n38313,n37256,n38298 );
   nor U39471 ( n38311,n38317,n38318 );
   nor U39472 ( n38318,n37259,n38301 );
   nor U39473 ( n38317,n37260,n38302 );
   nor U39474 ( n38320,n38321,n38322 );
   nand U39475 ( n38322,n38323,n38324 );
   nand U39476 ( n38324,n37267,n38296 );
   nand U39477 ( n38323,p2_instqueue_reg_3__4_,n38297 );
   nor U39478 ( n38321,n37268,n38298 );
   nor U39479 ( n38319,n38325,n38326 );
   nor U39480 ( n38326,n37271,n38301 );
   nor U39481 ( n38325,n37272,n38302 );
   nor U39482 ( n38328,n38329,n38330 );
   nand U39483 ( n38330,n38331,n38332 );
   nand U39484 ( n38332,n37279,n38296 );
   nand U39485 ( n38331,p2_instqueue_reg_3__3_,n38297 );
   nor U39486 ( n38329,n37280,n38298 );
   nor U39487 ( n38327,n38333,n38334 );
   nor U39488 ( n38334,n37283,n38301 );
   nor U39489 ( n38333,n37284,n38302 );
   nor U39490 ( n38336,n38337,n38338 );
   nand U39491 ( n38338,n38339,n38340 );
   nand U39492 ( n38340,n37291,n38296 );
   nand U39493 ( n38339,p2_instqueue_reg_3__2_,n38297 );
   nor U39494 ( n38337,n37292,n38298 );
   nor U39495 ( n38335,n38341,n38342 );
   nor U39496 ( n38342,n37295,n38301 );
   nor U39497 ( n38341,n37296,n38302 );
   nor U39498 ( n38344,n38345,n38346 );
   nand U39499 ( n38346,n38347,n38348 );
   nand U39500 ( n38348,n37303,n38296 );
   nand U39501 ( n38347,p2_instqueue_reg_3__1_,n38297 );
   nor U39502 ( n38345,n37304,n38298 );
   nor U39503 ( n38343,n38349,n38350 );
   nor U39504 ( n38350,n37307,n38301 );
   nor U39505 ( n38349,n37308,n38302 );
   nor U39506 ( n38352,n38353,n38354 );
   nand U39507 ( n38354,n38355,n38356 );
   nand U39508 ( n38356,n37315,n38296 );
   nand U39509 ( n38296,n38357,n38358 );
   nand U39510 ( n38358,p2_state2_reg_2_,n38359 );
   nand U39511 ( n38357,n38360,n37319 );
   nand U39512 ( n38355,p2_instqueue_reg_3__0_,n38297 );
   nand U39513 ( n38297,n38361,n38362 );
   nand U39514 ( n38362,p2_state2_reg_3_,n38302 );
   nor U39515 ( n38361,n38363,n38364 );
   nor U39516 ( n38364,n38365,n37326 );
   and U39517 ( n38365,n37327,n38359 );
   nand U39518 ( n38359,n38366,n38302 );
   nor U39519 ( n38363,n38360,n38367 );
   nand U39520 ( n38367,n38368,n37331 );
   nand U39521 ( n38368,n37332,n38369 );
   nand U39522 ( n38369,n38298,n38301 );
   nand U39523 ( n38360,n38302,n38370 );
   nand U39524 ( n38370,n38032,n37777 );
   nor U39525 ( n38353,n37337,n38298 );
   nand U39526 ( n38298,n38371,n37693 );
   nor U39527 ( n38351,n38372,n38373 );
   nor U39528 ( n38373,n37342,n38301 );
   nand U39529 ( n38301,n38374,n36702 );
   nor U39530 ( n36702,n36729,n38375 );
   nor U39531 ( n38372,n37344,n38302 );
   nand U39532 ( n38302,n38376,n37346 );
   nor U39533 ( n38378,n38379,n38380 );
   nand U39534 ( n38380,n38381,n38382 );
   nand U39535 ( n38382,n37226,n38383 );
   nand U39536 ( n38381,p2_instqueue_reg_2__7_,n38384 );
   nor U39537 ( n38379,n37229,n38385 );
   nor U39538 ( n38377,n38386,n38387 );
   nor U39539 ( n38387,n37236,n38388 );
   nor U39540 ( n38386,n37233,n38389 );
   nor U39541 ( n38391,n38392,n38393 );
   nand U39542 ( n38393,n38394,n38395 );
   nand U39543 ( n38395,n37243,n38383 );
   nand U39544 ( n38394,p2_instqueue_reg_2__6_,n38384 );
   nor U39545 ( n38392,n37244,n38385 );
   nor U39546 ( n38390,n38396,n38397 );
   nor U39547 ( n38397,n37248,n38388 );
   nor U39548 ( n38396,n37247,n38389 );
   nor U39549 ( n38399,n38400,n38401 );
   nand U39550 ( n38401,n38402,n38403 );
   nand U39551 ( n38403,n37255,n38383 );
   nand U39552 ( n38402,p2_instqueue_reg_2__5_,n38384 );
   nor U39553 ( n38400,n37256,n38385 );
   nor U39554 ( n38398,n38404,n38405 );
   nor U39555 ( n38405,n37260,n38388 );
   nor U39556 ( n38404,n37259,n38389 );
   nor U39557 ( n38407,n38408,n38409 );
   nand U39558 ( n38409,n38410,n38411 );
   nand U39559 ( n38411,n37267,n38383 );
   nand U39560 ( n38410,p2_instqueue_reg_2__4_,n38384 );
   nor U39561 ( n38408,n37268,n38385 );
   nor U39562 ( n38406,n38412,n38413 );
   nor U39563 ( n38413,n37272,n38388 );
   nor U39564 ( n38412,n37271,n38389 );
   nor U39565 ( n38415,n38416,n38417 );
   nand U39566 ( n38417,n38418,n38419 );
   nand U39567 ( n38419,n37279,n38383 );
   nand U39568 ( n38418,p2_instqueue_reg_2__3_,n38384 );
   nor U39569 ( n38416,n37280,n38385 );
   nor U39570 ( n38414,n38420,n38421 );
   nor U39571 ( n38421,n37284,n38388 );
   nor U39572 ( n38420,n37283,n38389 );
   nor U39573 ( n38423,n38424,n38425 );
   nand U39574 ( n38425,n38426,n38427 );
   nand U39575 ( n38427,n37291,n38383 );
   nand U39576 ( n38426,p2_instqueue_reg_2__2_,n38384 );
   nor U39577 ( n38424,n37292,n38385 );
   nor U39578 ( n38422,n38428,n38429 );
   nor U39579 ( n38429,n37296,n38388 );
   nor U39580 ( n38428,n37295,n38389 );
   nor U39581 ( n38431,n38432,n38433 );
   nand U39582 ( n38433,n38434,n38435 );
   nand U39583 ( n38435,n37303,n38383 );
   nand U39584 ( n38434,p2_instqueue_reg_2__1_,n38384 );
   nor U39585 ( n38432,n37304,n38385 );
   nor U39586 ( n38430,n38436,n38437 );
   nor U39587 ( n38437,n37308,n38388 );
   nor U39588 ( n38436,n37307,n38389 );
   nor U39589 ( n38439,n38440,n38441 );
   nand U39590 ( n38441,n38442,n38443 );
   nand U39591 ( n38443,n37315,n38383 );
   nand U39592 ( n38383,n38444,n38445 );
   nand U39593 ( n38445,n38104,n37777 );
   nand U39594 ( n38444,p2_state2_reg_2_,n38446 );
   nand U39595 ( n38442,p2_instqueue_reg_2__0_,n38384 );
   nand U39596 ( n38384,n38447,n38448 );
   nand U39597 ( n38448,p2_state2_reg_3_,n38388 );
   nor U39598 ( n38447,n38449,n38450 );
   nor U39599 ( n38450,n38451,n37326 );
   and U39600 ( n38451,n37327,n38446 );
   nand U39601 ( n38446,n38452,n38388 );
   nor U39602 ( n38449,n38453,n38454 );
   nand U39603 ( n38454,n38455,n37331 );
   nand U39604 ( n38455,n38115,n37777 );
   nor U39605 ( n37777,n38456,n38117 );
   nor U39606 ( n38453,n38457,n36712 );
   and U39607 ( n38457,n38385,n38389 );
   nor U39608 ( n38440,n37337,n38385 );
   nand U39609 ( n38385,n38371,n37430 );
   nor U39610 ( n38438,n38458,n38459 );
   nor U39611 ( n38459,n37344,n38388 );
   nand U39612 ( n38388,n38376,n37433 );
   nor U39613 ( n38458,n37342,n38389 );
   nand U39614 ( n38389,n38374,n36687 );
   nor U39615 ( n36687,n36674,n38375 );
   nor U39616 ( n38461,n38462,n38463 );
   nand U39617 ( n38463,n38464,n38465 );
   nand U39618 ( n38465,n37226,n38466 );
   nand U39619 ( n38464,p2_instqueue_reg_1__7_,n38467 );
   nor U39620 ( n38462,n37229,n38468 );
   nor U39621 ( n38460,n38469,n38470 );
   nor U39622 ( n38470,n37233,n38471 );
   not U39623 ( n37233,n38472 );
   nor U39624 ( n38469,n37236,n38473 );
   nor U39625 ( n38475,n38476,n38477 );
   nand U39626 ( n38477,n38478,n38479 );
   nand U39627 ( n38479,n37243,n38466 );
   nand U39628 ( n38478,p2_instqueue_reg_1__6_,n38467 );
   nor U39629 ( n38476,n37244,n38468 );
   nor U39630 ( n38474,n38480,n38481 );
   nor U39631 ( n38481,n37247,n38471 );
   not U39632 ( n37247,n38482 );
   nor U39633 ( n38480,n37248,n38473 );
   nor U39634 ( n38484,n38485,n38486 );
   nand U39635 ( n38486,n38487,n38488 );
   nand U39636 ( n38488,n37255,n38466 );
   nand U39637 ( n38487,p2_instqueue_reg_1__5_,n38467 );
   nor U39638 ( n38485,n37256,n38468 );
   nor U39639 ( n38483,n38489,n38490 );
   nor U39640 ( n38490,n37259,n38471 );
   not U39641 ( n37259,n38491 );
   nor U39642 ( n38489,n37260,n38473 );
   nor U39643 ( n38493,n38494,n38495 );
   nand U39644 ( n38495,n38496,n38497 );
   nand U39645 ( n38497,n37267,n38466 );
   nand U39646 ( n38496,p2_instqueue_reg_1__4_,n38467 );
   nor U39647 ( n38494,n37268,n38468 );
   nor U39648 ( n38492,n38498,n38499 );
   nor U39649 ( n38499,n37271,n38471 );
   not U39650 ( n37271,n38500 );
   nor U39651 ( n38498,n37272,n38473 );
   nor U39652 ( n38502,n38503,n38504 );
   nand U39653 ( n38504,n38505,n38506 );
   nand U39654 ( n38506,n37279,n38466 );
   nand U39655 ( n38505,p2_instqueue_reg_1__3_,n38467 );
   nor U39656 ( n38503,n37280,n38468 );
   nor U39657 ( n38501,n38507,n38508 );
   nor U39658 ( n38508,n37283,n38471 );
   not U39659 ( n37283,n38509 );
   nor U39660 ( n38507,n37284,n38473 );
   nor U39661 ( n38511,n38512,n38513 );
   nand U39662 ( n38513,n38514,n38515 );
   nand U39663 ( n38515,n37291,n38466 );
   nand U39664 ( n38514,p2_instqueue_reg_1__2_,n38467 );
   nor U39665 ( n38512,n37292,n38468 );
   nor U39666 ( n38510,n38516,n38517 );
   nor U39667 ( n38517,n37295,n38471 );
   not U39668 ( n37295,n38518 );
   nor U39669 ( n38516,n37296,n38473 );
   nor U39670 ( n38520,n38521,n38522 );
   nand U39671 ( n38522,n38523,n38524 );
   nand U39672 ( n38524,n37303,n38466 );
   nand U39673 ( n38523,p2_instqueue_reg_1__1_,n38467 );
   nor U39674 ( n38521,n37304,n38468 );
   nor U39675 ( n38519,n38525,n38526 );
   nor U39676 ( n38526,n37307,n38471 );
   not U39677 ( n37307,n38527 );
   nor U39678 ( n38525,n37308,n38473 );
   nor U39679 ( n38529,n38530,n38531 );
   nand U39680 ( n38531,n38532,n38533 );
   nand U39681 ( n38533,n37315,n38466 );
   nand U39682 ( n38466,n38534,n38535 );
   nand U39683 ( n38535,p2_state2_reg_2_,n38536 );
   nand U39684 ( n38534,n38537,n37319 );
   nand U39685 ( n38532,p2_instqueue_reg_1__0_,n38467 );
   nand U39686 ( n38467,n38538,n38539 );
   nand U39687 ( n38539,p2_state2_reg_3_,n38473 );
   nor U39688 ( n38538,n38540,n38541 );
   nor U39689 ( n38541,n38542,n28303 );
   and U39690 ( n38542,n37327,n38536 );
   nand U39691 ( n38536,n38543,n38473 );
   nor U39692 ( n38540,n38537,n38544 );
   nand U39693 ( n38544,n38545,n37331 );
   nand U39694 ( n38545,n37332,n38546 );
   nand U39695 ( n38546,n38468,n38471 );
   nand U39696 ( n38537,n38473,n38547 );
   nand U39697 ( n38547,n38032,n37944 );
   nor U39698 ( n38032,n37427,p2_instqueuewr_addr_reg_0_ );
   nor U39699 ( n38530,n37337,n38468 );
   nand U39700 ( n38468,n38371,n37517 );
   nor U39701 ( n38528,n38548,n38549 );
   nor U39702 ( n38549,n37342,n38471 );
   nand U39703 ( n38471,n38374,n36688 );
   nor U39704 ( n36688,n38550,n36729 );
   not U39705 ( n37342,n38551 );
   nor U39706 ( n38548,n37344,n38473 );
   nand U39707 ( n38473,n38376,n37520 );
   nor U39708 ( n38553,n38554,n38555 );
   nand U39709 ( n38555,n38556,n38557 );
   nand U39710 ( n38557,n38558,n38472 );
   nand U39711 ( n38472,n38559,n38560 );
   nand U39712 ( n38560,n38561,buf2_reg_31_ );
   nand U39713 ( n38559,n38562,buf1_reg_31_ );
   or U39714 ( n38556,n28193,n38563 );
   nand U39715 ( n37236,n38564,n38565 );
   nor U39716 ( n38554,n28197,n38566 );
   and U39717 ( n37229,n38567,n38568 );
   nand U39718 ( n38568,n38561,buf2_reg_23_ );
   nand U39719 ( n38567,n38562,buf1_reg_23_ );
   nor U39720 ( n38552,n38569,n38570 );
   nor U39721 ( n38570,n38571,n38572 );
   nor U39722 ( n38569,n38573,n38574 );
   not U39723 ( n38574,n37226 );
   nor U39724 ( n37226,n38575,n38576 );
   nor U39725 ( n38578,n38579,n38580 );
   nand U39726 ( n38580,n38581,n38582 );
   nand U39727 ( n38582,n38558,n38482 );
   nand U39728 ( n38482,n38583,n38584 );
   nand U39729 ( n38584,n38561,buf2_reg_30_ );
   nand U39730 ( n38583,n38562,buf1_reg_30_ );
   or U39731 ( n38581,n38563,n28199 );
   nand U39732 ( n37248,n38564,n38585 );
   nor U39733 ( n38579,n28203,n38566 );
   and U39734 ( n37244,n38586,n38587 );
   nand U39735 ( n38587,n38561,buf2_reg_22_ );
   nand U39736 ( n38586,n38562,buf1_reg_22_ );
   nor U39737 ( n38577,n38588,n38589 );
   nor U39738 ( n38589,n38571,n38590 );
   nor U39739 ( n38588,n38573,n38591 );
   not U39740 ( n38591,n37243 );
   nor U39741 ( n37243,n38592,n38576 );
   nor U39742 ( n38594,n38595,n38596 );
   nand U39743 ( n38596,n38597,n38598 );
   nand U39744 ( n38598,n38558,n38491 );
   nand U39745 ( n38491,n38599,n38600 );
   nand U39746 ( n38600,n38561,buf2_reg_29_ );
   nand U39747 ( n38599,n38562,buf1_reg_29_ );
   or U39748 ( n38597,n38563,n28206 );
   nand U39749 ( n37260,n38564,n28239 );
   nor U39750 ( n38595,n28210,n38566 );
   and U39751 ( n37256,n38602,n38603 );
   nand U39752 ( n38603,n38561,buf2_reg_21_ );
   nand U39753 ( n38602,n38562,buf1_reg_21_ );
   nor U39754 ( n38593,n38604,n38605 );
   nor U39755 ( n38605,n38571,n38606 );
   nor U39756 ( n38604,n38573,n38607 );
   not U39757 ( n38607,n37255 );
   nor U39758 ( n37255,n38608,n38576 );
   nor U39759 ( n38610,n38611,n38612 );
   nand U39760 ( n38612,n38613,n38614 );
   nand U39761 ( n38614,n38558,n38500 );
   nand U39762 ( n38500,n38615,n38616 );
   nand U39763 ( n38616,n38561,buf2_reg_28_ );
   nand U39764 ( n38615,n38562,buf1_reg_28_ );
   or U39765 ( n38613,n38563,n28214 );
   nand U39766 ( n37272,n38564,n38617 );
   nor U39767 ( n38611,n28218,n38566 );
   and U39768 ( n37268,n38618,n38619 );
   nand U39769 ( n38619,n38561,buf2_reg_20_ );
   nand U39770 ( n38618,n38562,buf1_reg_20_ );
   nor U39771 ( n38609,n38620,n38621 );
   nor U39772 ( n38621,n38571,n38622 );
   nor U39773 ( n38620,n38573,n38623 );
   not U39774 ( n38623,n37267 );
   nor U39775 ( n37267,n38624,n38576 );
   nor U39776 ( n38626,n38627,n38628 );
   nand U39777 ( n38628,n38629,n38630 );
   nand U39778 ( n38630,n38558,n38509 );
   nand U39779 ( n38509,n38631,n38632 );
   nand U39780 ( n38632,n38561,buf2_reg_27_ );
   nand U39781 ( n38631,n38562,buf1_reg_27_ );
   or U39782 ( n38629,n38563,n28226 );
   nand U39783 ( n37284,n38564,n38633 );
   nor U39784 ( n38627,n28230,n38566 );
   and U39785 ( n37280,n38634,n38635 );
   nand U39786 ( n38635,n38561,buf2_reg_19_ );
   nand U39787 ( n38634,n38562,buf1_reg_19_ );
   nor U39788 ( n38625,n38636,n38637 );
   nor U39789 ( n38637,n38571,n38638 );
   nor U39790 ( n38636,n38573,n38639 );
   not U39791 ( n38639,n37279 );
   nor U39792 ( n37279,n38640,n38576 );
   nor U39793 ( n38642,n38643,n38644 );
   nand U39794 ( n38644,n38645,n38646 );
   nand U39795 ( n38646,n38558,n38518 );
   nand U39796 ( n38518,n38647,n38648 );
   nand U39797 ( n38648,n38561,buf2_reg_26_ );
   nand U39798 ( n38647,n38562,buf1_reg_26_ );
   or U39799 ( n38645,n38563,n28267 );
   nand U39800 ( n37296,n38564,n38649 );
   nor U39801 ( n38643,n28248,n38566 );
   and U39802 ( n37292,n38650,n38651 );
   nand U39803 ( n38651,n38561,buf2_reg_18_ );
   nand U39804 ( n38650,n38562,buf1_reg_18_ );
   nor U39805 ( n38641,n38652,n38653 );
   nor U39806 ( n38653,n38571,n38654 );
   nor U39807 ( n38652,n38573,n38655 );
   not U39808 ( n38655,n37291 );
   nor U39809 ( n37291,n38656,n38576 );
   nor U39810 ( n38658,n38659,n38660 );
   nand U39811 ( n38660,n38661,n38662 );
   nand U39812 ( n38662,n38558,n38527 );
   nand U39813 ( n38527,n38663,n38664 );
   nand U39814 ( n38664,n38561,buf2_reg_25_ );
   nand U39815 ( n38663,n38562,buf1_reg_25_ );
   or U39816 ( n38661,n38563,n28244 );
   nand U39817 ( n37308,n38564,n28280 );
   nor U39818 ( n38659,n28272,n38566 );
   and U39819 ( n37304,n38665,n38666 );
   nand U39820 ( n38666,n38561,buf2_reg_17_ );
   nand U39821 ( n38665,n38562,buf1_reg_17_ );
   nor U39822 ( n38657,n38667,n38668 );
   nor U39823 ( n38668,n38571,n38669 );
   nor U39824 ( n38667,n38573,n38670 );
   not U39825 ( n38670,n37303 );
   nor U39826 ( n37303,n38671,n38576 );
   nor U39827 ( n38673,n38674,n38675 );
   nand U39828 ( n38675,n38676,n38677 );
   nand U39829 ( n38677,n38558,n38551 );
   nand U39830 ( n38551,n38678,n38679 );
   nand U39831 ( n38679,n38561,buf2_reg_24_ );
   nand U39832 ( n38678,n38562,buf1_reg_24_ );
   or U39833 ( n38676,n38563,n28324 );
   nand U39834 ( n37344,n38564,n38680 );
   nor U39835 ( n38564,n38681,n38576 );
   nor U39836 ( n38674,n28328,n38566 );
   and U39837 ( n37337,n38682,n38683 );
   nand U39838 ( n38683,n38561,buf2_reg_16_ );
   nor U39839 ( n38561,n38684,n28750 );
   nand U39840 ( n38682,n38562,buf1_reg_16_ );
   nor U39841 ( n38562,n38684,n28739 );
   nor U39842 ( n38672,n38685,n38686 );
   nor U39843 ( n38686,n38573,n38687 );
   not U39844 ( n38687,n37315 );
   nor U39845 ( n37315,n38688,n38576 );
   and U39846 ( n38573,n38689,n38690 );
   nand U39847 ( n38690,n38104,n37944 );
   and U39848 ( n38104,n38115,n37319 );
   nand U39849 ( n37319,n37332,n36686 );
   nand U39850 ( n38689,p2_state2_reg_2_,n38691 );
   nand U39851 ( n38691,n38692,n38563 );
   nor U39852 ( n38685,n38571,n38693 );
   and U39853 ( n38571,n38694,n38695 );
   nand U39854 ( n38695,p2_state2_reg_3_,n38563 );
   nor U39855 ( n38694,n38696,n38697 );
   nor U39856 ( n38697,n38698,n28303 );
   nor U39857 ( n37326,n38576,p2_state2_reg_2_ );
   nor U39858 ( n38698,n38576,n38699 );
   and U39859 ( n38699,n38563,n38692 );
   nand U39860 ( n38563,n38376,n37605 );
   nor U39861 ( n37605,p2_instqueuewr_addr_reg_1_,p2_instqueuewr_addr_reg_0_ );
   nor U39862 ( n38376,p2_instqueuewr_addr_reg_3_,p2_instqueuewr_addr_reg_2_ );
   nor U39863 ( n38696,n38700,n38701 );
   nand U39864 ( n38701,n38702,n37331 );
   nand U39865 ( n37331,n37332,n38684 );
   or U39866 ( n38684,n36686,n38576 );
   nand U39867 ( n36686,p2_statebs16_reg,n36628 );
   not U39868 ( n37332,n36712 );
   nand U39869 ( n38702,n38115,n37944 );
   nor U39870 ( n37944,n38456,n38286 );
   not U39871 ( n38286,n38117 );
   nor U39872 ( n38700,n38703,n36712 );
   nor U39873 ( n36712,n38704,p2_statebs16_reg );
   nor U39874 ( n38703,n38558,n38705 );
   not U39875 ( n38705,n38566 );
   nand U39876 ( n38566,n37946,n38371 );
   nor U39877 ( n38371,n36772,n36752 );
   nor U39878 ( n37946,n36729,n36740 );
   and U39879 ( n38558,n38374,n37608 );
   nor U39880 ( n37608,n38550,n36674 );
   not U39881 ( n38550,n38375 );
   nor U39882 ( n38375,n37430,n37517 );
   nor U39883 ( n37517,n36674,n36740 );
   nor U39884 ( n37430,n36684,n36729 );
   nor U39885 ( n38374,n37343,n36701 );
   xor U39886 ( n36701,n37693,n36752 );
   nand U39887 ( n37343,n38706,n38707 );
   nand U39888 ( n38707,n36772,n37339 );
   nor U39889 ( n38706,n37692,n38708 );
   not U39890 ( n38708,n37960 );
   nand U39891 ( n37960,n38709,n36752 );
   nor U39892 ( n38709,n36772,n37339 );
   not U39893 ( n37339,n37693 );
   nor U39894 ( n37692,n36711,n36752 );
   not U39895 ( n36665,n36667 );
   nand U39896 ( n36667,n38710,n38711 );
   or U39897 ( n38711,n36788,n37219 );
   nor U39898 ( n38710,n37327,n36784 );
   nor U39899 ( n36784,n38712,n36788 );
   nand U39900 ( n36788,n38713,p2_state2_reg_1_ );
   nor U39901 ( n38713,n37217,n36783 );
   not U39902 ( n37327,n38576 );
   nand U39903 ( n38576,n38714,n27895 );
   nand U39904 ( n38714,n38715,n38716 );
   nand U39905 ( n38716,p2_state2_reg_1_,n37217 );
   nor U39906 ( n38715,n37035,n36728 );
   nor U39907 ( n36728,n38681,n37168 );
   nor U39908 ( n38718,n38719,n38720 );
   nand U39909 ( n38720,n38721,n38722 );
   nand U39910 ( n38722,n38723,n28346 );
   nand U39911 ( n38721,n38725,n36670 );
   nor U39912 ( n38719,n38726,n28275 );
   nor U39913 ( n38717,n38728,n38729 );
   nand U39914 ( n38729,n38730,n38731 );
   nand U39915 ( n38731,n38732,p2_reip_reg_0_ );
   or U39916 ( n38730,n38733,n38734 );
   nand U39917 ( n38728,n38735,n38736 );
   nand U39918 ( n38736,n28304,p2_instaddrpointer_reg_0_ );
   nor U39919 ( n38739,n38740,n38741 );
   nand U39920 ( n38741,n38742,n38743 );
   nand U39921 ( n38743,n38725,n36680 );
   nand U39922 ( n38742,n38744,n38745 );
   nor U39923 ( n38740,n36961,n38746 );
   nor U39924 ( n38738,n38747,n38748 );
   nand U39925 ( n38748,n38749,n38750 );
   nand U39926 ( n38750,n38751,n28343 );
   nand U39927 ( n38749,n38753,n28346 );
   nand U39928 ( n38747,n38754,n38755 );
   nand U39929 ( n38755,p2_instaddrpointer_reg_1_,n38756 );
   nand U39930 ( n38756,n38757,n38735 );
   nand U39931 ( n38735,n38758,n36762 );
   nand U39932 ( n38754,n38759,n36758 );
   and U39933 ( n38759,n38758,p2_instaddrpointer_reg_0_ );
   nor U39934 ( n38761,n38762,n38763 );
   nand U39935 ( n38763,n38764,n38765 );
   nand U39936 ( n38765,n38744,n38766 );
   nand U39937 ( n38764,n38732,p2_reip_reg_2_ );
   nand U39938 ( n38762,n38767,n38768 );
   nand U39939 ( n38768,n38769,n38770 );
   nand U39940 ( n38770,n38771,n38772 );
   nand U39941 ( n38767,n38725,n36694 );
   nor U39942 ( n38760,n38773,n38774 );
   nand U39943 ( n38774,n38775,n38776 );
   nand U39944 ( n38776,n38777,n28343 );
   nand U39945 ( n38775,n38724,n38778 );
   nand U39946 ( n38773,n38779,n38780 );
   nand U39947 ( n38780,p2_instaddrpointer_reg_2_,n38781 );
   nand U39948 ( n38781,n38757,n38782 );
   nand U39949 ( n38782,n38783,n38784 );
   nand U39950 ( n38779,n38785,n38786 );
   nor U39951 ( n38785,n38784,n38787 );
   nor U39952 ( n38789,n38790,n38791 );
   nand U39953 ( n38791,n38792,n38793 );
   nand U39954 ( n38793,n38752,n38794 );
   nand U39955 ( n38792,n38725,n36708 );
   not U39956 ( n36708,n38795 );
   nor U39957 ( n38790,n37159,n28275 );
   nor U39958 ( n38788,n38796,n38797 );
   nand U39959 ( n38797,n38798,n38799 );
   nand U39960 ( n38799,n28269,p2_reip_reg_3_ );
   nand U39961 ( n38798,n38724,n38800 );
   nand U39962 ( n38796,n38801,n38802 );
   nand U39963 ( n38802,p2_instaddrpointer_reg_3_,n38803 );
   nand U39964 ( n38801,n38804,n38805 );
   nor U39965 ( n38807,n38808,n38809 );
   nand U39966 ( n38809,n38810,n38811 );
   nand U39967 ( n38811,n38812,n28326 );
   nand U39968 ( n38810,n38813,n38744 );
   nor U39969 ( n38808,n36945,n38746 );
   nor U39970 ( n38806,n38814,n38815 );
   nand U39971 ( n38815,n38816,n38817 );
   nand U39972 ( n38817,n38752,n38818 );
   nand U39973 ( n38816,n28346,n38819 );
   nand U39974 ( n38814,n38820,n38821 );
   nand U39975 ( n38821,p2_instaddrpointer_reg_4_,n38822 );
   nand U39976 ( n38822,n38823,n38824 );
   nand U39977 ( n38824,n28301,n38805 );
   not U39978 ( n38823,n38803 );
   nand U39979 ( n38803,n38825,n38826 );
   nand U39980 ( n38826,n38783,n38771 );
   nor U39981 ( n38825,n28304,n38827 );
   nor U39982 ( n38827,n38828,n38772 );
   nand U39983 ( n38820,n38829,n38830 );
   and U39984 ( n38829,n38804,p2_instaddrpointer_reg_3_ );
   nand U39985 ( n38804,n38831,n38832 );
   nand U39986 ( n38832,n38769,n38772 );
   or U39987 ( n38831,n38771,n38787 );
   nor U39988 ( n38834,n38835,n38836 );
   nand U39989 ( n38836,n38837,n38838 );
   nand U39990 ( n38838,n38839,n28326 );
   nand U39991 ( n38837,n38840,n38744 );
   nor U39992 ( n38835,n36940,n38746 );
   nor U39993 ( n38833,n38841,n38842 );
   nand U39994 ( n38842,n38843,n38844 );
   nand U39995 ( n38844,n38752,n38845 );
   nand U39996 ( n38843,n38724,n38846 );
   nand U39997 ( n38841,n38847,n38848 );
   nand U39998 ( n38848,p2_instaddrpointer_reg_5_,n38849 );
   nand U39999 ( n38847,n38850,n38851 );
   nor U40000 ( n38853,n38854,n38855 );
   nand U40001 ( n38855,n38856,n38857 );
   nand U40002 ( n38857,n38858,n38725 );
   nand U40003 ( n38856,n38859,n38744 );
   nor U40004 ( n38854,n36935,n38746 );
   nor U40005 ( n38852,n38860,n38861 );
   nand U40006 ( n38861,n38862,n38863 );
   nand U40007 ( n38863,n38752,n38864 );
   nand U40008 ( n38862,n38724,n38865 );
   nand U40009 ( n38860,n38866,n38867 );
   nand U40010 ( n38867,p2_instaddrpointer_reg_6_,n38868 );
   nand U40011 ( n38868,n38869,n38870 );
   nand U40012 ( n38870,n38758,n38851 );
   not U40013 ( n38869,n38849 );
   nand U40014 ( n38849,n38871,n38872 );
   nand U40015 ( n38872,n38783,n38873 );
   nor U40016 ( n38871,n28304,n38874 );
   nor U40017 ( n38874,n38875,n38828 );
   nand U40018 ( n38866,n38876,n38877 );
   and U40019 ( n38876,n38850,p2_instaddrpointer_reg_5_ );
   nand U40020 ( n38850,n38878,n38879 );
   nand U40021 ( n38879,n38875,n38769 );
   not U40022 ( n38875,n38880 );
   or U40023 ( n38878,n38873,n38787 );
   nor U40024 ( n38882,n38883,n38884 );
   nand U40025 ( n38884,n38885,n38886 );
   nand U40026 ( n38886,n38887,n28326 );
   nand U40027 ( n38885,n38888,n38744 );
   nor U40028 ( n38883,n36930,n38746 );
   nor U40029 ( n38881,n38889,n38890 );
   nand U40030 ( n38890,n38891,n38892 );
   nand U40031 ( n38892,n28343,n38893 );
   nand U40032 ( n38891,n38724,n38894 );
   nand U40033 ( n38889,n38895,n38896 );
   nand U40034 ( n38896,p2_instaddrpointer_reg_7_,n38897 );
   nand U40035 ( n38895,n38898,n38899 );
   nor U40036 ( n38901,n38902,n38903 );
   nand U40037 ( n38903,n38904,n38905 );
   nand U40038 ( n38905,n38724,n38906 );
   nand U40039 ( n38904,n38907,n38725 );
   nor U40040 ( n38902,n28275,n38908 );
   nor U40041 ( n38900,n38909,n38910 );
   nand U40042 ( n38910,n38911,n38912 );
   nand U40043 ( n38912,n38732,p2_reip_reg_8_ );
   nand U40044 ( n38911,n38752,n38913 );
   nand U40045 ( n38909,n38914,n38915 );
   nand U40046 ( n38915,p2_instaddrpointer_reg_8_,n38916 );
   nand U40047 ( n38916,n38917,n38918 );
   nand U40048 ( n38918,n38758,n38899 );
   not U40049 ( n38917,n38897 );
   nand U40050 ( n38897,n38919,n38920 );
   nand U40051 ( n38920,n38783,n38921 );
   nor U40052 ( n38919,n38737,n38922 );
   nor U40053 ( n38922,n38923,n38828 );
   nand U40054 ( n38914,n38924,n38925 );
   and U40055 ( n38924,n38898,p2_instaddrpointer_reg_7_ );
   nand U40056 ( n38898,n38926,n38927 );
   nand U40057 ( n38927,n38923,n38769 );
   not U40058 ( n38923,n38928 );
   or U40059 ( n38926,n38921,n38787 );
   nor U40060 ( n38930,n38931,n38932 );
   nand U40061 ( n38932,n38933,n38934 );
   nand U40062 ( n38934,n38752,n38935 );
   nand U40063 ( n38933,n38936,n28346 );
   nor U40064 ( n38931,n38937,n38938 );
   nor U40065 ( n38929,n38939,n38940 );
   nand U40066 ( n38940,n38941,n38942 );
   nand U40067 ( n38942,n38943,n38744 );
   nand U40068 ( n38941,n28269,p2_reip_reg_9_ );
   nand U40069 ( n38939,n38944,n38945 );
   nand U40070 ( n38945,p2_instaddrpointer_reg_9_,n38946 );
   nand U40071 ( n38944,n38947,n38948 );
   nor U40072 ( n38950,n38951,n38952 );
   nand U40073 ( n38952,n38953,n38954 );
   nand U40074 ( n38954,n38955,n28346 );
   nand U40075 ( n38953,n38956,n28343 );
   nor U40076 ( n38951,n38937,n38957 );
   nor U40077 ( n38949,n38958,n38959 );
   nand U40078 ( n38959,n38960,n38961 );
   nand U40079 ( n38961,n38962,n38744 );
   nand U40080 ( n38960,n28269,p2_reip_reg_10_ );
   nand U40081 ( n38958,n38963,n38964 );
   nand U40082 ( n38964,p2_instaddrpointer_reg_10_,n38965 );
   nand U40083 ( n38965,n38966,n38967 );
   nand U40084 ( n38967,n28301,n38948 );
   not U40085 ( n38966,n38946 );
   nand U40086 ( n38946,n38968,n38969 );
   nand U40087 ( n38969,n38783,n38970 );
   nor U40088 ( n38968,n38737,n38971 );
   nor U40089 ( n38971,n38972,n38828 );
   nand U40090 ( n38963,n38973,n38974 );
   and U40091 ( n38973,n38947,p2_instaddrpointer_reg_9_ );
   nand U40092 ( n38947,n38975,n38976 );
   nand U40093 ( n38976,n38972,n38769 );
   not U40094 ( n38972,n38977 );
   or U40095 ( n38975,n38970,n38787 );
   nor U40096 ( n38979,n38980,n38981 );
   nand U40097 ( n38981,n38982,n38983 );
   nand U40098 ( n38983,n28343,n38984 );
   nand U40099 ( n38982,n38724,n38985 );
   nor U40100 ( n38980,n38937,n38986 );
   nor U40101 ( n38978,n38987,n38988 );
   nand U40102 ( n38988,n38989,n38990 );
   nand U40103 ( n38990,n38991,n38744 );
   nand U40104 ( n38989,n28269,p2_reip_reg_11_ );
   nand U40105 ( n38987,n38992,n38993 );
   nand U40106 ( n38993,p2_instaddrpointer_reg_11_,n38994 );
   nand U40107 ( n38992,n38995,n38996 );
   nor U40108 ( n38998,n38999,n39000 );
   nand U40109 ( n39000,n39001,n39002 );
   nand U40110 ( n39002,n39003,n38725 );
   nand U40111 ( n39001,n39004,n38744 );
   nor U40112 ( n38999,n36905,n38746 );
   nor U40113 ( n38997,n39005,n39006 );
   nand U40114 ( n39006,n39007,n39008 );
   nand U40115 ( n39008,n38752,n39009 );
   nand U40116 ( n39007,n38724,n39010 );
   nand U40117 ( n39005,n39011,n39012 );
   nand U40118 ( n39012,p2_instaddrpointer_reg_12_,n39013 );
   nand U40119 ( n39013,n39014,n39015 );
   nand U40120 ( n39015,n38758,n38996 );
   not U40121 ( n39014,n38994 );
   nand U40122 ( n38994,n39016,n39017 );
   nand U40123 ( n39017,n38783,n39018 );
   nor U40124 ( n39016,n38737,n39019 );
   nor U40125 ( n39019,n39020,n38828 );
   nand U40126 ( n39011,n39021,n39022 );
   and U40127 ( n39021,n38995,p2_instaddrpointer_reg_11_ );
   nand U40128 ( n38995,n39023,n39024 );
   nand U40129 ( n39024,n39020,n38769 );
   nand U40130 ( n39023,n39025,n38783 );
   nor U40131 ( n39027,n39028,n39029 );
   nand U40132 ( n39029,n39030,n39031 );
   nand U40133 ( n39031,n39032,n28346 );
   nand U40134 ( n39030,n39033,n38725 );
   nor U40135 ( n39028,n38727,n39034 );
   nor U40136 ( n39026,n39035,n39036 );
   nand U40137 ( n39036,n39037,n39038 );
   nand U40138 ( n39038,n38732,p2_reip_reg_13_ );
   nand U40139 ( n39037,n28343,n39039 );
   nand U40140 ( n39035,n39040,n39041 );
   nand U40141 ( n39041,n39042,n39043 );
   nand U40142 ( n39040,p2_instaddrpointer_reg_13_,n39044 );
   nor U40143 ( n39046,n39047,n39048 );
   nand U40144 ( n39048,n39049,n39050 );
   nand U40145 ( n39050,n38724,n39051 );
   nand U40146 ( n39049,n39052,n38725 );
   nor U40147 ( n39047,n38727,n39053 );
   nor U40148 ( n39045,n39054,n39055 );
   nand U40149 ( n39055,n39056,n39057 );
   nand U40150 ( n39057,n38732,p2_reip_reg_14_ );
   nand U40151 ( n39056,n38752,n39058 );
   nand U40152 ( n39054,n39059,n39060 );
   nand U40153 ( n39060,p2_instaddrpointer_reg_14_,n39061 );
   nand U40154 ( n39061,n39062,n39063 );
   nand U40155 ( n39063,n38758,n39043 );
   not U40156 ( n39062,n39044 );
   nand U40157 ( n39044,n39064,n39065 );
   nand U40158 ( n39065,n38783,n39066 );
   nor U40159 ( n39064,n38737,n39067 );
   nor U40160 ( n39067,n39068,n38828 );
   nand U40161 ( n39059,n39069,n39070 );
   and U40162 ( n39069,n39042,p2_instaddrpointer_reg_13_ );
   nand U40163 ( n39042,n39071,n39072 );
   nand U40164 ( n39072,n39068,n38769 );
   nand U40165 ( n39071,n39073,n38783 );
   nor U40166 ( n39075,n39076,n39077 );
   nand U40167 ( n39077,n39078,n39079 );
   nand U40168 ( n39079,n39080,n38725 );
   nand U40169 ( n39078,n39081,n38744 );
   nor U40170 ( n39076,n36890,n38746 );
   nor U40171 ( n39074,n39082,n39083 );
   nand U40172 ( n39083,n39084,n39085 );
   nand U40173 ( n39085,n38752,n39086 );
   nand U40174 ( n39084,n38724,n39087 );
   nand U40175 ( n39082,n39088,n39089 );
   nand U40176 ( n39089,p2_instaddrpointer_reg_15_,n39090 );
   nand U40177 ( n39088,n39091,n39092 );
   nor U40178 ( n39094,n39095,n39096 );
   nand U40179 ( n39096,n39097,n39098 );
   nand U40180 ( n39098,n39099,n28346 );
   nand U40181 ( n39097,n39100,n38725 );
   nor U40182 ( n39095,n28275,n39101 );
   nor U40183 ( n39093,n39102,n39103 );
   nand U40184 ( n39103,n39104,n39105 );
   nand U40185 ( n39105,n38732,p2_reip_reg_16_ );
   nand U40186 ( n39104,n38752,n39106 );
   nand U40187 ( n39102,n39107,n39108 );
   nand U40188 ( n39108,p2_instaddrpointer_reg_16_,n39109 );
   nand U40189 ( n39109,n39110,n39111 );
   nand U40190 ( n39111,n38758,n39092 );
   not U40191 ( n39110,n39090 );
   nand U40192 ( n39090,n39112,n39113 );
   nand U40193 ( n39113,n38783,n39114 );
   nor U40194 ( n39112,n38737,n39115 );
   nor U40195 ( n39115,n39116,n38828 );
   nand U40196 ( n39107,n39117,n39118 );
   and U40197 ( n39117,n39091,p2_instaddrpointer_reg_15_ );
   nand U40198 ( n39091,n39119,n39120 );
   nand U40199 ( n39120,n39116,n38769 );
   not U40200 ( n39116,n39121 );
   or U40201 ( n39119,n39114,n38787 );
   nor U40202 ( n39123,n39124,n39125 );
   nand U40203 ( n39125,n39126,n39127 );
   nand U40204 ( n39127,n28346,n39128 );
   nand U40205 ( n39126,n39129,n38725 );
   nor U40206 ( n39124,n28275,n39130 );
   nor U40207 ( n39122,n39131,n39132 );
   nand U40208 ( n39132,n39133,n39134 );
   nand U40209 ( n39134,n38732,p2_reip_reg_17_ );
   nand U40210 ( n39133,n38752,n39135 );
   nand U40211 ( n39131,n39136,n39137 );
   nand U40212 ( n39137,p2_instaddrpointer_reg_17_,n39138 );
   nand U40213 ( n39136,n39139,n39140 );
   nor U40214 ( n39142,n39143,n39144 );
   nand U40215 ( n39144,n39145,n39146 );
   nand U40216 ( n39146,n39147,n28343 );
   nand U40217 ( n39145,n39148,n38725 );
   nor U40218 ( n39143,n28275,n39149 );
   nor U40219 ( n39141,n39150,n39151 );
   nand U40220 ( n39151,n39152,n39153 );
   nand U40221 ( n39153,n38732,p2_reip_reg_18_ );
   nand U40222 ( n39152,n28346,n39154 );
   nand U40223 ( n39150,n39155,n39156 );
   nand U40224 ( n39156,p2_instaddrpointer_reg_18_,n39157 );
   nand U40225 ( n39157,n39158,n39159 );
   nand U40226 ( n39159,n38758,n39140 );
   not U40227 ( n39158,n39138 );
   nand U40228 ( n39138,n39160,n39161 );
   nand U40229 ( n39161,n38783,n39162 );
   nor U40230 ( n39160,n38737,n39163 );
   nor U40231 ( n39163,n39164,n28236 );
   nand U40232 ( n39155,n39165,n39166 );
   and U40233 ( n39165,n39139,p2_instaddrpointer_reg_17_ );
   nand U40234 ( n39139,n39167,n39168 );
   nand U40235 ( n39168,n39164,n38769 );
   not U40236 ( n39164,n39169 );
   or U40237 ( n39167,n39162,n38787 );
   nor U40238 ( n39171,n39172,n39173 );
   nand U40239 ( n39173,n39174,n39175 );
   nand U40240 ( n39175,n39176,n28343 );
   nand U40241 ( n39174,n39177,n38725 );
   nor U40242 ( n39172,n28275,n39178 );
   nor U40243 ( n39170,n39179,n39180 );
   nand U40244 ( n39180,n39181,n39182 );
   nand U40245 ( n39182,n38732,p2_reip_reg_19_ );
   nand U40246 ( n39181,n39183,n28346 );
   nand U40247 ( n39179,n39184,n39185 );
   nand U40248 ( n39185,p2_instaddrpointer_reg_19_,n39186 );
   nand U40249 ( n39184,n39187,n39188 );
   nor U40250 ( n39190,n39191,n39192 );
   nand U40251 ( n39192,n39193,n39194 );
   nand U40252 ( n39194,n39195,n28346 );
   nand U40253 ( n39193,n39196,n38725 );
   nor U40254 ( n39191,n38727,n39197 );
   nor U40255 ( n39189,n39198,n39199 );
   nand U40256 ( n39199,n39200,n39201 );
   nand U40257 ( n39201,n38732,p2_reip_reg_20_ );
   nand U40258 ( n39200,n39202,n28343 );
   nand U40259 ( n39198,n39203,n39204 );
   nand U40260 ( n39204,p2_instaddrpointer_reg_20_,n39205 );
   nand U40261 ( n39205,n39206,n39207 );
   nand U40262 ( n39207,n38758,n39188 );
   not U40263 ( n39206,n39186 );
   nand U40264 ( n39186,n39208,n39209 );
   nand U40265 ( n39209,n38783,n39210 );
   nand U40266 ( n39203,n39211,n39212 );
   and U40267 ( n39211,n39187,p2_instaddrpointer_reg_19_ );
   nand U40268 ( n39187,n39213,n39214 );
   or U40269 ( n39214,n39215,n28236 );
   or U40270 ( n39213,n39210,n38787 );
   nor U40271 ( n39217,n39218,n39219 );
   nand U40272 ( n39219,n39220,n39221 );
   nand U40273 ( n39221,n38724,n39222 );
   nand U40274 ( n39220,n39223,n38725 );
   nor U40275 ( n39218,n38727,n39224 );
   nor U40276 ( n39216,n39225,n39226 );
   nand U40277 ( n39226,n39227,n39228 );
   nand U40278 ( n39228,n38732,p2_reip_reg_21_ );
   nand U40279 ( n39227,n39229,n28343 );
   nand U40280 ( n39225,n39230,n39231 );
   nand U40281 ( n39231,p2_instaddrpointer_reg_21_,n39232 );
   nand U40282 ( n39230,n39233,n39234 );
   nor U40283 ( n39236,n39237,n39238 );
   nand U40284 ( n39238,n39239,n39240 );
   nand U40285 ( n39240,n39241,n38725 );
   nand U40286 ( n39239,n39242,n38744 );
   nor U40287 ( n39237,n36855,n38746 );
   nor U40288 ( n39235,n39243,n39244 );
   nand U40289 ( n39244,n39245,n39246 );
   nand U40290 ( n39246,n38752,n39247 );
   nand U40291 ( n39245,n39248,n28346 );
   nand U40292 ( n39243,n39249,n39250 );
   nand U40293 ( n39250,p2_instaddrpointer_reg_22_,n39251 );
   nand U40294 ( n39251,n39252,n39253 );
   nand U40295 ( n39253,n38758,n39234 );
   not U40296 ( n39252,n39232 );
   nand U40297 ( n39232,n39254,n39208 );
   and U40298 ( n39208,n38757,n39255 );
   nand U40299 ( n39255,n38769,n39215 );
   nor U40300 ( n39254,n39256,n39257 );
   nor U40301 ( n39257,n39258,n38787 );
   nor U40302 ( n39256,n39259,n38828 );
   nand U40303 ( n39249,n39260,n39261 );
   and U40304 ( n39260,n39233,p2_instaddrpointer_reg_21_ );
   nand U40305 ( n39233,n39262,n39263 );
   nand U40306 ( n39263,n39264,n39259 );
   nor U40307 ( n39264,n38828,n39215 );
   nand U40308 ( n39262,n39258,n38783 );
   nor U40309 ( n39266,n39267,n39268 );
   nand U40310 ( n39268,n39269,n39270 );
   nand U40311 ( n39270,n39271,n28346 );
   nand U40312 ( n39269,n39272,n38725 );
   nor U40313 ( n39267,n38727,n39273 );
   nor U40314 ( n39265,n39274,n39275 );
   nand U40315 ( n39275,n39276,n39277 );
   nand U40316 ( n39277,n28269,p2_reip_reg_23_ );
   nand U40317 ( n39276,n39278,n28343 );
   nand U40318 ( n39274,n39279,n39280 );
   nand U40319 ( n39280,p2_instaddrpointer_reg_23_,n39281 );
   nand U40320 ( n39279,n39282,n39283 );
   nor U40321 ( n39285,n39286,n39287 );
   nand U40322 ( n39287,n39288,n39289 );
   nand U40323 ( n39289,n38724,n39290 );
   nand U40324 ( n39288,n39291,n38725 );
   nor U40325 ( n39286,n38727,n39292 );
   nor U40326 ( n39284,n39293,n39294 );
   nand U40327 ( n39294,n39295,n39296 );
   nand U40328 ( n39296,n38732,p2_reip_reg_24_ );
   nand U40329 ( n39295,n38752,n39297 );
   nand U40330 ( n39293,n39298,n39299 );
   nand U40331 ( n39299,p2_instaddrpointer_reg_24_,n39300 );
   nand U40332 ( n39300,n39301,n39302 );
   nand U40333 ( n39302,n38758,n39283 );
   not U40334 ( n39301,n39281 );
   nand U40335 ( n39281,n39303,n39304 );
   nand U40336 ( n39304,n38783,n39305 );
   nor U40337 ( n39303,n38737,n39306 );
   nor U40338 ( n39306,n39307,n38828 );
   nand U40339 ( n39298,n39308,n39309 );
   and U40340 ( n39308,n39282,p2_instaddrpointer_reg_23_ );
   nand U40341 ( n39282,n39310,n39311 );
   nand U40342 ( n39311,n39307,n38769 );
   not U40343 ( n39307,n39312 );
   or U40344 ( n39310,n39305,n38787 );
   nor U40345 ( n39314,n39315,n39316 );
   nand U40346 ( n39316,n39317,n39318 );
   nand U40347 ( n39318,n39319,n28326 );
   nand U40348 ( n39317,n39320,n38744 );
   nor U40349 ( n39315,n36840,n38746 );
   nor U40350 ( n39313,n39321,n39322 );
   nand U40351 ( n39322,n39323,n39324 );
   nand U40352 ( n39324,n39325,n28343 );
   nand U40353 ( n39323,n38724,n39326 );
   nand U40354 ( n39321,n39327,n39328 );
   nand U40355 ( n39328,p2_instaddrpointer_reg_25_,n39329 );
   nand U40356 ( n39327,n39330,n39331 );
   nor U40357 ( n39333,n39334,n39335 );
   nand U40358 ( n39335,n39336,n39337 );
   nand U40359 ( n39337,n38752,n39338 );
   nand U40360 ( n39336,n39339,n38725 );
   nor U40361 ( n39334,n38727,n39340 );
   nor U40362 ( n39332,n39341,n39342 );
   nand U40363 ( n39342,n39343,n39344 );
   nand U40364 ( n39344,n38732,p2_reip_reg_26_ );
   nand U40365 ( n39343,n38724,n39345 );
   nand U40366 ( n39341,n39346,n39347 );
   nand U40367 ( n39347,p2_instaddrpointer_reg_26_,n39348 );
   nand U40368 ( n39348,n39349,n39350 );
   nand U40369 ( n39350,n38758,n39331 );
   not U40370 ( n39349,n39329 );
   nand U40371 ( n39329,n39351,n39352 );
   nand U40372 ( n39352,n38783,n39353 );
   nor U40373 ( n39351,n38737,n39354 );
   nor U40374 ( n39354,n39355,n38828 );
   nand U40375 ( n39346,n39356,n39357 );
   and U40376 ( n39356,n39330,p2_instaddrpointer_reg_25_ );
   nand U40377 ( n39330,n39358,n39359 );
   nand U40378 ( n39359,n39355,n38769 );
   not U40379 ( n39355,n39360 );
   or U40380 ( n39358,n39353,n38787 );
   nor U40381 ( n39362,n39363,n39364 );
   nand U40382 ( n39364,n39365,n39366 );
   nand U40383 ( n39366,n38724,n39367 );
   nand U40384 ( n39365,n39368,n38725 );
   nor U40385 ( n39363,n38727,n39369 );
   nor U40386 ( n39361,n39370,n39371 );
   nand U40387 ( n39371,n39372,n39373 );
   nand U40388 ( n39373,n38732,p2_reip_reg_27_ );
   nand U40389 ( n39372,n39374,n28343 );
   nand U40390 ( n39370,n39375,n39376 );
   nand U40391 ( n39376,p2_instaddrpointer_reg_27_,n39377 );
   nand U40392 ( n39375,n39378,n39379 );
   nor U40393 ( n39381,n39382,n39383 );
   nand U40394 ( n39383,n39384,n39385 );
   nand U40395 ( n39385,n39386,n38725 );
   nand U40396 ( n39384,n39387,n38744 );
   nor U40397 ( n39382,n36825,n38746 );
   not U40398 ( n38746,n38732 );
   nor U40399 ( n39380,n39388,n39389 );
   nand U40400 ( n39389,n39390,n39391 );
   nand U40401 ( n39391,n39392,n28343 );
   nand U40402 ( n39390,n39393,n28346 );
   nand U40403 ( n39388,n39394,n39395 );
   or U40404 ( n39395,n39396,n39397 );
   nand U40405 ( n39394,n39398,n39396 );
   nor U40406 ( n39400,n39401,n39402 );
   nand U40407 ( n39402,n39403,n39404 );
   nand U40408 ( n39404,n39405,n28346 );
   nand U40409 ( n39403,n39406,n28326 );
   nor U40410 ( n39401,n38727,n39407 );
   nor U40411 ( n39399,n39408,n39409 );
   nand U40412 ( n39409,n39410,n39411 );
   nand U40413 ( n39411,n38732,p2_reip_reg_29_ );
   nand U40414 ( n39410,n39412,n28343 );
   nand U40415 ( n39408,n39413,n39414 );
   nand U40416 ( n39414,n39415,n39416 );
   nand U40417 ( n39413,p2_instaddrpointer_reg_29_,n39417 );
   nor U40418 ( n39419,n39420,n39421 );
   nand U40419 ( n39421,n39422,n39423 );
   nand U40420 ( n39423,n39424,n38744 );
   nand U40421 ( n39422,n38752,n39425 );
   not U40422 ( n38752,n38733 );
   nor U40423 ( n39420,n39426,n39427 );
   nor U40424 ( n39418,n39428,n39429 );
   nand U40425 ( n39429,n39430,n39431 );
   nand U40426 ( n39431,n39432,n28326 );
   not U40427 ( n38725,n38937 );
   nand U40428 ( n39430,n38732,p2_reip_reg_30_ );
   nand U40429 ( n39428,n39433,n39434 );
   or U40430 ( n39434,n39435,n39436 );
   nand U40431 ( n39433,n39437,n39435 );
   nor U40432 ( n39437,n39416,n39438 );
   nor U40433 ( n39440,n39441,n39442 );
   nand U40434 ( n39442,n39443,n39444 );
   nand U40435 ( n39444,n39445,n39446 );
   nor U40436 ( n39445,n39447,n38733 );
   nand U40437 ( n38733,n39448,n37202 );
   nand U40438 ( n39443,n38724,n39449 );
   not U40439 ( n38724,n39427 );
   nand U40440 ( n39427,n39450,n39448 );
   nor U40441 ( n39441,n38937,n39451 );
   nand U40442 ( n38937,n39448,n39452 );
   nand U40443 ( n39452,n39453,n39454 );
   nand U40444 ( n39454,n39455,n39456 );
   nor U40445 ( n39453,n37180,n37171 );
   nor U40446 ( n39439,n39457,n39458 );
   nand U40447 ( n39458,n39459,n39460 );
   nand U40448 ( n39460,n39461,n38744 );
   not U40449 ( n38744,n38727 );
   nand U40450 ( n38727,n39448,n39462 );
   nand U40451 ( n39462,n39463,n39464 );
   nor U40452 ( n39464,n37182,n37188 );
   nor U40453 ( n37188,n39465,n39466 );
   nand U40454 ( n39465,n38585,n39467 );
   nor U40455 ( n37182,n37133,n39466 );
   nand U40456 ( n37133,n39468,n39467 );
   nor U40457 ( n39468,n37195,n38585 );
   nor U40458 ( n39463,n37068,n36776 );
   nand U40459 ( n39459,n28269,p2_reip_reg_31_ );
   nor U40460 ( n38732,n38737,p2_state2_reg_2_ );
   nand U40461 ( n39457,n39469,n39470 );
   nand U40462 ( n39470,p2_instaddrpointer_reg_31_,n39471 );
   nand U40463 ( n39471,n39436,n39472 );
   nand U40464 ( n39472,n38758,n39435 );
   nor U40465 ( n39436,n39417,n39473 );
   and U40466 ( n39473,n38758,n39416 );
   nand U40467 ( n39417,n39397,n39474 );
   nand U40468 ( n39474,n28301,n39396 );
   nor U40469 ( n39397,n39377,n39475 );
   and U40470 ( n39475,n38758,n39379 );
   nand U40471 ( n38758,n38787,n28236 );
   nand U40472 ( n39377,n39476,n39477 );
   nand U40473 ( n39477,n38783,n39478 );
   not U40474 ( n38783,n38787 );
   nor U40475 ( n39476,n38737,n39479 );
   nor U40476 ( n39479,n39480,n38828 );
   nand U40477 ( n39469,n39481,n39482 );
   nor U40478 ( n39481,n39435,n39483 );
   nand U40479 ( n39483,n39415,p2_instaddrpointer_reg_29_ );
   not U40480 ( n39415,n39438 );
   nand U40481 ( n39438,n39398,p2_instaddrpointer_reg_28_ );
   nor U40482 ( n39398,n39484,n39379 );
   not U40483 ( n39484,n39378 );
   nand U40484 ( n39378,n39485,n39486 );
   nand U40485 ( n39486,n39480,n38769 );
   not U40486 ( n38769,n38828 );
   nand U40487 ( n38828,n39448,n37179 );
   and U40488 ( n39480,n39487,p2_instaddrpointer_reg_26_ );
   nor U40489 ( n39487,n39331,n39360 );
   nand U40490 ( n39360,n39488,p2_instaddrpointer_reg_24_ );
   nor U40491 ( n39488,n39283,n39312 );
   nand U40492 ( n39312,n39489,n39490 );
   nor U40493 ( n39489,n39215,n39491 );
   nand U40494 ( n39215,n39492,p2_instaddrpointer_reg_18_ );
   nor U40495 ( n39492,n39140,n39169 );
   nand U40496 ( n39169,n39493,p2_instaddrpointer_reg_16_ );
   nor U40497 ( n39493,n39092,n39121 );
   nand U40498 ( n39121,n39494,n39068 );
   and U40499 ( n39068,n39495,p2_instaddrpointer_reg_12_ );
   and U40500 ( n39495,p2_instaddrpointer_reg_11_,n39020 );
   nor U40501 ( n39020,n39496,n38977 );
   nand U40502 ( n38977,n39497,p2_instaddrpointer_reg_8_ );
   nor U40503 ( n39497,n38899,n38928 );
   nand U40504 ( n38928,n39498,p2_instaddrpointer_reg_6_ );
   nor U40505 ( n39498,n38851,n38880 );
   nand U40506 ( n38880,n39499,p2_instaddrpointer_reg_4_ );
   and U40507 ( n39499,n38772,p2_instaddrpointer_reg_3_ );
   nand U40508 ( n38772,n38786,n38784 );
   or U40509 ( n39485,n39478,n38787 );
   nand U40510 ( n38787,n39448,n39500 );
   nand U40511 ( n39500,n37190,n39501 );
   nor U40512 ( n39501,n37183,n39502 );
   nor U40513 ( n39502,n39503,n37194 );
   nor U40514 ( n39503,n39504,n38617 );
   nor U40515 ( n39504,n39505,n39506 );
   not U40516 ( n37183,n39507 );
   nor U40517 ( n37190,n39508,n39509 );
   nand U40518 ( n39509,n39510,n39511 );
   nand U40519 ( n39511,n39512,n39513 );
   nand U40520 ( n39513,n39514,n37130 );
   nor U40521 ( n39514,n39515,n38680 );
   nand U40522 ( n39512,n37113,n39516 );
   nor U40523 ( n39510,n39517,n39518 );
   nor U40524 ( n39518,n39519,n37136 );
   nor U40525 ( n39517,n39520,n39521 );
   nand U40526 ( n39521,n38633,n28280 );
   nand U40527 ( n39508,n39522,n39523 );
   nand U40528 ( n39523,n39524,n37130 );
   nor U40529 ( n39524,n39525,n38649 );
   nor U40530 ( n39525,n39526,n39527 );
   nor U40531 ( n39526,n39528,n39529 );
   nand U40532 ( n39522,n39530,n39531 );
   nand U40533 ( n39531,n38601,n38565 );
   nor U40534 ( n39448,n37217,n28304 );
   not U40535 ( n38737,n38757 );
   nand U40536 ( n38757,n39532,n39533 );
   nand U40537 ( n39533,n37045,n39534 );
   nand U40538 ( n39534,n39535,n39536 );
   nor U40539 ( n39536,n39537,n39538 );
   nand U40540 ( n39538,n39539,n39540 );
   nand U40541 ( n39539,n39541,n39542 );
   nand U40542 ( n39542,n39543,n39544 );
   nand U40543 ( n39544,n37213,n27896 );
   nor U40544 ( n39541,n37113,n37052 );
   nor U40545 ( n39537,n39545,n39546 );
   nor U40546 ( n39546,n39547,n39548 );
   nor U40547 ( n39548,n39506,n37201 );
   nor U40548 ( n39547,n37052,n39549 );
   nor U40549 ( n39535,n39550,n37173 );
   nand U40550 ( n37173,n39551,n39552 );
   nor U40551 ( n39552,n39553,n39554 );
   nand U40552 ( n39554,n39516,n39555 );
   nand U40553 ( n39555,n39556,n37170 );
   nand U40554 ( n39516,n39557,n39558 );
   nor U40555 ( n39551,n39559,n39560 );
   nand U40556 ( n39560,n39561,n39562 );
   nand U40557 ( n39562,n37113,n39563 );
   nand U40558 ( n39563,n39564,n39565 );
   nor U40559 ( n39565,n39530,n37130 );
   nor U40560 ( n39564,n39566,n39567 );
   nor U40561 ( n39567,n38617,n38680 );
   nand U40562 ( n39561,n39568,n38649 );
   or U40563 ( n39568,n39569,n38680 );
   nor U40564 ( n39550,n37195,n39570 );
   nand U40565 ( n39570,n39571,n39572 );
   nand U40566 ( n39572,n37168,n39573 );
   nand U40567 ( n39571,n37166,n28280 );
   nand U40568 ( n39532,n39574,n27895 );
   nand U40569 ( n39478,n39575,p2_instaddrpointer_reg_26_ );
   nor U40570 ( n39575,n39331,n39353 );
   nand U40571 ( n39353,n39576,p2_instaddrpointer_reg_24_ );
   nor U40572 ( n39576,n39283,n39305 );
   nand U40573 ( n39305,n39490,n39258 );
   nor U40574 ( n39258,n39491,n39210 );
   nand U40575 ( n39210,n39577,p2_instaddrpointer_reg_18_ );
   nor U40576 ( n39577,n39140,n39162 );
   nand U40577 ( n39162,n39578,p2_instaddrpointer_reg_16_ );
   nor U40578 ( n39578,n39092,n39114 );
   nand U40579 ( n39114,n39494,n39073 );
   not U40580 ( n39073,n39066 );
   nand U40581 ( n39066,n39579,p2_instaddrpointer_reg_12_ );
   nor U40582 ( n39579,n38996,n39018 );
   not U40583 ( n39018,n39025 );
   nor U40584 ( n39025,n39496,n38970 );
   nand U40585 ( n38970,n39580,p2_instaddrpointer_reg_8_ );
   nor U40586 ( n39580,n38899,n38921 );
   nand U40587 ( n38921,n39581,p2_instaddrpointer_reg_6_ );
   nor U40588 ( n39581,n38851,n38873 );
   nand U40589 ( n38873,n39582,p2_instaddrpointer_reg_4_ );
   nor U40590 ( n39582,n38805,n38771 );
   or U40591 ( n38771,n38784,n38786 );
   nand U40592 ( n38784,p2_instaddrpointer_reg_1_,p2_instaddrpointer_reg_0_ );
   nor U40593 ( n39584,n39585,n39586 );
   nand U40594 ( n39586,n39587,n39588 );
   nand U40595 ( n39588,n38723,n28285 );
   nor U40596 ( n38723,n39590,n39591 );
   and U40597 ( n39591,n39592,n36762 );
   nand U40598 ( n39587,p2_phyaddrpointer_reg_0_,n39593 );
   nand U40599 ( n39593,n28381,n39595 );
   nor U40600 ( n39585,n38734,n39596 );
   nand U40601 ( n38734,n39597,n39598 );
   nand U40602 ( n39598,n39599,n36762 );
   nor U40603 ( n39583,n39600,n39601 );
   nor U40604 ( n39601,n39602,n39603 );
   nor U40605 ( n39600,n38726,n39604 );
   nor U40606 ( n39606,n39607,n39608 );
   nand U40607 ( n39608,n39609,n39610 );
   nand U40608 ( n39610,n28353,n38751 );
   xor U40609 ( n38751,n39612,n39613 );
   xor U40610 ( n39612,n36758,n39597 );
   nand U40611 ( n39609,n39589,n38753 );
   xor U40612 ( n38753,n39614,n39615 );
   xor U40613 ( n39614,n39590,p2_instaddrpointer_reg_1_ );
   nor U40614 ( n39607,n37125,n28124 );
   nor U40615 ( n39605,n39616,n39617 );
   nand U40616 ( n39617,n39618,n39619 );
   nand U40617 ( n39619,n39620,n39621 );
   nand U40618 ( n39618,n39622,p2_phyaddrpointer_reg_1_ );
   nor U40619 ( n39616,n36961,n39603 );
   nor U40620 ( n39624,n39625,n39626 );
   nand U40621 ( n39626,n39627,n39628 );
   nand U40622 ( n39628,n39611,n38777 );
   xor U40623 ( n38777,n39629,n39630 );
   xor U40624 ( n39630,p2_instaddrpointer_reg_2_,n39631 );
   nand U40625 ( n39627,n39589,n38778 );
   xor U40626 ( n38778,n39632,n39633 );
   xor U40627 ( n39632,n39634,p2_instaddrpointer_reg_2_ );
   nor U40628 ( n39625,n37189,n39604 );
   nor U40629 ( n39623,n39635,n39636 );
   nand U40630 ( n39636,n39637,n39638 );
   nand U40631 ( n39638,n39639,n28345 );
   nand U40632 ( n39637,n28347,p2_reip_reg_2_ );
   nor U40633 ( n39635,n39641,n28382 );
   nor U40634 ( n39643,n39644,n39645 );
   nand U40635 ( n39645,n39646,n39647 );
   nand U40636 ( n39647,n28353,n38794 );
   xor U40637 ( n38794,n39648,n39649 );
   or U40638 ( n39648,n39650,n39651 );
   and U40639 ( n39650,n39652,p2_instaddrpointer_reg_3_ );
   nand U40640 ( n39646,n39589,n38800 );
   xor U40641 ( n38800,n39653,n39654 );
   xor U40642 ( n39653,n39655,p2_instaddrpointer_reg_3_ );
   nor U40643 ( n39644,n37159,n28124 );
   nor U40644 ( n39642,n39656,n39657 );
   nand U40645 ( n39657,n39658,n39659 );
   nand U40646 ( n39659,n39620,n39660 );
   nand U40647 ( n39658,n39640,p2_reip_reg_3_ );
   nor U40648 ( n39656,n39661,n28382 );
   nor U40649 ( n39663,n39664,n39665 );
   nand U40650 ( n39665,n39666,n39667 );
   nand U40651 ( n39667,n28353,n38818 );
   xor U40652 ( n38818,n39668,n39669 );
   xor U40653 ( n39668,n38830,n39670 );
   nand U40654 ( n39666,n39589,n38819 );
   xor U40655 ( n38819,n39671,n39672 );
   xor U40656 ( n39671,n39673,p2_instaddrpointer_reg_4_ );
   nor U40657 ( n39664,n39674,n28123 );
   nor U40658 ( n39662,n39675,n39676 );
   nand U40659 ( n39676,n39677,n39678 );
   nand U40660 ( n39678,n39679,n28345 );
   nand U40661 ( n39677,n28347,p2_reip_reg_4_ );
   nor U40662 ( n39675,n39680,n39594 );
   nor U40663 ( n39682,n39683,n39684 );
   nand U40664 ( n39684,n39685,n39686 );
   nand U40665 ( n39686,n28353,n38845 );
   xor U40666 ( n38845,n39687,n39688 );
   and U40667 ( n39687,n39689,n39690 );
   nand U40668 ( n39685,n39589,n38846 );
   xor U40669 ( n38846,n39691,n39692 );
   xor U40670 ( n39691,n39693,p2_instaddrpointer_reg_5_ );
   nor U40671 ( n39683,n39694,n28124 );
   nor U40672 ( n39681,n39695,n39696 );
   nand U40673 ( n39696,n39697,n39698 );
   nand U40674 ( n39698,n39620,n39699 );
   nand U40675 ( n39697,n28347,p2_reip_reg_5_ );
   nor U40676 ( n39695,n39700,n28381 );
   nor U40677 ( n39702,n39703,n39704 );
   nand U40678 ( n39704,n39705,n39706 );
   nand U40679 ( n39706,n28353,n38864 );
   xor U40680 ( n38864,n39707,n39708 );
   xor U40681 ( n39707,n38877,n39709 );
   nand U40682 ( n39705,n39589,n38865 );
   xor U40683 ( n38865,n39710,n39711 );
   xor U40684 ( n39710,n39712,p2_instaddrpointer_reg_6_ );
   nor U40685 ( n39703,n39713,n39604 );
   nor U40686 ( n39701,n39714,n39715 );
   nand U40687 ( n39715,n39716,n39717 );
   nand U40688 ( n39717,n39718,n28345 );
   nand U40689 ( n39716,n28347,p2_reip_reg_6_ );
   nor U40690 ( n39714,n39719,n28381 );
   nor U40691 ( n39721,n39722,n39723 );
   nand U40692 ( n39723,n39724,n39725 );
   nand U40693 ( n39725,n28353,n38893 );
   xor U40694 ( n38893,n39726,n39727 );
   and U40695 ( n39726,n39728,n39729 );
   nand U40696 ( n39724,n39589,n38894 );
   xor U40697 ( n38894,n39730,n39731 );
   xor U40698 ( n39730,n39732,p2_instaddrpointer_reg_7_ );
   nor U40699 ( n39722,n39733,n28123 );
   nor U40700 ( n39720,n39734,n39735 );
   nand U40701 ( n39735,n39736,n39737 );
   nand U40702 ( n39737,n39620,n39738 );
   nand U40703 ( n39736,n28347,p2_reip_reg_7_ );
   nor U40704 ( n39734,n39739,n28382 );
   nor U40705 ( n39741,n39742,n39743 );
   nand U40706 ( n39743,n39744,n39745 );
   nand U40707 ( n39745,n39589,n38906 );
   xor U40708 ( n38906,n39746,n39747 );
   or U40709 ( n39746,n39748,n39749 );
   nand U40710 ( n39744,n28353,n38913 );
   xor U40711 ( n38913,n39750,n39751 );
   xor U40712 ( n39750,n38925,n39752 );
   nor U40713 ( n39742,n38908,n28124 );
   nor U40714 ( n39740,n39753,n39754 );
   nand U40715 ( n39754,n39755,n39756 );
   nand U40716 ( n39756,n39757,n28345 );
   nand U40717 ( n39755,n28347,p2_reip_reg_8_ );
   nor U40718 ( n39753,n39758,n28381 );
   nor U40719 ( n39760,n39761,n39762 );
   nand U40720 ( n39762,n39763,n39764 );
   nand U40721 ( n39764,n28353,n38935 );
   xor U40722 ( n38935,n39765,n39766 );
   and U40723 ( n39765,n39767,n39768 );
   nand U40724 ( n39763,n28285,n38936 );
   xor U40725 ( n38936,n39769,p2_instaddrpointer_reg_9_ );
   nor U40726 ( n39761,n39770,n39604 );
   nor U40727 ( n39759,n39771,n39772 );
   nand U40728 ( n39772,n39773,n39774 );
   nand U40729 ( n39774,n39620,n39775 );
   nand U40730 ( n39773,n28347,p2_reip_reg_9_ );
   nor U40731 ( n39771,n39776,n39594 );
   nor U40732 ( n39778,n39779,n39780 );
   nand U40733 ( n39780,n39781,n39782 );
   nand U40734 ( n39782,n38955,n28285 );
   nor U40735 ( n38955,n39783,n39784 );
   and U40736 ( n39784,n38974,n39785 );
   nand U40737 ( n39785,p2_instaddrpointer_reg_9_,n39769 );
   nand U40738 ( n39781,n28353,n38956 );
   xor U40739 ( n38956,n39786,n39787 );
   nand U40740 ( n39787,n39788,n39789 );
   nor U40741 ( n39779,n39790,n28123 );
   nor U40742 ( n39777,n39791,n39792 );
   nand U40743 ( n39792,n39793,n39794 );
   nand U40744 ( n39794,n39795,n28345 );
   nand U40745 ( n39793,n28347,p2_reip_reg_10_ );
   nor U40746 ( n39791,n39796,n39594 );
   nor U40747 ( n39798,n39799,n39800 );
   nand U40748 ( n39800,n39801,n39802 );
   nand U40749 ( n39802,n28353,n38984 );
   xor U40750 ( n38984,n39803,n39804 );
   nand U40751 ( n39804,n39788,n39805 );
   nand U40752 ( n39805,n39786,n39789 );
   not U40753 ( n39786,n39806 );
   nand U40754 ( n39803,n39807,n39808 );
   nand U40755 ( n39801,n28285,n38985 );
   xor U40756 ( n38985,p2_instaddrpointer_reg_11_,n39783 );
   nor U40757 ( n39799,n39809,n28124 );
   nor U40758 ( n39797,n39810,n39811 );
   nand U40759 ( n39811,n39812,n39813 );
   nand U40760 ( n39813,n39620,n39814 );
   nand U40761 ( n39812,n28347,p2_reip_reg_11_ );
   nor U40762 ( n39810,n39815,n28381 );
   nor U40763 ( n39817,n39818,n39819 );
   nand U40764 ( n39819,n39820,n39821 );
   nand U40765 ( n39821,n28353,n39009 );
   nand U40766 ( n39009,n39822,n39823 );
   nand U40767 ( n39823,n39824,n39825 );
   nand U40768 ( n39824,n39826,n39827 );
   nand U40769 ( n39822,n39828,n39826 );
   nand U40770 ( n39820,n39589,n39010 );
   xor U40771 ( n39010,n39022,n39829 );
   nand U40772 ( n39829,n39783,p2_instaddrpointer_reg_11_ );
   nor U40773 ( n39783,n39496,n39830 );
   nor U40774 ( n39818,n39831,n28124 );
   nor U40775 ( n39816,n39832,n39833 );
   nand U40776 ( n39833,n39834,n39835 );
   nand U40777 ( n39835,n39836,n28345 );
   nand U40778 ( n39834,n28347,p2_reip_reg_12_ );
   nor U40779 ( n39832,n39837,n28382 );
   nor U40780 ( n39839,n39840,n39841 );
   nand U40781 ( n39841,n39842,n39843 );
   nand U40782 ( n39843,n39032,n28285 );
   nor U40783 ( n39032,n39844,n39845 );
   and U40784 ( n39845,n39043,n39846 );
   or U40785 ( n39846,n39847,n39830 );
   not U40786 ( n39844,n39848 );
   nand U40787 ( n39842,n28353,n39039 );
   xor U40788 ( n39039,n39849,n39850 );
   nand U40789 ( n39850,n39826,n39851 );
   not U40790 ( n39851,n39828 );
   nor U40791 ( n39828,n39825,n39852 );
   not U40792 ( n39852,n39827 );
   nand U40793 ( n39849,n39853,n39854 );
   nor U40794 ( n39840,n39034,n28123 );
   nor U40795 ( n39838,n39855,n39856 );
   nand U40796 ( n39856,n39857,n39858 );
   nand U40797 ( n39858,n39620,n39859 );
   nand U40798 ( n39857,n28347,p2_reip_reg_13_ );
   nor U40799 ( n39855,n39860,n28382 );
   nor U40800 ( n39862,n39863,n39864 );
   nand U40801 ( n39864,n39865,n39866 );
   nand U40802 ( n39866,n39589,n39051 );
   xor U40803 ( n39051,n39070,n39848 );
   nand U40804 ( n39865,n28353,n39058 );
   nand U40805 ( n39058,n39867,n39868 );
   nand U40806 ( n39868,n39869,n39870 );
   nand U40807 ( n39869,n39871,n39872 );
   nand U40808 ( n39867,n39873,n39871 );
   not U40809 ( n39873,n39874 );
   nor U40810 ( n39863,n39053,n39604 );
   nor U40811 ( n39861,n39875,n39876 );
   nand U40812 ( n39876,n39877,n39878 );
   nand U40813 ( n39878,n39879,n28345 );
   nand U40814 ( n39877,n39640,p2_reip_reg_14_ );
   nor U40815 ( n39875,n39880,n39594 );
   nor U40816 ( n39882,n39883,n39884 );
   nand U40817 ( n39884,n39885,n39886 );
   nand U40818 ( n39886,n28353,n39086 );
   xor U40819 ( n39086,n39887,n39888 );
   nand U40820 ( n39888,n39889,n39890 );
   nand U40821 ( n39887,n39874,n39871 );
   nand U40822 ( n39874,n39891,n39872 );
   not U40823 ( n39891,n39870 );
   nand U40824 ( n39885,n39589,n39087 );
   xor U40825 ( n39087,n39892,p2_instaddrpointer_reg_15_ );
   nor U40826 ( n39892,n39070,n39848 );
   nand U40827 ( n39848,n39893,p2_instaddrpointer_reg_13_ );
   nor U40828 ( n39893,n39830,n39847 );
   nor U40829 ( n39883,n39894,n39604 );
   nor U40830 ( n39881,n39895,n39896 );
   nand U40831 ( n39896,n39897,n39898 );
   nand U40832 ( n39898,n39620,n39899 );
   nand U40833 ( n39897,n39640,p2_reip_reg_15_ );
   nor U40834 ( n39895,n39900,n39594 );
   nor U40835 ( n39902,n39903,n39904 );
   nand U40836 ( n39904,n39905,n39906 );
   nand U40837 ( n39906,n39099,n28285 );
   nor U40838 ( n39099,n39907,n39908 );
   and U40839 ( n39908,n39118,n39909 );
   or U40840 ( n39909,n39910,n39830 );
   not U40841 ( n39907,n39911 );
   nand U40842 ( n39905,n39611,n39106 );
   nand U40843 ( n39106,n39912,n39913 );
   nand U40844 ( n39913,n39914,n39915 );
   nand U40845 ( n39914,n39916,n39917 );
   nand U40846 ( n39912,n39918,n39916 );
   not U40847 ( n39918,n39919 );
   nor U40848 ( n39903,n39101,n28123 );
   nor U40849 ( n39901,n39920,n39921 );
   nand U40850 ( n39921,n39922,n39923 );
   nand U40851 ( n39923,n39924,n28345 );
   nand U40852 ( n39922,n39640,p2_reip_reg_16_ );
   nor U40853 ( n39920,n39925,n28382 );
   nor U40854 ( n39927,n39928,n39929 );
   nand U40855 ( n39929,n39930,n39931 );
   nand U40856 ( n39931,n39589,n39128 );
   xor U40857 ( n39128,n39140,n39911 );
   nand U40858 ( n39930,n39611,n39135 );
   xor U40859 ( n39135,n39932,n39933 );
   nand U40860 ( n39933,n39934,n39935 );
   nand U40861 ( n39932,n39919,n39916 );
   nand U40862 ( n39919,n39936,n39917 );
   not U40863 ( n39936,n39915 );
   nor U40864 ( n39928,n39130,n28124 );
   nor U40865 ( n39926,n39937,n39938 );
   nand U40866 ( n39938,n39939,n39940 );
   nand U40867 ( n39940,n39620,n39941 );
   nand U40868 ( n39939,n39640,p2_reip_reg_17_ );
   nor U40869 ( n39937,n39942,n28382 );
   nor U40870 ( n39944,n39945,n39946 );
   nand U40871 ( n39946,n39947,n39948 );
   nand U40872 ( n39948,n39611,n39147 );
   xor U40873 ( n39147,n39949,n39950 );
   and U40874 ( n39949,n39951,n39952 );
   nand U40875 ( n39947,n28285,n39154 );
   xor U40876 ( n39154,n39953,p2_instaddrpointer_reg_18_ );
   nor U40877 ( n39953,n39140,n39911 );
   nand U40878 ( n39911,n39954,p2_instaddrpointer_reg_16_ );
   nor U40879 ( n39954,n39830,n39910 );
   nor U40880 ( n39945,n39149,n28124 );
   nor U40881 ( n39943,n39955,n39956 );
   nand U40882 ( n39956,n39957,n39958 );
   nand U40883 ( n39958,n39959,n28345 );
   nand U40884 ( n39957,n39640,p2_reip_reg_18_ );
   nor U40885 ( n39955,n39960,n28382 );
   nor U40886 ( n39962,n39963,n39964 );
   nand U40887 ( n39964,n39965,n39966 );
   nand U40888 ( n39966,n39611,n39176 );
   xor U40889 ( n39176,n39967,n39968 );
   nand U40890 ( n39968,n39951,n39969 );
   nand U40891 ( n39969,n39952,n39950 );
   nor U40892 ( n39967,n39970,n39971 );
   and U40893 ( n39971,n39972,n39188 );
   nand U40894 ( n39965,n28285,n39183 );
   and U40895 ( n39183,n39973,n39974 );
   nand U40896 ( n39974,n39975,n39188 );
   nor U40897 ( n39963,n39178,n28123 );
   nor U40898 ( n39961,n39976,n39977 );
   nand U40899 ( n39977,n39978,n39979 );
   nand U40900 ( n39979,n39620,n39980 );
   nand U40901 ( n39978,n39640,p2_reip_reg_19_ );
   nor U40902 ( n39976,n39981,n39594 );
   nor U40903 ( n39983,n39984,n39985 );
   nand U40904 ( n39985,n39986,n39987 );
   nand U40905 ( n39987,n39195,n28285 );
   nor U40906 ( n39195,n39988,n39989 );
   and U40907 ( n39989,n39212,n39973 );
   or U40908 ( n39973,n39975,n39188 );
   nand U40909 ( n39986,n39611,n39202 );
   not U40910 ( n39202,n39990 );
   xor U40911 ( n39990,n39991,n39992 );
   nand U40912 ( n39992,n39993,n39994 );
   nor U40913 ( n39984,n39197,n39604 );
   nor U40914 ( n39982,n39995,n39996 );
   nand U40915 ( n39996,n39997,n39998 );
   nand U40916 ( n39998,n39999,n28345 );
   nand U40917 ( n39997,n39640,p2_reip_reg_20_ );
   nor U40918 ( n39995,n40000,n28381 );
   nor U40919 ( n40002,n40003,n40004 );
   nand U40920 ( n40004,n40005,n40006 );
   nand U40921 ( n40006,n28285,n39222 );
   xor U40922 ( n39222,p2_instaddrpointer_reg_21_,n39988 );
   nand U40923 ( n40005,n39611,n39229 );
   xor U40924 ( n39229,n40007,n40008 );
   nand U40925 ( n40008,n40009,n40010 );
   nor U40926 ( n40003,n39224,n39604 );
   nor U40927 ( n40001,n40011,n40012 );
   nand U40928 ( n40012,n40013,n40014 );
   nand U40929 ( n40014,n39620,n40015 );
   nand U40930 ( n40013,n39640,p2_reip_reg_21_ );
   nor U40931 ( n40011,n40016,n28381 );
   nor U40932 ( n40018,n40019,n40020 );
   nand U40933 ( n40020,n40021,n40022 );
   nand U40934 ( n40022,n39611,n39247 );
   nand U40935 ( n39247,n40023,n40024 );
   nand U40936 ( n40024,n40025,n40026 );
   nor U40937 ( n40023,n40027,n40028 );
   nor U40938 ( n40028,n39261,n40029 );
   xor U40939 ( n40029,n40026,n40030 );
   not U40940 ( n40026,n40031 );
   nor U40941 ( n40027,p2_instaddrpointer_reg_22_,n40032 );
   nand U40942 ( n40032,n40030,n40031 );
   nand U40943 ( n40031,n40009,n40033 );
   nand U40944 ( n40033,n40007,n40010 );
   not U40945 ( n40007,n40034 );
   nand U40946 ( n40021,n28285,n39248 );
   and U40947 ( n39248,n40035,n40036 );
   nand U40948 ( n40036,n40037,n39261 );
   nand U40949 ( n40037,n39988,p2_instaddrpointer_reg_21_ );
   nor U40950 ( n40019,n40038,n28123 );
   nor U40951 ( n40017,n40039,n40040 );
   nand U40952 ( n40040,n40041,n40042 );
   nand U40953 ( n40042,n40043,n28345 );
   nand U40954 ( n40041,n39640,p2_reip_reg_22_ );
   nor U40955 ( n40039,n40044,n39594 );
   nor U40956 ( n40046,n40047,n40048 );
   nand U40957 ( n40048,n40049,n40050 );
   nand U40958 ( n40050,n39271,n28285 );
   nor U40959 ( n39271,n40051,n40052 );
   and U40960 ( n40052,n39283,n40035 );
   nand U40961 ( n40049,n39611,n39278 );
   xor U40962 ( n39278,n40053,n40054 );
   nand U40963 ( n40054,n40055,n40056 );
   nor U40964 ( n40047,n39273,n28124 );
   nor U40965 ( n40045,n40057,n40058 );
   nand U40966 ( n40058,n40059,n40060 );
   nand U40967 ( n40060,n39620,n40061 );
   nand U40968 ( n40059,n39640,p2_reip_reg_23_ );
   nor U40969 ( n40057,n40062,n28382 );
   nor U40970 ( n40064,n40065,n40066 );
   nand U40971 ( n40066,n40067,n40068 );
   nand U40972 ( n40068,n28285,n39290 );
   xor U40973 ( n39290,n39309,n40069 );
   nand U40974 ( n40067,n39611,n39297 );
   nand U40975 ( n39297,n40070,n40071 );
   nand U40976 ( n40071,n40072,n40073 );
   nor U40977 ( n40070,n40074,n40075 );
   nor U40978 ( n40075,n39309,n40076 );
   xor U40979 ( n40076,n40073,n40077 );
   not U40980 ( n40073,n40078 );
   nor U40981 ( n40074,p2_instaddrpointer_reg_24_,n40079 );
   nand U40982 ( n40079,n40077,n40078 );
   nand U40983 ( n40078,n40055,n40080 );
   nand U40984 ( n40080,n40053,n40056 );
   not U40985 ( n40053,n40081 );
   nor U40986 ( n40065,n39292,n39604 );
   nor U40987 ( n40063,n40082,n40083 );
   nand U40988 ( n40083,n40084,n40085 );
   nand U40989 ( n40085,n40086,n28345 );
   nand U40990 ( n40084,n39640,p2_reip_reg_24_ );
   nor U40991 ( n40082,n40087,n28382 );
   nor U40992 ( n40089,n40090,n40091 );
   nand U40993 ( n40091,n40092,n40093 );
   nand U40994 ( n40093,n39611,n39325 );
   xor U40995 ( n39325,n40094,n40095 );
   xor U40996 ( n40094,n39331,n40096 );
   nand U40997 ( n40092,n28285,n39326 );
   xor U40998 ( n39326,n40097,p2_instaddrpointer_reg_25_ );
   nor U40999 ( n40097,n39309,n40069 );
   nor U41000 ( n40090,n40098,n28123 );
   nor U41001 ( n40088,n40099,n40100 );
   nand U41002 ( n40100,n40101,n40102 );
   nand U41003 ( n40102,n39620,n40103 );
   nand U41004 ( n40101,n39640,p2_reip_reg_25_ );
   nor U41005 ( n40099,n40104,n39594 );
   nor U41006 ( n40106,n40107,n40108 );
   nand U41007 ( n40108,n40109,n40110 );
   nand U41008 ( n40110,n39611,n39338 );
   xor U41009 ( n39338,n40111,n40112 );
   nor U41010 ( n40111,n40113,n40114 );
   not U41011 ( n40114,n40115 );
   nor U41012 ( n40113,p2_instaddrpointer_reg_26_,n40116 );
   nand U41013 ( n40109,n39589,n39345 );
   nand U41014 ( n39345,n40117,n40118 );
   nand U41015 ( n40118,n40119,n40120 );
   nor U41016 ( n40120,n40121,n39309 );
   nor U41017 ( n40119,n40069,n39331 );
   not U41018 ( n40069,n40051 );
   nor U41019 ( n40051,n39283,n40035 );
   nand U41020 ( n40035,n39490,n39988 );
   nor U41021 ( n39988,n39491,n39975 );
   nand U41022 ( n39975,n40122,n39769 );
   not U41023 ( n39491,n39259 );
   nand U41024 ( n40117,p2_instaddrpointer_reg_26_,n40123 );
   nor U41025 ( n40107,n39340,n28124 );
   nor U41026 ( n40105,n40124,n40125 );
   nand U41027 ( n40125,n40126,n40127 );
   nand U41028 ( n40127,n40128,n28345 );
   nand U41029 ( n40126,n39640,p2_reip_reg_26_ );
   nor U41030 ( n40124,n40129,n28381 );
   nor U41031 ( n40131,n40132,n40133 );
   nand U41032 ( n40133,n40134,n40135 );
   nand U41033 ( n40135,n39589,n39367 );
   xor U41034 ( n39367,n39379,n40123 );
   nand U41035 ( n40134,n39611,n39374 );
   xor U41036 ( n39374,n40136,n40137 );
   and U41037 ( n40136,n40138,n40139 );
   nor U41038 ( n40132,n39369,n39604 );
   nor U41039 ( n40130,n40140,n40141 );
   nand U41040 ( n40141,n40142,n40143 );
   nand U41041 ( n40143,n39620,n40144 );
   nand U41042 ( n40142,n39640,p2_reip_reg_27_ );
   nor U41043 ( n40140,n40145,n28381 );
   nor U41044 ( n40147,n40148,n40149 );
   nand U41045 ( n40149,n40150,n40151 );
   nand U41046 ( n40151,n39611,n39392 );
   xor U41047 ( n39392,n40152,n40153 );
   and U41048 ( n40152,n40154,n40155 );
   nand U41049 ( n40150,n39589,n39393 );
   and U41050 ( n39393,n40156,n40157 );
   nand U41051 ( n40157,n40158,n39396 );
   nor U41052 ( n40148,n40159,n28123 );
   nor U41053 ( n40146,n40160,n40161 );
   nand U41054 ( n40161,n40162,n40163 );
   nand U41055 ( n40163,n40164,n28345 );
   nand U41056 ( n40162,n39640,p2_reip_reg_28_ );
   nor U41057 ( n40160,n40165,n39594 );
   nor U41058 ( n40167,n40168,n40169 );
   nand U41059 ( n40169,n40170,n40171 );
   nand U41060 ( n40171,n39405,n28285 );
   nor U41061 ( n39405,n40172,n40173 );
   nor U41062 ( n40173,p2_instaddrpointer_reg_29_,n40174 );
   nand U41063 ( n40170,n39611,n39412 );
   xor U41064 ( n39412,n40175,n40176 );
   and U41065 ( n40175,n40177,n40178 );
   nor U41066 ( n40168,n39407,n39604 );
   nor U41067 ( n40166,n40179,n40180 );
   nand U41068 ( n40180,n40181,n40182 );
   nand U41069 ( n40182,n39620,n40183 );
   nand U41070 ( n40181,n39640,p2_reip_reg_29_ );
   nor U41071 ( n40179,n40184,n39594 );
   nor U41072 ( n40186,n40187,n40188 );
   nand U41073 ( n40188,n40189,n40190 );
   or U41074 ( n40190,n28123,n40191 );
   nand U41075 ( n40189,n28353,n39425 );
   xor U41076 ( n39425,n40192,n40193 );
   nand U41077 ( n40193,n40194,n40195 );
   not U41078 ( n39611,n39596 );
   nor U41079 ( n40187,n39426,n40196 );
   not U41080 ( n40196,n39589 );
   xor U41081 ( n39426,n39435,n40172 );
   nor U41082 ( n40185,n40197,n40198 );
   nand U41083 ( n40198,n40199,n40200 );
   nand U41084 ( n40200,n40201,n28345 );
   nand U41085 ( n40199,n28347,p2_reip_reg_30_ );
   not U41086 ( n39640,n39603 );
   nor U41087 ( n40197,n40202,n28381 );
   nor U41088 ( n40204,n40205,n40206 );
   nand U41089 ( n40206,n40207,n40208 );
   nand U41090 ( n40208,n40209,n39446 );
   nor U41091 ( n39446,n40210,n40211 );
   and U41092 ( n40211,n40212,n40213 );
   nand U41093 ( n40213,n40214,n40194 );
   nand U41094 ( n40214,n40215,n40216 );
   nand U41095 ( n40216,n40178,n40176 );
   and U41096 ( n40215,n40177,n40195 );
   nor U41097 ( n40210,n40195,n40212 );
   nand U41098 ( n40195,n40217,n40218 );
   nor U41099 ( n40217,n28370,n39435 );
   nor U41100 ( n40209,n39447,n39596 );
   nand U41101 ( n39596,n40220,n39594 );
   nor U41102 ( n39447,n40221,n40192 );
   nand U41103 ( n40192,n40178,n40222 );
   nand U41104 ( n40222,n40223,n40177 );
   nand U41105 ( n40177,n40224,n40225 );
   nor U41106 ( n40224,n28371,n39416 );
   not U41107 ( n40223,n40176 );
   nand U41108 ( n40176,n40154,n40226 );
   nand U41109 ( n40226,n40153,n40155 );
   nand U41110 ( n40155,n39396,n40227 );
   nand U41111 ( n40227,n40228,n28282 );
   nand U41112 ( n40153,n40138,n40230 );
   nand U41113 ( n40230,n40137,n40139 );
   nand U41114 ( n40139,n39379,n40231 );
   nand U41115 ( n40231,n40232,n28282 );
   nand U41116 ( n40137,n40233,n40115 );
   nand U41117 ( n40115,n40116,p2_instaddrpointer_reg_26_ );
   nor U41118 ( n40116,n28371,n40234 );
   nand U41119 ( n40233,n40112,n40235 );
   nand U41120 ( n40235,n39357,n40236 );
   nand U41121 ( n40236,n40237,n40229 );
   and U41122 ( n40112,n40238,n40239 );
   nand U41123 ( n40239,n40240,n39331 );
   nand U41124 ( n40240,n40241,n40096 );
   or U41125 ( n40238,n40096,n40241 );
   not U41126 ( n40241,n40095 );
   nand U41127 ( n40095,n40242,n40243 );
   nor U41128 ( n40242,n40219,n40244 );
   nand U41129 ( n40096,n40245,n40246 );
   nand U41130 ( n40246,n40247,n40248 );
   not U41131 ( n40248,n40072 );
   nor U41132 ( n40072,p2_instaddrpointer_reg_24_,n40077 );
   nand U41133 ( n40247,n40056,n40249 );
   nand U41134 ( n40249,n40055,n40081 );
   nand U41135 ( n40081,n40250,n40251 );
   nand U41136 ( n40251,n40252,n40253 );
   not U41137 ( n40253,n40025 );
   nor U41138 ( n40025,p2_instaddrpointer_reg_22_,n40030 );
   nand U41139 ( n40252,n40010,n40254 );
   nand U41140 ( n40254,n40009,n40034 );
   nand U41141 ( n40034,n39994,n40255 );
   nand U41142 ( n40255,n39991,n39993 );
   nand U41143 ( n39993,n40256,n39212 );
   nand U41144 ( n39991,n40257,n40258 );
   nand U41145 ( n40258,n40259,n40260 );
   nand U41146 ( n40259,n39951,n40261 );
   not U41147 ( n40261,n39970 );
   nor U41148 ( n39970,n39188,n39972 );
   nand U41149 ( n39951,n40262,p2_instaddrpointer_reg_18_ );
   and U41150 ( n40262,n40229,n40263 );
   nand U41151 ( n40257,n40264,n40260 );
   nand U41152 ( n40260,n39972,n39188 );
   nand U41153 ( n39972,n40265,n40266 );
   nor U41154 ( n40265,n28371,n40267 );
   and U41155 ( n40264,n39950,n39952 );
   nand U41156 ( n39952,n39166,n40268 );
   nand U41157 ( n40268,n40263,n40229 );
   nand U41158 ( n39950,n39935,n40269 );
   nand U41159 ( n40269,n40270,n39934 );
   nand U41160 ( n39934,n39140,n40271 );
   nand U41161 ( n40271,n40272,n28282 );
   nand U41162 ( n40270,n39917,n40273 );
   nand U41163 ( n40273,n39915,n39916 );
   nand U41164 ( n39916,n39118,n40274 );
   nand U41165 ( n40274,n40275,n40229 );
   nand U41166 ( n39915,n39890,n40276 );
   nand U41167 ( n40276,n40277,n39889 );
   nand U41168 ( n39889,n39092,n40278 );
   nand U41169 ( n40278,n40279,n28282 );
   nand U41170 ( n40277,n39872,n40280 );
   nand U41171 ( n40280,n39870,n39871 );
   nand U41172 ( n39871,n39070,n40281 );
   nand U41173 ( n40281,n40282,n40229 );
   nand U41174 ( n39870,n39853,n40283 );
   nand U41175 ( n40283,n40284,n39854 );
   nand U41176 ( n39854,n39043,n40285 );
   nand U41177 ( n40285,n40286,n28282 );
   nand U41178 ( n40284,n39827,n40287 );
   nand U41179 ( n40287,n39825,n39826 );
   nand U41180 ( n39826,n39022,n40288 );
   nand U41181 ( n40288,n40289,n28282 );
   nand U41182 ( n39825,n39807,n40290 );
   nand U41183 ( n40290,n40291,n39808 );
   nand U41184 ( n39808,n40292,n38996 );
   nand U41185 ( n40292,n40293,n40229 );
   nand U41186 ( n40291,n39789,n40294 );
   nand U41187 ( n40294,n39788,n39806 );
   nand U41188 ( n39806,n39767,n40295 );
   nand U41189 ( n40295,n39766,n39768 );
   nand U41190 ( n39768,n38948,n40296 );
   nand U41191 ( n40296,n40297,n40229 );
   and U41192 ( n39766,n40298,n40299 );
   nand U41193 ( n40299,n40300,n38925 );
   nand U41194 ( n40300,n40301,n39752 );
   or U41195 ( n40298,n39752,n40301 );
   not U41196 ( n40301,n39751 );
   nand U41197 ( n39751,n40302,n40303 );
   nand U41198 ( n40303,n40219,n40304 );
   nand U41199 ( n40302,n40305,n40229 );
   xor U41200 ( n40305,n40306,n40307 );
   nand U41201 ( n39752,n39729,n40308 );
   nand U41202 ( n40308,n39727,n39728 );
   or U41203 ( n39728,n40309,p2_instaddrpointer_reg_7_ );
   and U41204 ( n39727,n40310,n40311 );
   nand U41205 ( n40311,n40312,n38877 );
   nand U41206 ( n40312,n40313,n39709 );
   or U41207 ( n40310,n39709,n40313 );
   not U41208 ( n40313,n39708 );
   nand U41209 ( n39708,n40314,n40315 );
   nand U41210 ( n40315,n28371,n39712 );
   nand U41211 ( n40314,n40316,n28282 );
   xor U41212 ( n40316,n40317,n40318 );
   nand U41213 ( n39709,n39690,n40319 );
   nand U41214 ( n40319,n39688,n39689 );
   or U41215 ( n39689,n40320,p2_instaddrpointer_reg_5_ );
   and U41216 ( n39688,n40321,n40322 );
   nand U41217 ( n40322,n40323,n38830 );
   nand U41218 ( n40323,n40324,n39670 );
   or U41219 ( n40321,n39670,n40324 );
   not U41220 ( n40324,n39669 );
   nand U41221 ( n39669,n40325,n40326 );
   nand U41222 ( n40326,n40327,n28282 );
   xor U41223 ( n40327,n40328,n40329 );
   nand U41224 ( n40325,n39672,n28371 );
   nand U41225 ( n39670,n40330,n40331 );
   nand U41226 ( n40331,p2_instaddrpointer_reg_3_,n39652 );
   or U41227 ( n40330,n39649,n39651 );
   nor U41228 ( n39651,n39652,p2_instaddrpointer_reg_3_ );
   nand U41229 ( n39652,n40332,n40333 );
   nand U41230 ( n40333,n40334,n28282 );
   nand U41231 ( n40332,n39654,n28370 );
   nand U41232 ( n39649,n40335,n40336 );
   nand U41233 ( n40336,n40337,n38786 );
   or U41234 ( n40337,n39629,n39631 );
   nand U41235 ( n40335,n39629,n39631 );
   nand U41236 ( n39631,n40338,n40339 );
   nand U41237 ( n40339,n40340,n36758 );
   nand U41238 ( n40340,n39613,n40341 );
   not U41239 ( n39613,n40342 );
   nand U41240 ( n40338,n40342,n39597 );
   not U41241 ( n39597,n40341 );
   nor U41242 ( n40341,n39599,n36762 );
   nand U41243 ( n39599,n40343,n40344 );
   nand U41244 ( n40344,n40229,n40345 );
   nand U41245 ( n40343,n39592,n28370 );
   nand U41246 ( n40342,n40346,n40347 );
   nand U41247 ( n40347,n40348,n40229 );
   or U41248 ( n40346,n39615,n40229 );
   nand U41249 ( n39629,n40349,n40350 );
   nand U41250 ( n40350,n40351,n40229 );
   nand U41251 ( n40351,n40352,n40353 );
   nand U41252 ( n40353,n40354,n40355 );
   nand U41253 ( n40349,n39633,n28370 );
   nand U41254 ( n39690,p2_instaddrpointer_reg_5_,n40320 );
   nand U41255 ( n40320,n40356,n40357 );
   nand U41256 ( n40357,n40358,n40229 );
   and U41257 ( n40358,n40359,n40360 );
   nand U41258 ( n40356,n39693,n40219 );
   nand U41259 ( n39729,p2_instaddrpointer_reg_7_,n40309 );
   nand U41260 ( n40309,n40361,n40362 );
   nand U41261 ( n40362,n40363,n40229 );
   and U41262 ( n40363,n40364,n40365 );
   nand U41263 ( n40361,n39732,n28371 );
   nand U41264 ( n39767,n40366,p2_instaddrpointer_reg_9_ );
   nor U41265 ( n40366,n40219,n40367 );
   nand U41266 ( n39788,n38974,n40368 );
   nand U41267 ( n40368,n40369,n28282 );
   nand U41268 ( n39789,n40370,n40369 );
   nor U41269 ( n40370,n40219,n38974 );
   nand U41270 ( n39807,n40371,p2_instaddrpointer_reg_11_ );
   nor U41271 ( n40371,n28370,n40372 );
   nand U41272 ( n39827,n40373,n40289 );
   nor U41273 ( n40373,n28371,n39022 );
   nand U41274 ( n39853,n40374,n40286 );
   nor U41275 ( n40374,n28370,n39043 );
   nand U41276 ( n39872,n40375,n40282 );
   nor U41277 ( n40375,n40219,n39070 );
   nand U41278 ( n39890,n40376,n40279 );
   nor U41279 ( n40376,n28370,n39092 );
   nand U41280 ( n39917,n40377,n40275 );
   nor U41281 ( n40377,n40219,n39118 );
   nand U41282 ( n39935,n40378,n40272 );
   nor U41283 ( n40378,n28371,n39140 );
   or U41284 ( n39994,n40256,n39212 );
   nand U41285 ( n40256,n40379,n28282 );
   nand U41286 ( n40009,n39234,n40380 );
   nand U41287 ( n40380,n40381,n40382 );
   nand U41288 ( n40010,n40383,n40381 );
   nor U41289 ( n40381,n28371,n40384 );
   nor U41290 ( n40383,n40385,n39234 );
   nand U41291 ( n40250,n40030,p2_instaddrpointer_reg_22_ );
   and U41292 ( n40030,n40386,n40229 );
   nand U41293 ( n40055,n39283,n40387 );
   nand U41294 ( n40387,n40388,n40389 );
   nand U41295 ( n40056,n40390,n40388 );
   nor U41296 ( n40388,n40219,n40391 );
   nor U41297 ( n40390,n40392,n39283 );
   nand U41298 ( n40245,n40077,p2_instaddrpointer_reg_24_ );
   and U41299 ( n40077,n40393,n40229 );
   nand U41300 ( n40138,n40394,n40232 );
   nor U41301 ( n40394,n28370,n39379 );
   nand U41302 ( n40154,n40395,n40228 );
   nor U41303 ( n40395,n28370,n39396 );
   nand U41304 ( n40178,n39416,n40396 );
   nand U41305 ( n40396,n40225,n40229 );
   nand U41306 ( n40221,n40194,n40397 );
   not U41307 ( n40397,n40212 );
   xor U41308 ( n40212,n40398,n39482 );
   nor U41309 ( n40398,n28361,n40400 );
   nand U41310 ( n40400,n40401,n28282 );
   nand U41311 ( n40194,n39435,n40402 );
   nand U41312 ( n40402,n40218,n40229 );
   nand U41313 ( n40207,n39589,n39449 );
   xor U41314 ( n39449,n40403,p2_instaddrpointer_reg_31_ );
   and U41315 ( n40403,p2_instaddrpointer_reg_30_,n40172 );
   nor U41316 ( n40172,n39416,n40156 );
   not U41317 ( n40156,n40174 );
   nor U41318 ( n40174,n40158,n39396 );
   or U41319 ( n40158,n40123,n39379 );
   nand U41320 ( n40123,n40121,n39769 );
   not U41321 ( n39769,n39830 );
   nor U41322 ( n39830,n39748,n40404 );
   nor U41323 ( n40404,n39747,n39749 );
   nor U41324 ( n39749,p2_instaddrpointer_reg_8_,n40405 );
   nand U41325 ( n39747,n40406,n40407 );
   nand U41326 ( n40407,n40408,n38899 );
   nand U41327 ( n40408,n39731,n39732 );
   not U41328 ( n39732,n40409 );
   not U41329 ( n39731,n40410 );
   nand U41330 ( n40406,n40410,n40409 );
   nand U41331 ( n40409,n40304,n40411 );
   nand U41332 ( n40411,n40412,n40413 );
   nand U41333 ( n40410,n40414,n40415 );
   nand U41334 ( n40415,n40416,n38877 );
   or U41335 ( n40416,n39711,n39712 );
   nand U41336 ( n40414,n39711,n39712 );
   nand U41337 ( n39712,n40413,n40417 );
   nand U41338 ( n40417,n40418,n40419 );
   nand U41339 ( n39711,n40420,n40421 );
   nand U41340 ( n40421,n40422,n38851 );
   nand U41341 ( n40422,n39692,n39693 );
   not U41342 ( n39693,n40423 );
   not U41343 ( n39692,n40424 );
   nand U41344 ( n40420,n40424,n40423 );
   nand U41345 ( n40423,n40419,n40425 );
   nand U41346 ( n40425,n40426,n40427 );
   nand U41347 ( n40427,n40428,n40429 );
   nand U41348 ( n40424,n40430,n40431 );
   nand U41349 ( n40431,n40432,n38830 );
   or U41350 ( n40432,n39673,n39672 );
   nand U41351 ( n40430,n39672,n39673 );
   nand U41352 ( n39673,n40433,n40434 );
   nand U41353 ( n40434,n40435,n38805 );
   nand U41354 ( n40435,n39655,n39654 );
   or U41355 ( n40433,n39654,n39655 );
   and U41356 ( n39655,n40436,n40437 );
   nand U41357 ( n40437,n40438,n38786 );
   or U41358 ( n40438,n39634,n39633 );
   nand U41359 ( n40436,n39633,n39634 );
   nand U41360 ( n39634,n40439,n40440 );
   nand U41361 ( n40440,n40441,n36758 );
   nand U41362 ( n40441,n39615,n39590 );
   or U41363 ( n40439,n39615,n39590 );
   nor U41364 ( n39590,n36762,n39592 );
   xor U41365 ( n39592,n36646,n40442 );
   xor U41366 ( n39615,n40443,n40444 );
   xor U41367 ( n39633,n40445,n40446 );
   xor U41368 ( n40446,n36646,n40447 );
   xor U41369 ( n39654,n40448,n40449 );
   xor U41370 ( n39672,n40428,n40450 );
   nor U41371 ( n39748,n38925,n40304 );
   not U41372 ( n40304,n40405 );
   nor U41373 ( n40405,n40413,n40412 );
   and U41374 ( n40412,n28371,n40451 );
   nand U41375 ( n40451,n40452,n28280 );
   nand U41376 ( n40452,n40453,n40454 );
   nor U41377 ( n40454,n40455,n40456 );
   nand U41378 ( n40456,n40457,n40458 );
   nor U41379 ( n40458,n40459,n40460 );
   nor U41380 ( n40460,n40461,n37423 );
   nor U41381 ( n40459,n40462,n37511 );
   nor U41382 ( n40457,n40463,n40464 );
   nor U41383 ( n40464,n40465,n37597 );
   nor U41384 ( n40463,n40466,n37774 );
   nand U41385 ( n40455,n40467,n40468 );
   nor U41386 ( n40468,n40469,n40470 );
   nor U41387 ( n40470,n40471,n37857 );
   nor U41388 ( n40469,n40472,n37941 );
   nor U41389 ( n40467,n40473,n40474 );
   nor U41390 ( n40474,n40475,n38111 );
   nor U41391 ( n40473,n40476,n38200 );
   nor U41392 ( n40453,n40477,n40478 );
   nand U41393 ( n40478,n40479,n40480 );
   nor U41394 ( n40480,n40481,n40482 );
   nor U41395 ( n40482,n40483,n38282 );
   nor U41396 ( n40481,n40484,n38452 );
   nor U41397 ( n40479,n40485,n40486 );
   nor U41398 ( n40486,n40487,n38543 );
   nor U41399 ( n40485,n38572,n38692 );
   nand U41400 ( n40477,n40488,n40489 );
   nor U41401 ( n40489,n40490,n40491 );
   nor U41402 ( n40491,n40492,n37328 );
   nor U41403 ( n40490,n40493,n37686 );
   nor U41404 ( n40488,n40494,n40495 );
   nor U41405 ( n40495,n40496,n38019 );
   nor U41406 ( n40494,n40497,n38366 );
   or U41407 ( n40413,n40419,n40418 );
   and U41408 ( n40418,n40498,n40499 );
   nand U41409 ( n40499,n39545,n40500 );
   nand U41410 ( n40498,n40501,n28280 );
   nand U41411 ( n40501,n40502,n40503 );
   nor U41412 ( n40503,n40504,n40505 );
   nand U41413 ( n40505,n40506,n40507 );
   nor U41414 ( n40507,n40508,n40509 );
   nor U41415 ( n40509,n40510,n37423 );
   nor U41416 ( n40508,n40511,n37511 );
   nor U41417 ( n40506,n40512,n40513 );
   nor U41418 ( n40513,n40514,n37597 );
   nor U41419 ( n40512,n40515,n37774 );
   nand U41420 ( n40504,n40516,n40517 );
   nor U41421 ( n40517,n40518,n40519 );
   nor U41422 ( n40519,n40520,n37857 );
   nor U41423 ( n40518,n40521,n37941 );
   nor U41424 ( n40516,n40522,n40523 );
   nor U41425 ( n40523,n40524,n38111 );
   nor U41426 ( n40522,n40525,n38200 );
   nor U41427 ( n40502,n40526,n40527 );
   nand U41428 ( n40527,n40528,n40529 );
   nor U41429 ( n40529,n40530,n40531 );
   nor U41430 ( n40531,n40532,n38282 );
   nor U41431 ( n40530,n40533,n38452 );
   nor U41432 ( n40528,n40534,n40535 );
   nor U41433 ( n40535,n40536,n38543 );
   nor U41434 ( n40534,n38590,n38692 );
   nand U41435 ( n40526,n40537,n40538 );
   nor U41436 ( n40538,n40539,n40540 );
   nor U41437 ( n40540,n40541,n37328 );
   nor U41438 ( n40539,n40542,n37686 );
   nor U41439 ( n40537,n40543,n40544 );
   nor U41440 ( n40544,n40545,n38019 );
   nor U41441 ( n40543,n40546,n38366 );
   nand U41442 ( n40419,n40547,n40428 );
   nor U41443 ( n40428,n40449,n40448 );
   and U41444 ( n40448,n40548,n40549 );
   nand U41445 ( n40549,n39545,n40550 );
   nand U41446 ( n40548,n40551,n28280 );
   nand U41447 ( n40551,n40552,n40553 );
   nor U41448 ( n40553,n40554,n40555 );
   nand U41449 ( n40555,n40556,n40557 );
   nor U41450 ( n40557,n40558,n40559 );
   nor U41451 ( n40559,n40560,n37328 );
   nor U41452 ( n40558,n40561,n37686 );
   nor U41453 ( n40556,n40562,n40563 );
   nor U41454 ( n40563,n40564,n38019 );
   nor U41455 ( n40562,n40565,n38366 );
   nand U41456 ( n40554,n40566,n40567 );
   nor U41457 ( n40567,n40568,n40569 );
   nor U41458 ( n40569,n40570,n38282 );
   nor U41459 ( n40568,n40571,n38452 );
   nor U41460 ( n40566,n40572,n40573 );
   nor U41461 ( n40573,n40574,n38543 );
   nor U41462 ( n40572,n38638,n38692 );
   nor U41463 ( n40552,n40575,n40576 );
   nand U41464 ( n40576,n40577,n40578 );
   nor U41465 ( n40578,n40579,n40580 );
   nor U41466 ( n40580,n40581,n37857 );
   nor U41467 ( n40579,n40582,n37941 );
   nor U41468 ( n40577,n40583,n40584 );
   nor U41469 ( n40584,n40585,n38111 );
   nor U41470 ( n40583,n40586,n38200 );
   nand U41471 ( n40575,n40587,n40588 );
   nor U41472 ( n40588,n40589,n40590 );
   nor U41473 ( n40590,n40591,n37423 );
   nor U41474 ( n40589,n40592,n37511 );
   nor U41475 ( n40587,n40593,n40594 );
   nor U41476 ( n40594,n40595,n37597 );
   nor U41477 ( n40593,n40596,n37774 );
   nand U41478 ( n40449,n40597,n40598 );
   nand U41479 ( n40598,n40599,n28280 );
   nand U41480 ( n40599,n40447,n40445 );
   or U41481 ( n40597,n40445,n40447 );
   and U41482 ( n40447,n40444,n40443 );
   or U41483 ( n40443,n40442,n28280 );
   nand U41484 ( n40442,n40600,n40601 );
   nand U41485 ( n40601,n27896,n40602 );
   nand U41486 ( n40600,n40603,n28280 );
   nand U41487 ( n40603,n40604,n40605 );
   nor U41488 ( n40605,n40606,n40607 );
   nand U41489 ( n40607,n40608,n40609 );
   nor U41490 ( n40609,n40610,n40611 );
   nor U41491 ( n40611,n40612,n37423 );
   nor U41492 ( n40610,n40613,n37511 );
   nor U41493 ( n40608,n40614,n40615 );
   nor U41494 ( n40615,n40616,n37597 );
   nor U41495 ( n40614,n40617,n37774 );
   nand U41496 ( n40606,n40618,n40619 );
   nor U41497 ( n40619,n40620,n40621 );
   nor U41498 ( n40621,n40622,n37857 );
   nor U41499 ( n40620,n40623,n37941 );
   nor U41500 ( n40618,n40624,n40625 );
   nor U41501 ( n40625,n40626,n38111 );
   nor U41502 ( n40624,n40627,n38200 );
   nor U41503 ( n40604,n40628,n40629 );
   nand U41504 ( n40629,n40630,n40631 );
   nor U41505 ( n40631,n40632,n40633 );
   nor U41506 ( n40633,n40634,n38282 );
   nor U41507 ( n40632,n40635,n38452 );
   nor U41508 ( n40630,n40636,n40637 );
   nor U41509 ( n40637,n40638,n38543 );
   nor U41510 ( n40636,n38693,n38692 );
   nand U41511 ( n40628,n40639,n40640 );
   nor U41512 ( n40640,n40641,n40642 );
   nor U41513 ( n40642,n40643,n37328 );
   nor U41514 ( n40641,n40644,n37686 );
   nor U41515 ( n40639,n40645,n40646 );
   nor U41516 ( n40646,n40647,n38019 );
   nor U41517 ( n40645,n40648,n38366 );
   nand U41518 ( n40444,n40649,n40650 );
   nand U41519 ( n40650,n27896,n40651 );
   nand U41520 ( n40649,n40652,n28280 );
   nand U41521 ( n40652,n40653,n40654 );
   nor U41522 ( n40654,n40655,n40656 );
   nand U41523 ( n40656,n40657,n40658 );
   nor U41524 ( n40658,n40659,n40660 );
   nor U41525 ( n40660,n40661,n37423 );
   nor U41526 ( n40659,n40662,n37511 );
   nor U41527 ( n40657,n40663,n40664 );
   nor U41528 ( n40664,n40665,n37597 );
   nor U41529 ( n40663,n40666,n37774 );
   nand U41530 ( n40655,n40667,n40668 );
   nor U41531 ( n40668,n40669,n40670 );
   nor U41532 ( n40670,n40671,n37857 );
   nor U41533 ( n40669,n40672,n37941 );
   nor U41534 ( n40667,n40673,n40674 );
   nor U41535 ( n40674,n40675,n38111 );
   nor U41536 ( n40673,n40676,n38200 );
   nor U41537 ( n40653,n40677,n40678 );
   nand U41538 ( n40678,n40679,n40680 );
   nor U41539 ( n40680,n40681,n40682 );
   nor U41540 ( n40682,n40683,n38282 );
   nor U41541 ( n40681,n40684,n38452 );
   nor U41542 ( n40679,n40685,n40686 );
   nor U41543 ( n40686,n40687,n38543 );
   nor U41544 ( n40685,n38669,n38692 );
   nand U41545 ( n40677,n40688,n40689 );
   nor U41546 ( n40689,n40690,n40691 );
   nor U41547 ( n40691,n40692,n37328 );
   nor U41548 ( n40690,n40693,n37686 );
   nor U41549 ( n40688,n40694,n40695 );
   nor U41550 ( n40695,n40696,n38019 );
   nor U41551 ( n40694,n40697,n38366 );
   nand U41552 ( n40445,n40698,n40699 );
   nand U41553 ( n40699,n27896,n40700 );
   nand U41554 ( n40698,n40701,n28280 );
   nand U41555 ( n40701,n40702,n40703 );
   nor U41556 ( n40703,n40704,n40705 );
   nand U41557 ( n40705,n40706,n40707 );
   nor U41558 ( n40707,n40708,n40709 );
   nor U41559 ( n40709,n40710,n37423 );
   nor U41560 ( n40708,n40711,n37511 );
   nor U41561 ( n40706,n40712,n40713 );
   nor U41562 ( n40713,n40714,n37597 );
   nor U41563 ( n40712,n40715,n37774 );
   nand U41564 ( n40704,n40716,n40717 );
   nor U41565 ( n40717,n40718,n40719 );
   nor U41566 ( n40719,n40720,n37857 );
   nor U41567 ( n40718,n40721,n37941 );
   nor U41568 ( n40716,n40722,n40723 );
   nor U41569 ( n40723,n40724,n38111 );
   nor U41570 ( n40722,n40725,n38200 );
   nor U41571 ( n40702,n40726,n40727 );
   nand U41572 ( n40727,n40728,n40729 );
   nor U41573 ( n40729,n40730,n40731 );
   nor U41574 ( n40731,n40732,n38282 );
   nor U41575 ( n40730,n40733,n38452 );
   nor U41576 ( n40728,n40734,n40735 );
   nor U41577 ( n40735,n40736,n38543 );
   nor U41578 ( n40734,n38654,n38692 );
   nand U41579 ( n40726,n40737,n40738 );
   nor U41580 ( n40738,n40739,n40740 );
   nor U41581 ( n40740,n40741,n37328 );
   nor U41582 ( n40739,n40742,n37686 );
   nor U41583 ( n40737,n40743,n40744 );
   nor U41584 ( n40744,n40745,n38019 );
   nor U41585 ( n40743,n40746,n38366 );
   nor U41586 ( n40547,n40450,n40426 );
   and U41587 ( n40426,n40747,n40748 );
   nand U41588 ( n40748,n39545,n40749 );
   nand U41589 ( n40747,n40750,n28280 );
   nand U41590 ( n40750,n40751,n40752 );
   nor U41591 ( n40752,n40753,n40754 );
   nand U41592 ( n40754,n40755,n40756 );
   nor U41593 ( n40756,n40757,n40758 );
   nor U41594 ( n40758,n40759,n37328 );
   nor U41595 ( n40757,n40760,n37686 );
   nor U41596 ( n40755,n40761,n40762 );
   nor U41597 ( n40762,n40763,n38019 );
   nor U41598 ( n40761,n40764,n38366 );
   nand U41599 ( n40753,n40765,n40766 );
   nor U41600 ( n40766,n40767,n40768 );
   nor U41601 ( n40768,n40769,n38282 );
   nor U41602 ( n40767,n40770,n38452 );
   nor U41603 ( n40765,n40771,n40772 );
   nor U41604 ( n40772,n40773,n38543 );
   nor U41605 ( n40771,n38606,n38692 );
   nor U41606 ( n40751,n40774,n40775 );
   nand U41607 ( n40775,n40776,n40777 );
   nor U41608 ( n40777,n40778,n40779 );
   nor U41609 ( n40779,n40780,n37857 );
   nor U41610 ( n40778,n40781,n37941 );
   nor U41611 ( n40776,n40782,n40783 );
   nor U41612 ( n40783,n40784,n38111 );
   nor U41613 ( n40782,n40785,n38200 );
   nand U41614 ( n40774,n40786,n40787 );
   nor U41615 ( n40787,n40788,n40789 );
   nor U41616 ( n40789,n40790,n37423 );
   nor U41617 ( n40788,n40791,n37511 );
   nor U41618 ( n40786,n40792,n40793 );
   nor U41619 ( n40793,n40794,n37597 );
   nor U41620 ( n40792,n40795,n37774 );
   not U41621 ( n40450,n40429 );
   nand U41622 ( n40429,n40796,n40797 );
   nand U41623 ( n40797,n39545,n40798 );
   nand U41624 ( n40796,n40799,n28280 );
   nand U41625 ( n40799,n40800,n40801 );
   nor U41626 ( n40801,n40802,n40803 );
   nand U41627 ( n40803,n40804,n40805 );
   nor U41628 ( n40805,n40806,n40807 );
   nor U41629 ( n40807,n40808,n37423 );
   nand U41630 ( n37423,n40809,n40810 );
   nor U41631 ( n40806,n40811,n37511 );
   nand U41632 ( n37511,n40812,n40813 );
   nor U41633 ( n40804,n40814,n40815 );
   nor U41634 ( n40815,n40816,n37597 );
   nand U41635 ( n37597,n40812,n40809 );
   nor U41636 ( n40814,n40817,n37774 );
   nand U41637 ( n37774,n40818,n40810 );
   nand U41638 ( n40802,n40819,n40820 );
   nor U41639 ( n40820,n40821,n40822 );
   nor U41640 ( n40822,n40823,n37857 );
   nand U41641 ( n37857,n40824,n40812 );
   nor U41642 ( n40821,n40825,n37941 );
   nand U41643 ( n37941,n40818,n40812 );
   nor U41644 ( n40812,n38745,n37159 );
   nor U41645 ( n40819,n40826,n40827 );
   nor U41646 ( n40827,n40828,n38111 );
   nand U41647 ( n38111,n40829,n40809 );
   nor U41648 ( n40826,n40830,n38200 );
   nand U41649 ( n38200,n40831,n40813 );
   nor U41650 ( n40800,n40832,n40833 );
   nand U41651 ( n40833,n40834,n40835 );
   nor U41652 ( n40835,n40836,n40837 );
   nor U41653 ( n40837,n40838,n38282 );
   nand U41654 ( n38282,n40831,n40809 );
   nor U41655 ( n40809,n37189,n37116 );
   nor U41656 ( n40836,n40839,n38452 );
   nand U41657 ( n38452,n40829,n40818 );
   nor U41658 ( n40834,n40840,n40841 );
   nor U41659 ( n40841,n40842,n38543 );
   nand U41660 ( n38543,n40831,n40824 );
   nor U41661 ( n40840,n38622,n38692 );
   nand U41662 ( n38692,n40831,n40818 );
   nor U41663 ( n40818,n38766,n37116 );
   nor U41664 ( n40831,n40843,n38745 );
   nand U41665 ( n40832,n40844,n40845 );
   nor U41666 ( n40845,n40846,n40847 );
   nor U41667 ( n40847,n40848,n37328 );
   nand U41668 ( n37328,n40813,n40810 );
   nor U41669 ( n40846,n40849,n37686 );
   nand U41670 ( n37686,n40824,n40810 );
   nor U41671 ( n40810,n37159,n37125 );
   nor U41672 ( n40844,n40850,n40851 );
   nor U41673 ( n40851,n40852,n38019 );
   nand U41674 ( n38019,n40829,n40813 );
   nor U41675 ( n40813,n37189,n38726 );
   nor U41676 ( n40850,n40853,n38366 );
   nand U41677 ( n38366,n40829,n40824 );
   nor U41678 ( n40824,n38726,n38766 );
   nor U41679 ( n40829,n40843,n37125 );
   and U41680 ( n40121,n40854,n40855 );
   nor U41681 ( n40855,n40856,n40857 );
   nand U41682 ( n40857,p2_instaddrpointer_reg_23_,n39490 );
   nor U41683 ( n39490,n39261,n39234 );
   nand U41684 ( n40856,n39259,n40122 );
   and U41685 ( n40122,n40858,n40859 );
   nor U41686 ( n40859,n39910,n39118 );
   nand U41687 ( n39910,n40860,n39494 );
   nor U41688 ( n39494,n39070,n39043 );
   nor U41689 ( n40860,n39847,n39092 );
   nand U41690 ( n39847,n40861,p2_instaddrpointer_reg_12_ );
   nor U41691 ( n40861,n39496,n38996 );
   nand U41692 ( n39496,p2_instaddrpointer_reg_10_,p2_instaddrpointer_reg_9_ );
   nor U41693 ( n40858,n39140,n39166 );
   nor U41694 ( n39259,n39212,n39188 );
   nor U41695 ( n40854,n39357,n40862 );
   nand U41696 ( n40862,p2_instaddrpointer_reg_25_,p2_instaddrpointer_reg_24_ );
   nor U41697 ( n39589,n39622,n40863 );
   nor U41698 ( n40205,n40864,n28123 );
   nand U41699 ( n39604,n40865,p2_statebs16_reg );
   nor U41700 ( n40865,n39622,n28178 );
   not U41701 ( n39622,n28381 );
   not U41702 ( n40864,n39461 );
   nor U41703 ( n40203,n40866,n40867 );
   nand U41704 ( n40867,n40868,n40869 );
   nand U41705 ( n40869,p2_phyaddrpointer_reg_31_,n40870 );
   nand U41706 ( n40870,n28382,n40871 );
   nand U41707 ( n40871,n39620,n40872 );
   not U41708 ( n39620,n39595 );
   nand U41709 ( n40868,n40873,n40874 );
   not U41710 ( n40874,p2_phyaddrpointer_reg_31_ );
   nor U41711 ( n40873,n40872,n39595 );
   nand U41712 ( n39595,n39594,n40875 );
   nand U41713 ( n40875,n40876,n40877 );
   nand U41714 ( n40876,p2_state2_reg_1_,n36648 );
   nor U41715 ( n40866,n36813,n39603 );
   nand U41716 ( n39603,n36653,n28381 );
   nand U41717 ( n39594,n40878,n40879 );
   or U41718 ( n40879,n36673,p2_state2_reg_0_ );
   nor U41719 ( n36673,n36628,n36713 );
   nor U41720 ( n36713,p2_state2_reg_1_,p2_state2_reg_3_ );
   nand U41721 ( n40878,n37045,n37196 );
   nand U41722 ( n37196,n39540,n40880 );
   nand U41723 ( n40880,n37219,n37202 );
   nor U41724 ( n37202,n39506,n37132 );
   not U41725 ( n37219,n37201 );
   nand U41726 ( n39540,n39450,n40881 );
   not U41727 ( n40881,n37205 );
   nor U41728 ( n39450,n39506,n37203 );
   nor U41729 ( n36653,p2_state2_reg_2_,p2_state2_reg_1_ );
   nand U41730 ( n40883,p2_lword_reg_15_,n28336 );
   nor U41731 ( n40882,n40885,n40886 );
   nor U41732 ( n40886,n40887,n28106 );
   nor U41733 ( n40885,n40888,n28225 );
   nand U41734 ( n40891,p2_lword_reg_14_,n28336 );
   nor U41735 ( n40890,n40892,n40893 );
   nor U41736 ( n40893,n40894,n28104 );
   nand U41737 ( n40896,p2_lword_reg_13_,n40884 );
   nor U41738 ( n40895,n40897,n40898 );
   nor U41739 ( n40898,n40899,n28105 );
   nand U41740 ( n40901,p2_lword_reg_12_,n40884 );
   nor U41741 ( n40900,n40902,n40903 );
   nor U41742 ( n40903,n40904,n28106 );
   nand U41743 ( n40906,p2_lword_reg_11_,n40884 );
   nor U41744 ( n40905,n40907,n40908 );
   nor U41745 ( n40908,n40909,n28104 );
   nand U41746 ( n40911,p2_lword_reg_10_,n40884 );
   nor U41747 ( n40910,n40912,n40913 );
   nor U41748 ( n40913,n40914,n28105 );
   nand U41749 ( n40916,p2_lword_reg_9_,n40884 );
   nor U41750 ( n40915,n40917,n40918 );
   nor U41751 ( n40918,n40919,n28106 );
   nand U41752 ( n40921,p2_lword_reg_8_,n40884 );
   nor U41753 ( n40920,n40922,n40923 );
   nor U41754 ( n40923,n40924,n28104 );
   nand U41755 ( n40926,p2_lword_reg_7_,n40884 );
   nor U41756 ( n40925,n40927,n40928 );
   nor U41757 ( n40928,n40929,n28105 );
   nand U41758 ( n40931,p2_lword_reg_6_,n40884 );
   nor U41759 ( n40930,n40932,n40933 );
   nor U41760 ( n40933,n40934,n28106 );
   nand U41761 ( n40936,p2_lword_reg_5_,n40884 );
   nor U41762 ( n40935,n40937,n40938 );
   nor U41763 ( n40938,n40939,n28104 );
   nand U41764 ( n40941,p2_lword_reg_4_,n40884 );
   nor U41765 ( n40940,n40942,n40943 );
   nor U41766 ( n40943,n40944,n28105 );
   nand U41767 ( n40946,p2_lword_reg_3_,n40884 );
   nor U41768 ( n40945,n40947,n40948 );
   nor U41769 ( n40948,n40949,n28106 );
   nand U41770 ( n40951,p2_lword_reg_2_,n40884 );
   nor U41771 ( n40950,n40952,n40953 );
   nor U41772 ( n40953,n40954,n28104 );
   nand U41773 ( n40956,p2_lword_reg_1_,n40884 );
   nor U41774 ( n40955,n40957,n40958 );
   nor U41775 ( n40958,n40959,n28105 );
   nand U41776 ( n40961,p2_lword_reg_0_,n40884 );
   nor U41777 ( n40960,n40962,n40963 );
   nor U41778 ( n40963,n40964,n28106 );
   nand U41779 ( n40966,p2_uword_reg_14_,n40884 );
   nor U41780 ( n40965,n40892,n40967 );
   nor U41781 ( n40967,n40968,n28104 );
   nor U41782 ( n40892,n40889,n40969 );
   nand U41783 ( n40971,p2_uword_reg_13_,n40884 );
   nor U41784 ( n40970,n40897,n40972 );
   nor U41785 ( n40972,n40973,n28105 );
   nor U41786 ( n40897,n40889,n40974 );
   nand U41787 ( n40976,p2_uword_reg_12_,n40884 );
   nor U41788 ( n40975,n40902,n40977 );
   nor U41789 ( n40977,n40978,n28106 );
   nor U41790 ( n40902,n40889,n40979 );
   nand U41791 ( n40981,p2_uword_reg_11_,n40884 );
   nor U41792 ( n40980,n40907,n40982 );
   nor U41793 ( n40982,n40983,n28104 );
   nor U41794 ( n40907,n40889,n40984 );
   nand U41795 ( n40986,p2_uword_reg_10_,n40884 );
   nor U41796 ( n40985,n40912,n40987 );
   nor U41797 ( n40987,n40988,n28105 );
   nor U41798 ( n40912,n40889,n40989 );
   nand U41799 ( n40991,p2_uword_reg_9_,n28336 );
   nor U41800 ( n40990,n40917,n40992 );
   nor U41801 ( n40992,n40993,n28106 );
   nor U41802 ( n40917,n40889,n40994 );
   nand U41803 ( n40996,p2_uword_reg_8_,n28336 );
   nor U41804 ( n40995,n40922,n40997 );
   nor U41805 ( n40997,n40998,n28104 );
   nor U41806 ( n40922,n40889,n40999 );
   nand U41807 ( n41001,p2_uword_reg_7_,n28336 );
   nor U41808 ( n41000,n40927,n41002 );
   nor U41809 ( n41002,n41003,n28105 );
   nor U41810 ( n40927,n38575,n28225 );
   nand U41811 ( n41005,p2_uword_reg_6_,n28336 );
   nor U41812 ( n41004,n40932,n41006 );
   nor U41813 ( n41006,n41007,n28106 );
   nor U41814 ( n40932,n38592,n28225 );
   nand U41815 ( n41009,p2_uword_reg_5_,n28336 );
   nor U41816 ( n41008,n40937,n41010 );
   nor U41817 ( n41010,n41011,n28104 );
   nor U41818 ( n40937,n38608,n40889 );
   nand U41819 ( n41013,p2_uword_reg_4_,n28336 );
   nor U41820 ( n41012,n40942,n41014 );
   nor U41821 ( n41014,n41015,n28105 );
   nor U41822 ( n40942,n38624,n40889 );
   nand U41823 ( n41017,p2_uword_reg_3_,n28336 );
   nor U41824 ( n41016,n40947,n41018 );
   nor U41825 ( n41018,n41019,n28106 );
   nor U41826 ( n40947,n38640,n40889 );
   nand U41827 ( n41021,p2_uword_reg_2_,n28336 );
   nor U41828 ( n41020,n40952,n41022 );
   nor U41829 ( n41022,n41023,n28104 );
   nor U41830 ( n40952,n38656,n28225 );
   nand U41831 ( n41025,p2_uword_reg_1_,n28336 );
   nor U41832 ( n41024,n40957,n41026 );
   nor U41833 ( n41026,n41027,n28105 );
   nor U41834 ( n40957,n38671,n28225 );
   nand U41835 ( n41029,p2_uword_reg_0_,n28336 );
   nor U41836 ( n41028,n40962,n41030 );
   nor U41837 ( n41030,n41031,n28105 );
   nor U41838 ( n40962,n38688,n28225 );
   nand U41839 ( n40889,n41032,n28280 );
   not U41840 ( n41032,n40884 );
   nand U41841 ( n40884,n41033,n41034 );
   nor U41842 ( n41034,n41035,n41036 );
   nor U41843 ( n41035,n39545,n36635 );
   nor U41844 ( n41033,n41037,n39549 );
   nand U41845 ( n41039,n28357,p2_datao_reg_0_ );
   nor U41846 ( n41038,n41041,n41042 );
   nor U41847 ( n41042,n41043,n28101 );
   not U41848 ( n41043,p2_lword_reg_0_ );
   nor U41849 ( n41041,n40964,n41045 );
   nand U41850 ( n41047,n41040,p2_datao_reg_1_ );
   nor U41851 ( n41046,n41048,n41049 );
   nor U41852 ( n41049,n41050,n28101 );
   not U41853 ( n41050,p2_lword_reg_1_ );
   nor U41854 ( n41048,n40959,n28255 );
   nand U41855 ( n41052,n41040,p2_datao_reg_2_ );
   nor U41856 ( n41051,n41053,n41054 );
   nor U41857 ( n41054,n41055,n28100 );
   not U41858 ( n41055,p2_lword_reg_2_ );
   nor U41859 ( n41053,n40954,n28255 );
   nand U41860 ( n41057,n41040,p2_datao_reg_3_ );
   nor U41861 ( n41056,n41058,n41059 );
   nor U41862 ( n41059,n41060,n28101 );
   not U41863 ( n41060,p2_lword_reg_3_ );
   nor U41864 ( n41058,n40949,n28255 );
   nand U41865 ( n41062,n41040,p2_datao_reg_4_ );
   nor U41866 ( n41061,n41063,n41064 );
   nor U41867 ( n41064,n41065,n41044 );
   not U41868 ( n41065,p2_lword_reg_4_ );
   nor U41869 ( n41063,n40944,n41045 );
   nand U41870 ( n41067,n41040,p2_datao_reg_5_ );
   nor U41871 ( n41066,n41068,n41069 );
   nor U41872 ( n41069,n41070,n28100 );
   not U41873 ( n41070,p2_lword_reg_5_ );
   nor U41874 ( n41068,n40939,n41045 );
   nand U41875 ( n41072,n41040,p2_datao_reg_6_ );
   nor U41876 ( n41071,n41073,n41074 );
   nor U41877 ( n41074,n41075,n28101 );
   not U41878 ( n41075,p2_lword_reg_6_ );
   nor U41879 ( n41073,n40934,n41045 );
   nand U41880 ( n41077,n41040,p2_datao_reg_7_ );
   nor U41881 ( n41076,n41078,n41079 );
   nor U41882 ( n41079,n41080,n41044 );
   not U41883 ( n41080,p2_lword_reg_7_ );
   nor U41884 ( n41078,n40929,n41045 );
   nand U41885 ( n41082,n41040,p2_datao_reg_8_ );
   nor U41886 ( n41081,n41083,n41084 );
   nor U41887 ( n41084,n41085,n28100 );
   not U41888 ( n41085,p2_lword_reg_8_ );
   nor U41889 ( n41083,n40924,n41045 );
   nand U41890 ( n41087,n41040,p2_datao_reg_9_ );
   nor U41891 ( n41086,n41088,n41089 );
   nor U41892 ( n41089,n41090,n28101 );
   not U41893 ( n41090,p2_lword_reg_9_ );
   nor U41894 ( n41088,n40919,n41045 );
   nand U41895 ( n41092,n41040,p2_datao_reg_10_ );
   nor U41896 ( n41091,n41093,n41094 );
   nor U41897 ( n41094,n41095,n41044 );
   not U41898 ( n41095,p2_lword_reg_10_ );
   nor U41899 ( n41093,n40914,n41045 );
   nand U41900 ( n41097,n41040,p2_datao_reg_11_ );
   nor U41901 ( n41096,n41098,n41099 );
   nor U41902 ( n41099,n41100,n28100 );
   not U41903 ( n41100,p2_lword_reg_11_ );
   nor U41904 ( n41098,n40909,n41045 );
   nand U41905 ( n41102,n41040,p2_datao_reg_12_ );
   nor U41906 ( n41101,n41103,n41104 );
   nor U41907 ( n41104,n41105,n28101 );
   not U41908 ( n41105,p2_lword_reg_12_ );
   nor U41909 ( n41103,n40904,n41045 );
   nand U41910 ( n41107,n41040,p2_datao_reg_13_ );
   nor U41911 ( n41106,n41108,n41109 );
   nor U41912 ( n41109,n41110,n41044 );
   not U41913 ( n41110,p2_lword_reg_13_ );
   nor U41914 ( n41108,n40899,n41045 );
   nand U41915 ( n41112,n41040,p2_datao_reg_14_ );
   nor U41916 ( n41111,n41113,n41114 );
   nor U41917 ( n41114,n41115,n28100 );
   not U41918 ( n41115,p2_lword_reg_14_ );
   nor U41919 ( n41113,n40894,n28255 );
   nand U41920 ( n41117,n41040,p2_datao_reg_15_ );
   nor U41921 ( n41116,n41118,n41119 );
   nor U41922 ( n41119,n41120,n28101 );
   not U41923 ( n41120,p2_lword_reg_15_ );
   nor U41924 ( n41118,n40887,n41045 );
   nand U41925 ( n41045,p2_state2_reg_0_,n41121 );
   nand U41926 ( n41123,n41040,p2_datao_reg_16_ );
   nor U41927 ( n41122,n41124,n41125 );
   nor U41928 ( n41125,n41031,n41126 );
   nor U41929 ( n41124,n41127,n41044 );
   not U41930 ( n41127,p2_uword_reg_0_ );
   nand U41931 ( n41129,n28357,p2_datao_reg_17_ );
   nor U41932 ( n41128,n41130,n41131 );
   nor U41933 ( n41131,n41027,n27880 );
   nor U41934 ( n41130,n41132,n28100 );
   not U41935 ( n41132,p2_uword_reg_1_ );
   nand U41936 ( n41134,n28357,p2_datao_reg_18_ );
   nor U41937 ( n41133,n41135,n41136 );
   nor U41938 ( n41136,n41023,n27880 );
   nor U41939 ( n41135,n41137,n28101 );
   not U41940 ( n41137,p2_uword_reg_2_ );
   nand U41941 ( n41139,n28357,p2_datao_reg_19_ );
   nor U41942 ( n41138,n41140,n41141 );
   nor U41943 ( n41141,n41019,n27880 );
   nor U41944 ( n41140,n41142,n41044 );
   not U41945 ( n41142,p2_uword_reg_3_ );
   nand U41946 ( n41144,n28357,p2_datao_reg_20_ );
   nor U41947 ( n41143,n41145,n41146 );
   nor U41948 ( n41146,n41015,n41126 );
   nor U41949 ( n41145,n41147,n28100 );
   not U41950 ( n41147,p2_uword_reg_4_ );
   nand U41951 ( n41149,n28357,p2_datao_reg_21_ );
   nor U41952 ( n41148,n41150,n41151 );
   nor U41953 ( n41151,n41011,n41126 );
   nor U41954 ( n41150,n41152,n28101 );
   not U41955 ( n41152,p2_uword_reg_5_ );
   nand U41956 ( n41154,n28357,p2_datao_reg_22_ );
   nor U41957 ( n41153,n41155,n41156 );
   nor U41958 ( n41156,n41007,n41126 );
   nor U41959 ( n41155,n41157,n41044 );
   not U41960 ( n41157,p2_uword_reg_6_ );
   nand U41961 ( n41159,n28357,p2_datao_reg_23_ );
   nor U41962 ( n41158,n41160,n41161 );
   nor U41963 ( n41161,n41003,n41126 );
   nor U41964 ( n41160,n41162,n28100 );
   not U41965 ( n41162,p2_uword_reg_7_ );
   nand U41966 ( n41164,n28357,p2_datao_reg_24_ );
   nor U41967 ( n41163,n41165,n41166 );
   nor U41968 ( n41166,n40998,n41126 );
   nor U41969 ( n41165,n41167,n28101 );
   not U41970 ( n41167,p2_uword_reg_8_ );
   nand U41971 ( n41169,n28357,p2_datao_reg_25_ );
   nor U41972 ( n41168,n41170,n41171 );
   nor U41973 ( n41171,n40993,n41126 );
   nor U41974 ( n41170,n41172,n41044 );
   not U41975 ( n41172,p2_uword_reg_9_ );
   nand U41976 ( n41174,n28357,p2_datao_reg_26_ );
   nor U41977 ( n41173,n41175,n41176 );
   nor U41978 ( n41176,n40988,n41126 );
   nor U41979 ( n41175,n41177,n28100 );
   not U41980 ( n41177,p2_uword_reg_10_ );
   nand U41981 ( n41179,n28357,p2_datao_reg_27_ );
   nor U41982 ( n41178,n41180,n41181 );
   nor U41983 ( n41181,n40983,n41126 );
   nor U41984 ( n41180,n41182,n28101 );
   not U41985 ( n41182,p2_uword_reg_11_ );
   nand U41986 ( n41184,n28357,p2_datao_reg_28_ );
   nor U41987 ( n41183,n41185,n41186 );
   nor U41988 ( n41186,n40978,n41126 );
   nor U41989 ( n41185,n41187,n41044 );
   not U41990 ( n41187,p2_uword_reg_12_ );
   nand U41991 ( n41189,n28357,p2_datao_reg_29_ );
   nor U41992 ( n41188,n41190,n41191 );
   nor U41993 ( n41191,n40973,n41126 );
   nor U41994 ( n41190,n41192,n28100 );
   not U41995 ( n41192,p2_uword_reg_13_ );
   nand U41996 ( n41194,n28357,p2_datao_reg_30_ );
   not U41997 ( n41040,n41121 );
   nor U41998 ( n41193,n41195,n41196 );
   nor U41999 ( n41196,n40968,n41126 );
   nand U42000 ( n41126,n36644,n41121 );
   nor U42001 ( n41195,n41197,n28100 );
   nand U42002 ( n41044,n36783,n41121 );
   not U42003 ( n41197,p2_uword_reg_14_ );
   nand U42004 ( n41121,n41198,n41199 );
   nand U42005 ( n41199,p2_state2_reg_1_,n36634 );
   nor U42006 ( n41198,n41200,n41201 );
   nor U42007 ( n41201,n41202,n41203 );
   or U42008 ( n41203,n39543,n41036 );
   nand U42009 ( n39543,n41204,n36654 );
   nor U42010 ( n41204,n39545,n37168 );
   nor U42011 ( n41200,n41205,n41206 );
   nand U42012 ( n41206,n39556,n39557 );
   not U42013 ( n39556,n39549 );
   nand U42014 ( n41205,n36654,n37045 );
   not U42015 ( n36654,n36647 );
   not U42016 ( n28737,p2_datao_reg_31_ );
   nor U42017 ( n41208,n41209,n41210 );
   nor U42018 ( n41210,n36670,n41211 );
   nand U42019 ( n41211,n41212,n36729 );
   nor U42020 ( n41209,n41213,n41214 );
   not U42021 ( n41214,n36670 );
   nor U42022 ( n41213,n41215,n41216 );
   nor U42023 ( n41215,n36729,n41217 );
   nor U42024 ( n41207,n41218,n41219 );
   nor U42025 ( n41219,n28373,n40964 );
   nor U42026 ( n41218,n38688,n41221 );
   nor U42027 ( n41223,n41224,n41225 );
   nor U42028 ( n41225,n38671,n28256 );
   nor U42029 ( n41224,n41217,n41226 );
   xor U42030 ( n41226,n41227,n41228 );
   xor U42031 ( n41227,n36684,n41229 );
   nor U42032 ( n41222,n41230,n41231 );
   nor U42033 ( n41231,n28372,n40959 );
   not U42034 ( n40959,p2_eax_reg_1_ );
   nor U42035 ( n41230,n41228,n41232 );
   nor U42036 ( n41234,n41235,n41236 );
   nor U42037 ( n41236,n38656,n28256 );
   nor U42038 ( n41235,n41217,n41237 );
   xor U42039 ( n41237,n41238,n41239 );
   xor U42040 ( n41239,n41240,n36697 );
   nor U42041 ( n41233,n41241,n41242 );
   nor U42042 ( n41242,n28373,n40954 );
   nor U42043 ( n41241,n41238,n41232 );
   nor U42044 ( n41244,n41245,n41246 );
   nor U42045 ( n41246,n38640,n28256 );
   nor U42046 ( n41245,n41217,n41247 );
   xor U42047 ( n41247,n41248,n38795 );
   xor U42048 ( n41248,n41249,n36711 );
   nor U42049 ( n41243,n41250,n41251 );
   nor U42050 ( n41251,n28372,n40949 );
   nor U42051 ( n41250,n38795,n41232 );
   nor U42052 ( n41253,n41254,n41255 );
   nor U42053 ( n41255,n38624,n41221 );
   nor U42054 ( n41254,n41217,n41256 );
   xor U42055 ( n41256,n41257,n41258 );
   nand U42056 ( n41258,n41259,n41260 );
   nor U42057 ( n41252,n41261,n41262 );
   nor U42058 ( n41262,n41220,n40944 );
   nor U42059 ( n41261,n41257,n41232 );
   nor U42060 ( n41264,n41265,n41266 );
   nor U42061 ( n41266,n38839,n41267 );
   nand U42062 ( n41267,n41268,n41212 );
   nor U42063 ( n41265,n41269,n41270 );
   nor U42064 ( n41269,n41271,n41216 );
   nor U42065 ( n41271,n41268,n41217 );
   nor U42066 ( n41263,n41272,n41273 );
   nor U42067 ( n41273,n28372,n40939 );
   nor U42068 ( n41272,n38608,n41221 );
   nor U42069 ( n41275,n41276,n41277 );
   nor U42070 ( n41277,n38858,n41278 );
   nand U42071 ( n41278,n41279,n41212 );
   nor U42072 ( n41276,n41280,n41281 );
   nor U42073 ( n41280,n41282,n41216 );
   nor U42074 ( n41282,n41279,n41217 );
   nor U42075 ( n41274,n41283,n41284 );
   nor U42076 ( n41284,n41220,n40934 );
   nor U42077 ( n41283,n38592,n41221 );
   nor U42078 ( n41286,n41287,n41288 );
   nor U42079 ( n41288,n41289,n41217 );
   nor U42080 ( n41287,n38575,n41221 );
   nor U42081 ( n41285,n41290,n41291 );
   nor U42082 ( n41291,n41220,n40929 );
   nor U42083 ( n41290,n41292,n41232 );
   nand U42084 ( n41294,p2_eax_reg_8_,n41295 );
   nor U42085 ( n41293,n41296,n41297 );
   nor U42086 ( n41297,n40999,n41221 );
   nor U42087 ( n41296,n41298,n41299 );
   nand U42088 ( n41301,p2_eax_reg_9_,n41295 );
   nor U42089 ( n41300,n41302,n41303 );
   nor U42090 ( n41303,n40994,n41221 );
   nor U42091 ( n41302,n41298,n38938 );
   nand U42092 ( n41305,p2_eax_reg_10_,n41295 );
   nor U42093 ( n41304,n41306,n41307 );
   nor U42094 ( n41307,n40989,n41221 );
   nor U42095 ( n41306,n41298,n38957 );
   nand U42096 ( n41309,p2_eax_reg_11_,n41295 );
   nor U42097 ( n41308,n41310,n41311 );
   nor U42098 ( n41311,n40984,n41221 );
   nor U42099 ( n41310,n41298,n38986 );
   nand U42100 ( n41313,p2_eax_reg_12_,n41295 );
   nor U42101 ( n41312,n41314,n41315 );
   nor U42102 ( n41315,n40979,n41221 );
   nor U42103 ( n41314,n41298,n41316 );
   nand U42104 ( n41318,p2_eax_reg_13_,n41295 );
   nor U42105 ( n41317,n41319,n41320 );
   nor U42106 ( n41320,n40974,n41221 );
   nor U42107 ( n41319,n41298,n41321 );
   nand U42108 ( n41323,p2_eax_reg_14_,n41295 );
   nor U42109 ( n41322,n41324,n41325 );
   nor U42110 ( n41325,n40969,n28256 );
   nor U42111 ( n41324,n41298,n41326 );
   nand U42112 ( n41328,p2_eax_reg_15_,n41295 );
   nor U42113 ( n41327,n41329,n41330 );
   nor U42114 ( n41330,n41298,n41331 );
   nor U42115 ( n41298,n41216,n41212 );
   nor U42116 ( n41329,n40888,n41221 );
   nand U42117 ( n41221,n41332,n28373 );
   and U42118 ( n40888,n41333,n41334 );
   nand U42119 ( n41334,buf2_reg_15_,n28188 );
   nand U42120 ( n41333,buf1_reg_15_,n27891 );
   nor U42121 ( n41336,n41337,n41338 );
   nand U42122 ( n41338,n41339,n41340 );
   nand U42123 ( n41340,n41341,n41342 );
   not U42124 ( n41342,n38688 );
   nand U42125 ( n38688,n41343,n41344 );
   nand U42126 ( n41344,n27891,n28550 );
   not U42127 ( n28550,buf1_reg_0_ );
   nand U42128 ( n41343,n28188,n30737 );
   not U42129 ( n30737,buf2_reg_0_ );
   nand U42130 ( n41339,n41345,n41212 );
   nor U42131 ( n41337,n28647,n41346 );
   nor U42132 ( n41335,n41347,n41348 );
   nand U42133 ( n41348,n41349,n41350 );
   nand U42134 ( n41350,n41351,buf2_reg_16_ );
   nand U42135 ( n41349,n28259,n39100 );
   nor U42136 ( n41347,n28373,n41031 );
   not U42137 ( n41031,p2_eax_reg_16_ );
   nor U42138 ( n41353,n41354,n41355 );
   nand U42139 ( n41355,n41356,n41357 );
   nand U42140 ( n41357,n41212,n41358 );
   xor U42141 ( n41358,n41359,n41360 );
   nand U42142 ( n41356,n41341,n41361 );
   not U42143 ( n41361,n38671 );
   nand U42144 ( n38671,n41362,n41363 );
   nand U42145 ( n41363,n27891,n28557 );
   not U42146 ( n28557,buf1_reg_1_ );
   nand U42147 ( n41362,n28739,n30712 );
   not U42148 ( n30712,buf2_reg_1_ );
   nor U42149 ( n41354,n28653,n28237 );
   nor U42150 ( n41352,n41364,n41365 );
   nand U42151 ( n41365,n41366,n41367 );
   nand U42152 ( n41367,n41351,buf2_reg_17_ );
   nand U42153 ( n41366,n41216,n39129 );
   nor U42154 ( n41364,n28372,n41027 );
   not U42155 ( n41027,p2_eax_reg_17_ );
   nor U42156 ( n41369,n41370,n41371 );
   nand U42157 ( n41371,n41372,n41373 );
   nand U42158 ( n41373,n41212,n41374 );
   xor U42159 ( n41374,n41375,n41376 );
   nand U42160 ( n41372,n41341,n41377 );
   not U42161 ( n41377,n38656 );
   nand U42162 ( n38656,n41378,n41379 );
   nand U42163 ( n41379,n27891,n28563 );
   not U42164 ( n28563,buf1_reg_2_ );
   nand U42165 ( n41378,n28188,n30701 );
   not U42166 ( n30701,buf2_reg_2_ );
   nor U42167 ( n41370,n28659,n28237 );
   nor U42168 ( n41368,n41380,n41381 );
   nand U42169 ( n41381,n41382,n41383 );
   nand U42170 ( n41383,n41351,buf2_reg_18_ );
   nand U42171 ( n41382,n41216,n39148 );
   nor U42172 ( n41380,n41220,n41023 );
   not U42173 ( n41023,p2_eax_reg_18_ );
   nor U42174 ( n41385,n41386,n41387 );
   nand U42175 ( n41387,n41388,n41389 );
   nand U42176 ( n41389,n41212,n41390 );
   xor U42177 ( n41390,n41391,n41392 );
   nand U42178 ( n41388,n41341,n41393 );
   not U42179 ( n41393,n38640 );
   nand U42180 ( n38640,n41394,n41395 );
   nand U42181 ( n41395,n27891,n28569 );
   not U42182 ( n28569,buf1_reg_3_ );
   nand U42183 ( n41394,n28739,n30690 );
   not U42184 ( n30690,buf2_reg_3_ );
   nor U42185 ( n41386,n28665,n28237 );
   nor U42186 ( n41384,n41396,n41397 );
   nand U42187 ( n41397,n41398,n41399 );
   nand U42188 ( n41399,n41351,buf2_reg_19_ );
   nand U42189 ( n41398,n28259,n39177 );
   nor U42190 ( n41396,n28373,n41019 );
   not U42191 ( n41019,p2_eax_reg_19_ );
   nor U42192 ( n41401,n41402,n41403 );
   nand U42193 ( n41403,n41404,n41405 );
   nand U42194 ( n41405,n41212,n41406 );
   xor U42195 ( n41406,n41407,n41408 );
   nand U42196 ( n41404,n41341,n41409 );
   not U42197 ( n41409,n38624 );
   nand U42198 ( n38624,n41410,n41411 );
   nand U42199 ( n41411,n27891,n28575 );
   not U42200 ( n28575,buf1_reg_4_ );
   nand U42201 ( n41410,n28188,n30680 );
   not U42202 ( n30680,buf2_reg_4_ );
   nor U42203 ( n41402,n28671,n41346 );
   nor U42204 ( n41400,n41412,n41413 );
   nand U42205 ( n41413,n41414,n41415 );
   nand U42206 ( n41415,n41351,buf2_reg_20_ );
   nand U42207 ( n41414,n41216,n39196 );
   nor U42208 ( n41412,n41220,n41015 );
   not U42209 ( n41015,p2_eax_reg_20_ );
   nor U42210 ( n41417,n41418,n41419 );
   nand U42211 ( n41419,n41420,n41421 );
   nand U42212 ( n41421,n41212,n41422 );
   xor U42213 ( n41422,n41423,n41424 );
   nand U42214 ( n41420,n41341,n41425 );
   not U42215 ( n41425,n38608 );
   nand U42216 ( n38608,n41426,n41427 );
   nand U42217 ( n41427,n27891,n28581 );
   not U42218 ( n28581,buf1_reg_5_ );
   nand U42219 ( n41426,n28739,n30669 );
   not U42220 ( n30669,buf2_reg_5_ );
   nor U42221 ( n41418,n28677,n41346 );
   nor U42222 ( n41416,n41428,n41429 );
   nand U42223 ( n41429,n41430,n41431 );
   nand U42224 ( n41431,n41351,buf2_reg_21_ );
   nand U42225 ( n41430,n41216,n39223 );
   nor U42226 ( n41428,n41220,n41011 );
   not U42227 ( n41011,p2_eax_reg_21_ );
   nor U42228 ( n41433,n41434,n41435 );
   nand U42229 ( n41435,n41436,n41437 );
   nand U42230 ( n41437,n41212,n41438 );
   xor U42231 ( n41438,n41439,n41440 );
   nand U42232 ( n41436,n41341,n41441 );
   not U42233 ( n41441,n38592 );
   nand U42234 ( n38592,n41442,n41443 );
   nand U42235 ( n41443,n27891,n28587 );
   not U42236 ( n28587,buf1_reg_6_ );
   nand U42237 ( n41442,n28188,n30658 );
   not U42238 ( n30658,buf2_reg_6_ );
   nor U42239 ( n41434,n28683,n41346 );
   nor U42240 ( n41432,n41444,n41445 );
   nand U42241 ( n41445,n41446,n41447 );
   nand U42242 ( n41447,n41351,buf2_reg_22_ );
   nand U42243 ( n41446,n41216,n39241 );
   nor U42244 ( n41444,n28372,n41007 );
   not U42245 ( n41007,p2_eax_reg_22_ );
   nor U42246 ( n41449,n41450,n41451 );
   nand U42247 ( n41451,n41452,n41453 );
   nand U42248 ( n41453,n41212,n41454 );
   xor U42249 ( n41454,n41455,n41456 );
   nand U42250 ( n41452,n41341,n41457 );
   not U42251 ( n41457,n38575 );
   nand U42252 ( n38575,n41458,n41459 );
   nand U42253 ( n41459,n27891,n28593 );
   not U42254 ( n28593,buf1_reg_7_ );
   nand U42255 ( n41458,n28739,n30643 );
   not U42256 ( n30643,buf2_reg_7_ );
   nor U42257 ( n41450,n28689,n41346 );
   nor U42258 ( n41448,n41460,n41461 );
   nand U42259 ( n41461,n41462,n41463 );
   nand U42260 ( n41463,n41351,buf2_reg_23_ );
   nand U42261 ( n41462,n28259,n39272 );
   nor U42262 ( n41460,n28373,n41003 );
   not U42263 ( n41003,p2_eax_reg_23_ );
   nor U42264 ( n41465,n41466,n41467 );
   nand U42265 ( n41467,n41468,n41469 );
   nand U42266 ( n41469,n41212,n41470 );
   xor U42267 ( n41470,n41471,n41472 );
   nand U42268 ( n41468,n41341,n41473 );
   not U42269 ( n41473,n40999 );
   nand U42270 ( n40999,n41474,n41475 );
   nand U42271 ( n41475,n27891,n28599 );
   not U42272 ( n28599,buf1_reg_8_ );
   nand U42273 ( n41474,n28739,n33208 );
   not U42274 ( n33208,buf2_reg_8_ );
   nor U42275 ( n41466,n28695,n41346 );
   nor U42276 ( n41464,n41476,n41477 );
   nand U42277 ( n41477,n41478,n41479 );
   nand U42278 ( n41479,n41351,buf2_reg_24_ );
   nand U42279 ( n41478,n28259,n39291 );
   nor U42280 ( n41476,n41220,n40998 );
   not U42281 ( n40998,p2_eax_reg_24_ );
   nor U42282 ( n41481,n41482,n41483 );
   nand U42283 ( n41483,n41484,n41485 );
   nand U42284 ( n41485,n41212,n41486 );
   xor U42285 ( n41486,n41487,n41488 );
   nand U42286 ( n41484,n41341,n41489 );
   not U42287 ( n41489,n40994 );
   nand U42288 ( n40994,n41490,n41491 );
   nand U42289 ( n41491,n27891,n28605 );
   not U42290 ( n28605,buf1_reg_9_ );
   nand U42291 ( n41490,n28739,n33203 );
   not U42292 ( n33203,buf2_reg_9_ );
   nor U42293 ( n41482,n28701,n41346 );
   nor U42294 ( n41480,n41492,n41493 );
   nand U42295 ( n41493,n41494,n41495 );
   nand U42296 ( n41495,n41351,buf2_reg_25_ );
   nand U42297 ( n41494,n28259,n39319 );
   nor U42298 ( n41492,n28372,n40993 );
   not U42299 ( n40993,p2_eax_reg_25_ );
   nor U42300 ( n41497,n41498,n41499 );
   nand U42301 ( n41499,n41500,n41501 );
   nand U42302 ( n41501,n41212,n41502 );
   xor U42303 ( n41502,n41503,n41504 );
   nand U42304 ( n41500,n41341,n41505 );
   not U42305 ( n41505,n40989 );
   nand U42306 ( n40989,n41506,n41507 );
   nand U42307 ( n41507,n27891,n28611 );
   not U42308 ( n28611,buf1_reg_10_ );
   nand U42309 ( n41506,n28739,n33198 );
   not U42310 ( n33198,buf2_reg_10_ );
   nor U42311 ( n41498,n28707,n41346 );
   nor U42312 ( n41496,n41508,n41509 );
   nand U42313 ( n41509,n41510,n41511 );
   nand U42314 ( n41511,n41351,buf2_reg_26_ );
   nand U42315 ( n41510,n41216,n39339 );
   nor U42316 ( n41508,n28373,n40988 );
   not U42317 ( n40988,p2_eax_reg_26_ );
   nor U42318 ( n41513,n41514,n41515 );
   nand U42319 ( n41515,n41516,n41517 );
   nand U42320 ( n41517,n41212,n41518 );
   xor U42321 ( n41518,n41519,n41520 );
   nand U42322 ( n41516,n41341,n41521 );
   not U42323 ( n41521,n40984 );
   nand U42324 ( n40984,n41522,n41523 );
   nand U42325 ( n41523,n27891,n28617 );
   not U42326 ( n28617,buf1_reg_11_ );
   nand U42327 ( n41522,n28739,n33193 );
   not U42328 ( n33193,buf2_reg_11_ );
   nor U42329 ( n41514,n28713,n41346 );
   nor U42330 ( n41512,n41524,n41525 );
   nand U42331 ( n41525,n41526,n41527 );
   nand U42332 ( n41527,n41351,buf2_reg_27_ );
   nand U42333 ( n41526,n41216,n39368 );
   nor U42334 ( n41524,n28372,n40983 );
   not U42335 ( n40983,p2_eax_reg_27_ );
   nor U42336 ( n41529,n41530,n41531 );
   nand U42337 ( n41531,n41532,n41533 );
   nand U42338 ( n41533,n41212,n41534 );
   xor U42339 ( n41534,n41535,n41536 );
   nand U42340 ( n41532,n41341,n41537 );
   not U42341 ( n41537,n40979 );
   nand U42342 ( n40979,n41538,n41539 );
   nand U42343 ( n41539,n27891,n28623 );
   not U42344 ( n28623,buf1_reg_12_ );
   nand U42345 ( n41538,n28739,n33188 );
   not U42346 ( n33188,buf2_reg_12_ );
   nor U42347 ( n41530,n28719,n41346 );
   nor U42348 ( n41528,n41540,n41541 );
   nand U42349 ( n41541,n41542,n41543 );
   nand U42350 ( n41543,n41351,buf2_reg_28_ );
   nand U42351 ( n41542,n41216,n39386 );
   nor U42352 ( n41540,n41220,n40978 );
   not U42353 ( n40978,p2_eax_reg_28_ );
   nor U42354 ( n41545,n41546,n41547 );
   nand U42355 ( n41547,n41548,n41549 );
   nand U42356 ( n41549,n41550,n41212 );
   not U42357 ( n41212,n41217 );
   xor U42358 ( n41550,n41551,n41552 );
   nand U42359 ( n41548,n41341,n41553 );
   not U42360 ( n41553,n40974 );
   nand U42361 ( n40974,n41554,n41555 );
   nand U42362 ( n41555,n27891,n28629 );
   not U42363 ( n28629,buf1_reg_13_ );
   nand U42364 ( n41554,n28188,n33183 );
   not U42365 ( n33183,buf2_reg_13_ );
   nor U42366 ( n41546,n28725,n41346 );
   nor U42367 ( n41544,n41556,n41557 );
   nand U42368 ( n41557,n41558,n41559 );
   nand U42369 ( n41559,n41351,buf2_reg_29_ );
   nand U42370 ( n41558,n41216,n39406 );
   nor U42371 ( n41556,n28373,n40973 );
   not U42372 ( n40973,p2_eax_reg_29_ );
   nor U42373 ( n41561,n41562,n41563 );
   nand U42374 ( n41563,n41564,n41565 );
   or U42375 ( n41565,n41566,n41217 );
   nand U42376 ( n41217,n28372,n41567 );
   xor U42377 ( n41566,n41568,n41569 );
   nand U42378 ( n41569,n41552,n41551 );
   and U42379 ( n41552,n41570,n41571 );
   nand U42380 ( n41571,n41572,n41573 );
   or U42381 ( n41572,n41535,n41536 );
   nand U42382 ( n41570,n41535,n41536 );
   nand U42383 ( n41535,n41574,n41575 );
   nand U42384 ( n41575,n41576,n41577 );
   or U42385 ( n41577,n41519,n41520 );
   nand U42386 ( n41574,n41519,n41520 );
   nand U42387 ( n41519,n41578,n41579 );
   nand U42388 ( n41579,n41580,n41581 );
   or U42389 ( n41580,n41503,n41504 );
   nand U42390 ( n41578,n41503,n41504 );
   nand U42391 ( n41503,n41582,n41583 );
   nand U42392 ( n41583,n41584,n41585 );
   or U42393 ( n41585,n41487,n41488 );
   nand U42394 ( n41582,n41487,n41488 );
   nand U42395 ( n41487,n41586,n41587 );
   nand U42396 ( n41587,n41588,n41589 );
   or U42397 ( n41588,n41471,n41472 );
   nand U42398 ( n41586,n41471,n41472 );
   nand U42399 ( n41471,n41590,n41591 );
   nand U42400 ( n41591,n41592,n41593 );
   nand U42401 ( n41593,n41456,n41455 );
   or U42402 ( n41590,n41455,n41456 );
   and U42403 ( n41456,n41594,n41595 );
   nand U42404 ( n41595,n41596,n41597 );
   or U42405 ( n41596,n41439,n41440 );
   nand U42406 ( n41594,n41439,n41440 );
   not U42407 ( n41440,n41598 );
   nand U42408 ( n41439,n41599,n41600 );
   nand U42409 ( n41600,n41601,n41602 );
   nand U42410 ( n41602,n41424,n41423 );
   or U42411 ( n41599,n41423,n41424 );
   and U42412 ( n41424,n41603,n41604 );
   nand U42413 ( n41604,n41605,n41606 );
   or U42414 ( n41605,n41407,n41408 );
   nand U42415 ( n41603,n41407,n41408 );
   not U42416 ( n41408,n41607 );
   nand U42417 ( n41407,n41608,n41609 );
   nand U42418 ( n41609,n41610,n41611 );
   nand U42419 ( n41611,n41392,n41391 );
   or U42420 ( n41608,n41391,n41392 );
   and U42421 ( n41392,n41612,n41613 );
   nand U42422 ( n41613,n41614,n41615 );
   or U42423 ( n41614,n41375,n41376 );
   nand U42424 ( n41612,n41375,n41376 );
   not U42425 ( n41376,n41616 );
   nand U42426 ( n41375,n41617,n41618 );
   nand U42427 ( n41618,n41619,n41620 );
   or U42428 ( n41620,n41359,n41360 );
   nand U42429 ( n41617,n41360,n41359 );
   nand U42430 ( n41359,n41621,n41622 );
   nand U42431 ( n41622,n41623,n41624 );
   nand U42432 ( n41624,n39080,n41625 );
   nor U42433 ( n41623,n41626,n41627 );
   nor U42434 ( n41627,n41628,n41629 );
   nor U42435 ( n41626,n41630,n41631 );
   nand U42436 ( n41631,n41632,n41633 );
   nand U42437 ( n41633,n41634,n41635 );
   nand U42438 ( n41635,n39052,n41636 );
   nor U42439 ( n41634,n41637,n41638 );
   nor U42440 ( n41638,n41639,n41640 );
   nor U42441 ( n41637,n41641,n41321 );
   and U42442 ( n41641,n41639,n41640 );
   nand U42443 ( n41639,n41642,n41643 );
   nand U42444 ( n41643,n41644,n41645 );
   nand U42445 ( n41645,n41646,n41647 );
   nor U42446 ( n41644,n41648,n41649 );
   nor U42447 ( n41649,n41650,n41316 );
   nor U42448 ( n41648,n41651,n41652 );
   nand U42449 ( n41652,n41653,n41654 );
   nand U42450 ( n41654,n41655,n41656 );
   nand U42451 ( n41656,n41657,n41658 );
   nor U42452 ( n41655,n41659,n41660 );
   and U42453 ( n41660,n41661,n41662 );
   nor U42454 ( n41659,n41663,n38938 );
   nor U42455 ( n41663,n41662,n41661 );
   nand U42456 ( n41661,n41664,n41665 );
   nand U42457 ( n41665,n38907,n41666 );
   or U42458 ( n41666,n41667,n41668 );
   nand U42459 ( n41664,n41668,n41667 );
   nand U42460 ( n41667,n41669,n41670 );
   nand U42461 ( n41670,n41671,n41672 );
   not U42462 ( n41672,n41289 );
   nor U42463 ( n41289,n41673,n38887 );
   nand U42464 ( n41671,n41674,n41675 );
   nand U42465 ( n41675,n38858,n41676 );
   nand U42466 ( n41676,n41677,n41678 );
   nand U42467 ( n41674,n41279,n41679 );
   not U42468 ( n41279,n41678 );
   nand U42469 ( n41678,n41680,n41681 );
   nand U42470 ( n41681,n41682,n41683 );
   nand U42471 ( n41682,n41268,n38839 );
   not U42472 ( n41268,n41684 );
   nand U42473 ( n41680,n41270,n41684 );
   nand U42474 ( n41684,n41685,n41686 );
   nand U42475 ( n41686,n41687,n41260 );
   or U42476 ( n41687,n41259,n41257 );
   nand U42477 ( n41685,n41257,n41259 );
   nand U42478 ( n41259,n41688,n41689 );
   nand U42479 ( n41689,n36711,n41690 );
   or U42480 ( n41690,n41249,n38795 );
   not U42481 ( n36711,n36772 );
   nand U42482 ( n41688,n38795,n41249 );
   nand U42483 ( n41249,n41691,n41692 );
   nand U42484 ( n41692,n41693,n36697 );
   or U42485 ( n41693,n41240,n41238 );
   nand U42486 ( n41691,n41238,n41240 );
   nand U42487 ( n41240,n41694,n41695 );
   nand U42488 ( n41695,n41228,n41696 );
   nand U42489 ( n41696,n37693,n36670 );
   nor U42490 ( n37693,n36684,n36674 );
   not U42491 ( n41228,n36680 );
   nand U42492 ( n41694,n36684,n41229 );
   nand U42493 ( n41229,n36670,n36729 );
   nand U42494 ( n41669,n38887,n41673 );
   or U42495 ( n41653,n41658,n41657 );
   nor U42496 ( n41651,n41646,n41647 );
   nand U42497 ( n41642,n41650,n41316 );
   not U42498 ( n41650,n41697 );
   nand U42499 ( n41632,n41698,n41326 );
   nor U42500 ( n41630,n39080,n41625 );
   nand U42501 ( n41621,n41629,n41628 );
   not U42502 ( n41629,n41345 );
   not U42503 ( n41360,n41699 );
   nand U42504 ( n41564,n41341,n41700 );
   not U42505 ( n41700,n40969 );
   nand U42506 ( n40969,n41701,n41702 );
   nand U42507 ( n41702,n27891,n28635 );
   not U42508 ( n28635,buf1_reg_14_ );
   nand U42509 ( n41701,n28188,n33178 );
   not U42510 ( n33178,buf2_reg_14_ );
   and U42511 ( n41341,n41703,n41220 );
   nor U42512 ( n41703,n39566,n38601 );
   nor U42513 ( n41562,n28731,n28237 );
   nor U42514 ( n41560,n41704,n41705 );
   nand U42515 ( n41705,n41706,n41707 );
   nand U42516 ( n41707,n41351,buf2_reg_30_ );
   nand U42517 ( n41706,n41216,n39432 );
   nor U42518 ( n41704,n28372,n40968 );
   nor U42519 ( n41709,n41710,n41711 );
   and U42520 ( n41711,buf2_reg_31_,n41351 );
   and U42521 ( n41351,n41712,n41713 );
   nor U42522 ( n41713,n28750,n39515 );
   not U42523 ( n28750,n28739 );
   nor U42524 ( n41712,n39566,n41295 );
   nor U42525 ( n41710,n28736,n41346 );
   nand U42526 ( n41346,n41714,n41715 );
   nor U42527 ( n41714,n28739,n41295 );
   nand U42528 ( n28739,p2_address_reg_29_,n41716 );
   nand U42529 ( n41716,n41717,n41718 );
   nor U42530 ( n41718,n41719,n41720 );
   nand U42531 ( n41720,n41721,n41722 );
   nor U42532 ( n41722,n41723,n41724 );
   or U42533 ( n41724,p2_address_reg_25_,p2_address_reg_26_ );
   or U42534 ( n41723,p2_address_reg_27_,p2_address_reg_28_ );
   nor U42535 ( n41721,p2_address_reg_22_,n41725 );
   or U42536 ( n41725,p2_address_reg_23_,p2_address_reg_24_ );
   nand U42537 ( n41719,n41726,n41727 );
   nor U42538 ( n41727,n41728,n41729 );
   or U42539 ( n41729,p2_address_reg_6_,p2_address_reg_7_ );
   or U42540 ( n41728,p2_address_reg_8_,p2_address_reg_9_ );
   nor U42541 ( n41726,n41730,n41731 );
   or U42542 ( n41731,p2_address_reg_2_,p2_address_reg_3_ );
   or U42543 ( n41730,p2_address_reg_4_,p2_address_reg_5_ );
   nor U42544 ( n41717,n41732,n41733 );
   nand U42545 ( n41733,n41734,n41735 );
   nor U42546 ( n41735,n41736,n41737 );
   or U42547 ( n41737,p2_address_reg_12_,p2_address_reg_13_ );
   or U42548 ( n41736,p2_address_reg_14_,p2_address_reg_15_ );
   nor U42549 ( n41734,p2_address_reg_0_,n41738 );
   or U42550 ( n41738,p2_address_reg_10_,p2_address_reg_11_ );
   nand U42551 ( n41732,n41739,n41740 );
   nor U42552 ( n41740,n41741,n41742 );
   or U42553 ( n41742,p2_address_reg_19_,p2_address_reg_1_ );
   or U42554 ( n41741,p2_address_reg_20_,p2_address_reg_21_ );
   nor U42555 ( n41739,p2_address_reg_16_,n41743 );
   or U42556 ( n41743,p2_address_reg_17_,p2_address_reg_18_ );
   nor U42557 ( n41708,n41744,n41745 );
   nor U42558 ( n41745,n28373,n41746 );
   not U42559 ( n41220,n41295 );
   nor U42560 ( n41744,n39451,n41232 );
   not U42561 ( n41232,n41216 );
   nor U42562 ( n41216,n41295,n38565 );
   nand U42563 ( n41295,n37045,n41747 );
   nand U42564 ( n41747,n41748,n41749 );
   nand U42565 ( n41749,n41750,n39467 );
   not U42566 ( n41748,n37172 );
   nand U42567 ( n37172,n41751,n41752 );
   nand U42568 ( n41752,n41753,n37213 );
   nor U42569 ( n41753,n37052,n41754 );
   nor U42570 ( n41754,n41755,n36776 );
   not U42571 ( n36776,n37078 );
   nor U42572 ( n41755,n41756,n37132 );
   nand U42573 ( n41751,n37179,n37166 );
   not U42574 ( n37179,n37212 );
   nand U42575 ( n37212,n41757,n37134 );
   nor U42576 ( n41757,n38649,n37136 );
   not U42577 ( n39451,n41758 );
   nand U42578 ( n41760,n41761,n36729 );
   nor U42579 ( n41759,n41762,n41763 );
   nor U42580 ( n41763,n38726,n28148 );
   nor U42581 ( n41762,n28154,n41766 );
   nand U42582 ( n41768,n41761,n36740 );
   nor U42583 ( n41767,n41769,n41770 );
   nor U42584 ( n41770,n37125,n41764 );
   nor U42585 ( n41769,n28153,n41771 );
   nand U42586 ( n41773,n41761,n36752 );
   nor U42587 ( n41772,n41774,n41775 );
   nor U42588 ( n41775,n28148,n37189 );
   nor U42589 ( n41774,n28152,n41776 );
   nand U42590 ( n41778,n41761,n36772 );
   nor U42591 ( n41777,n41779,n41780 );
   nor U42592 ( n41780,n37159,n28148 );
   nor U42593 ( n41779,n28154,n41781 );
   nand U42594 ( n41783,n41761,n41784 );
   not U42595 ( n41784,n41260 );
   nor U42596 ( n41782,n41785,n41786 );
   nor U42597 ( n41786,n41764,n39674 );
   nor U42598 ( n41785,n28152,n41787 );
   nand U42599 ( n41789,n41790,n28091 );
   nor U42600 ( n41788,n41791,n41792 );
   nor U42601 ( n41792,n28148,n39694 );
   not U42602 ( n39694,n38840 );
   nor U42603 ( n41791,n41765,n41793 );
   nand U42604 ( n41795,n41761,n41679 );
   not U42605 ( n41679,n41677 );
   xor U42606 ( n41677,n41796,n41797 );
   nand U42607 ( n41797,n41798,p2_instqueue_reg_0__6_ );
   nor U42608 ( n41794,n41799,n41800 );
   nor U42609 ( n41800,n39713,n28147 );
   nor U42610 ( n41799,n28153,n41801 );
   nand U42611 ( n41803,n41761,n41673 );
   xor U42612 ( n41673,n41804,n41805 );
   nor U42613 ( n41802,n41806,n41807 );
   nor U42614 ( n41807,n28147,n39733 );
   nor U42615 ( n41806,n28154,n41808 );
   nand U42616 ( n41810,n41761,n41668 );
   xor U42617 ( n41668,n41811,n41812 );
   nor U42618 ( n41809,n41813,n41814 );
   nor U42619 ( n41814,n38908,n28147 );
   nor U42620 ( n41813,n28154,n41815 );
   nand U42621 ( n41817,n41761,n41662 );
   and U42622 ( n41662,n41818,n41819 );
   nand U42623 ( n41819,n41820,n41821 );
   nand U42624 ( n41820,n41812,n41811 );
   not U42625 ( n41811,n41822 );
   nor U42626 ( n41816,n41823,n41824 );
   nor U42627 ( n41824,n28148,n39770 );
   nor U42628 ( n41823,n28152,n41825 );
   nand U42629 ( n41827,n41761,n41658 );
   xor U42630 ( n41658,n41818,n41828 );
   nand U42631 ( n41828,n41798,n41829 );
   nor U42632 ( n41826,n41830,n41831 );
   nor U42633 ( n41831,n39790,n28148 );
   nor U42634 ( n41830,n41765,n41832 );
   nand U42635 ( n41834,n41761,n41647 );
   xor U42636 ( n41647,n41835,n41836 );
   nor U42637 ( n41833,n41837,n41838 );
   nor U42638 ( n41838,n41764,n39809 );
   nor U42639 ( n41837,n28153,n41839 );
   nand U42640 ( n41841,n41761,n41697 );
   xor U42641 ( n41697,n41842,n41843 );
   nor U42642 ( n41840,n41844,n41845 );
   nor U42643 ( n41845,n39831,n28148 );
   nor U42644 ( n41844,n28152,n41846 );
   nand U42645 ( n41848,n41761,n41849 );
   not U42646 ( n41849,n41640 );
   nand U42647 ( n41640,n41850,n41851 );
   nand U42648 ( n41851,n41852,n41853 );
   nand U42649 ( n41852,n41842,n41843 );
   not U42650 ( n41843,n41854 );
   nor U42651 ( n41847,n41855,n41856 );
   nor U42652 ( n41856,n28147,n39034 );
   nor U42653 ( n41855,n41765,n41857 );
   nand U42654 ( n41859,n41761,n41636 );
   not U42655 ( n41636,n41698 );
   xor U42656 ( n41698,n41860,n41850 );
   nor U42657 ( n41860,n41861,n41862 );
   nor U42658 ( n41858,n41863,n41864 );
   nor U42659 ( n41864,n39053,n28148 );
   nor U42660 ( n41863,n28153,n41865 );
   nand U42661 ( n41867,n41761,n41625 );
   xor U42662 ( n41625,n41868,n41869 );
   nand U42663 ( n41869,n41798,n41870 );
   not U42664 ( n41868,n41871 );
   nor U42665 ( n41866,n41872,n41873 );
   nor U42666 ( n41873,n41764,n39894 );
   nor U42667 ( n41872,n28154,n41874 );
   nand U42668 ( n41876,n41761,n41345 );
   nor U42669 ( n41345,n41877,n41878 );
   and U42670 ( n41877,n41879,n41880 );
   nor U42671 ( n41875,n41881,n41882 );
   nor U42672 ( n41882,n39101,n28147 );
   nor U42673 ( n41881,n28152,n41883 );
   nand U42674 ( n41885,n28091,n41699 );
   xor U42675 ( n41699,n41886,n41878 );
   nor U42676 ( n41884,n41887,n41888 );
   nor U42677 ( n41888,n28148,n39130 );
   nor U42678 ( n41887,n41765,n41889 );
   nand U42679 ( n41891,n28091,n41616 );
   nor U42680 ( n41616,n41892,n41893 );
   and U42681 ( n41893,n41894,n41895 );
   nor U42682 ( n41890,n41896,n41897 );
   nor U42683 ( n41897,n39149,n41764 );
   nor U42684 ( n41896,n28153,n41898 );
   nand U42685 ( n41900,n28091,n41391 );
   xor U42686 ( n41391,n41901,n41892 );
   nor U42687 ( n41899,n41902,n41903 );
   nor U42688 ( n41903,n41764,n39178 );
   nor U42689 ( n41902,n28154,n41904 );
   nand U42690 ( n41906,n28091,n41607 );
   nor U42691 ( n41607,n41907,n41908 );
   and U42692 ( n41908,n41909,n41910 );
   nor U42693 ( n41905,n41911,n41912 );
   nor U42694 ( n41912,n39197,n28148 );
   nor U42695 ( n41911,n28152,n41913 );
   nand U42696 ( n41915,n28091,n41423 );
   xor U42697 ( n41423,n41916,n41907 );
   nor U42698 ( n41914,n41917,n41918 );
   nor U42699 ( n41918,n28147,n39224 );
   nor U42700 ( n41917,n41765,n41919 );
   nand U42701 ( n41921,n28091,n41598 );
   nor U42702 ( n41598,n41922,n41923 );
   and U42703 ( n41923,n41924,n41925 );
   nor U42704 ( n41920,n41926,n41927 );
   nor U42705 ( n41927,n40038,n41764 );
   nor U42706 ( n41926,n28153,n41928 );
   nand U42707 ( n41930,n28091,n41455 );
   xor U42708 ( n41455,n41931,n41922 );
   nor U42709 ( n41931,n41932,n41933 );
   not U42710 ( n41933,n41934 );
   nor U42711 ( n41932,n41935,n41936 );
   nor U42712 ( n41929,n41937,n41938 );
   nor U42713 ( n41938,n28147,n39273 );
   nor U42714 ( n41937,n28154,n41939 );
   nand U42715 ( n41941,n28091,n41942 );
   not U42716 ( n41942,n41472 );
   nand U42717 ( n41472,n41943,n41944 );
   nand U42718 ( n41944,n41945,n41946 );
   not U42719 ( n41946,n41947 );
   nor U42720 ( n41945,n41948,n41949 );
   nor U42721 ( n41940,n41950,n41951 );
   nor U42722 ( n41951,n39292,n41764 );
   nor U42723 ( n41950,n28152,n41952 );
   nand U42724 ( n41954,n28091,n41955 );
   not U42725 ( n41955,n41488 );
   nand U42726 ( n41488,n41956,n41957 );
   nand U42727 ( n41957,n41958,n41959 );
   and U42728 ( n41958,n41943,n41960 );
   nor U42729 ( n41953,n41961,n41962 );
   nor U42730 ( n41962,n28148,n40098 );
   nor U42731 ( n41961,n41765,n41963 );
   nand U42732 ( n41965,n28091,n41966 );
   not U42733 ( n41966,n41504 );
   nand U42734 ( n41504,n41967,n41968 );
   nand U42735 ( n41968,n41969,n41970 );
   and U42736 ( n41969,n41956,n41971 );
   not U42737 ( n41956,n41972 );
   nor U42738 ( n41964,n41973,n41974 );
   nor U42739 ( n41974,n39340,n28147 );
   nor U42740 ( n41973,n28153,n41975 );
   nand U42741 ( n41977,n28091,n41978 );
   not U42742 ( n41978,n41520 );
   nand U42743 ( n41520,n41979,n41980 );
   nand U42744 ( n41980,n41981,n41982 );
   and U42745 ( n41981,n41967,n41983 );
   nor U42746 ( n41976,n41984,n41985 );
   nor U42747 ( n41985,n28147,n39369 );
   nor U42748 ( n41984,n28154,n41986 );
   nand U42749 ( n41988,n28091,n41989 );
   not U42750 ( n41989,n41536 );
   nand U42751 ( n41536,n41990,n41991 );
   nand U42752 ( n41991,n41992,n41993 );
   and U42753 ( n41992,n41979,n41994 );
   not U42754 ( n41979,n41995 );
   nor U42755 ( n41987,n41996,n41997 );
   nor U42756 ( n41997,n40159,n28147 );
   nor U42757 ( n41996,n28152,n41998 );
   nand U42758 ( n42000,n28091,n41551 );
   xor U42759 ( n41551,n42001,n42002 );
   nor U42760 ( n41999,n42003,n42004 );
   nor U42761 ( n42004,n41764,n39407 );
   nor U42762 ( n42003,n41765,n42005 );
   nand U42763 ( n42007,n28091,n41568 );
   xor U42764 ( n41568,n42008,n42009 );
   nand U42765 ( n42009,n42002,n42001 );
   nand U42766 ( n42001,n42010,n42011 );
   nand U42767 ( n42011,n42012,n28306 );
   xor U42768 ( n42012,n42013,n42014 );
   nand U42769 ( n42010,n42015,n42013 );
   not U42770 ( n42002,n41990 );
   nand U42771 ( n41990,n41995,n42016 );
   nand U42772 ( n42016,n41993,n41994 );
   nand U42773 ( n41994,n42017,n41798 );
   nor U42774 ( n42017,n42014,n42018 );
   nor U42775 ( n42018,n42019,n42020 );
   nand U42776 ( n41993,n42015,n42020 );
   nor U42777 ( n41995,n41967,n42021 );
   and U42778 ( n42021,n41983,n41982 );
   nand U42779 ( n41982,n42015,n42022 );
   nand U42780 ( n41983,n42023,n41798 );
   nor U42781 ( n42023,n42019,n42024 );
   nor U42782 ( n42024,n42025,n42022 );
   and U42783 ( n42025,n42026,n42027 );
   nand U42784 ( n41967,n41972,n42028 );
   nand U42785 ( n42028,n41971,n41970 );
   nand U42786 ( n41970,n42015,n42026 );
   nand U42787 ( n41971,n42029,n41798 );
   xor U42788 ( n42029,n42026,n42027 );
   nor U42789 ( n41972,n41943,n42030 );
   and U42790 ( n42030,n41960,n41959 );
   nand U42791 ( n41959,n42015,n42031 );
   nand U42792 ( n41960,n42032,n28306 );
   nor U42793 ( n42032,n42027,n42033 );
   nor U42794 ( n42033,n42034,n42031 );
   nor U42795 ( n42034,n42035,n42036 );
   nand U42796 ( n41943,n42037,n41947 );
   nand U42797 ( n41947,n41934,n42038 );
   nand U42798 ( n42038,n41922,n41935 );
   nor U42799 ( n41922,n41924,n41925 );
   nand U42800 ( n41925,n42039,n42040 );
   nand U42801 ( n42040,n42041,n42042 );
   nor U42802 ( n42042,n42043,n42044 );
   nand U42803 ( n42044,n42045,n42046 );
   nor U42804 ( n42046,n42047,n42048 );
   nor U42805 ( n42048,n40541,n42049 );
   nor U42806 ( n42047,n40542,n42050 );
   nor U42807 ( n42045,n42051,n42052 );
   nor U42808 ( n42052,n40545,n42053 );
   nor U42809 ( n42051,n40546,n42054 );
   nand U42810 ( n42043,n42055,n42056 );
   nor U42811 ( n42056,n42057,n42058 );
   nor U42812 ( n42058,n40532,n42059 );
   nor U42813 ( n42057,n40533,n42060 );
   nor U42814 ( n42055,n42061,n42062 );
   nor U42815 ( n42062,n40536,n42063 );
   nor U42816 ( n42061,n38590,n42064 );
   nor U42817 ( n42041,n42065,n42066 );
   nand U42818 ( n42066,n42067,n42068 );
   nor U42819 ( n42068,n42069,n42070 );
   nor U42820 ( n42070,n40520,n42071 );
   nor U42821 ( n42069,n40521,n42072 );
   nor U42822 ( n42067,n42073,n42074 );
   nor U42823 ( n42074,n40524,n42075 );
   nor U42824 ( n42073,n40525,n42076 );
   nand U42825 ( n42065,n42077,n42078 );
   nor U42826 ( n42078,n42079,n42080 );
   nor U42827 ( n42080,n40510,n42081 );
   nor U42828 ( n42079,n40511,n42082 );
   nor U42829 ( n42077,n42083,n42084 );
   nor U42830 ( n42084,n40514,n42085 );
   nor U42831 ( n42083,n40515,n42086 );
   nand U42832 ( n41924,n41907,n41916 );
   and U42833 ( n41916,n42087,n42039 );
   nand U42834 ( n42087,n42088,n42089 );
   nor U42835 ( n42089,n42090,n42091 );
   nand U42836 ( n42091,n42092,n42093 );
   nor U42837 ( n42093,n42094,n42095 );
   nor U42838 ( n42095,n40790,n42081 );
   nor U42839 ( n42094,n40791,n42082 );
   nor U42840 ( n42092,n42096,n42097 );
   nor U42841 ( n42097,n40794,n42085 );
   nor U42842 ( n42096,n40795,n42086 );
   nand U42843 ( n42090,n42098,n42099 );
   nor U42844 ( n42099,n42100,n42101 );
   nor U42845 ( n42101,n40780,n42071 );
   nor U42846 ( n42100,n40781,n42072 );
   nor U42847 ( n42098,n42102,n42103 );
   nor U42848 ( n42103,n40784,n42075 );
   nor U42849 ( n42102,n40785,n42076 );
   nor U42850 ( n42088,n42104,n42105 );
   nand U42851 ( n42105,n42106,n42107 );
   nor U42852 ( n42107,n42108,n42109 );
   nor U42853 ( n42109,n40769,n42059 );
   nor U42854 ( n42108,n40770,n42060 );
   nor U42855 ( n42106,n42110,n42111 );
   nor U42856 ( n42111,n40773,n42063 );
   nor U42857 ( n42110,n38606,n42064 );
   nand U42858 ( n42104,n42112,n42113 );
   nor U42859 ( n42113,n42114,n42115 );
   nor U42860 ( n42115,n40759,n42049 );
   nor U42861 ( n42114,n40760,n42050 );
   nor U42862 ( n42112,n42116,n42117 );
   nor U42863 ( n42117,n40763,n42053 );
   nor U42864 ( n42116,n40764,n42054 );
   nor U42865 ( n41907,n41909,n41910 );
   nand U42866 ( n41910,n42039,n42118 );
   nand U42867 ( n42118,n42119,n42120 );
   nor U42868 ( n42120,n42121,n42122 );
   nand U42869 ( n42122,n42123,n42124 );
   nor U42870 ( n42124,n42125,n42126 );
   nor U42871 ( n42126,n40848,n42049 );
   nor U42872 ( n42125,n40849,n42050 );
   nor U42873 ( n42123,n42127,n42128 );
   nor U42874 ( n42128,n40852,n42053 );
   nor U42875 ( n42127,n40853,n42054 );
   nand U42876 ( n42121,n42129,n42130 );
   nor U42877 ( n42130,n42131,n42132 );
   nor U42878 ( n42132,n40838,n42059 );
   nor U42879 ( n42131,n40839,n42060 );
   nor U42880 ( n42129,n42133,n42134 );
   nor U42881 ( n42134,n40842,n42063 );
   nor U42882 ( n42133,n38622,n42064 );
   nor U42883 ( n42119,n42135,n42136 );
   nand U42884 ( n42136,n42137,n42138 );
   nor U42885 ( n42138,n42139,n42140 );
   nor U42886 ( n42140,n40823,n42071 );
   nor U42887 ( n42139,n40825,n42072 );
   nor U42888 ( n42137,n42141,n42142 );
   nor U42889 ( n42142,n40828,n42075 );
   nor U42890 ( n42141,n40830,n42076 );
   nand U42891 ( n42135,n42143,n42144 );
   nor U42892 ( n42144,n42145,n42146 );
   nor U42893 ( n42146,n40808,n42081 );
   nor U42894 ( n42145,n40811,n42082 );
   nor U42895 ( n42143,n42147,n42148 );
   nor U42896 ( n42148,n40816,n42085 );
   nor U42897 ( n42147,n40817,n42086 );
   nand U42898 ( n41909,n41892,n41901 );
   and U42899 ( n41901,n42149,n42039 );
   nand U42900 ( n42149,n42150,n42151 );
   nor U42901 ( n42151,n42152,n42153 );
   nand U42902 ( n42153,n42154,n42155 );
   nor U42903 ( n42155,n42156,n42157 );
   nor U42904 ( n42157,n40591,n42081 );
   nor U42905 ( n42156,n40592,n42082 );
   nor U42906 ( n42154,n42158,n42159 );
   nor U42907 ( n42159,n40595,n42085 );
   nor U42908 ( n42158,n40596,n42086 );
   nand U42909 ( n42152,n42160,n42161 );
   nor U42910 ( n42161,n42162,n42163 );
   nor U42911 ( n42163,n40581,n42071 );
   nor U42912 ( n42162,n40582,n42072 );
   nor U42913 ( n42160,n42164,n42165 );
   nor U42914 ( n42165,n40585,n42075 );
   nor U42915 ( n42164,n40586,n42076 );
   nor U42916 ( n42150,n42166,n42167 );
   nand U42917 ( n42167,n42168,n42169 );
   nor U42918 ( n42169,n42170,n42171 );
   nor U42919 ( n42171,n40570,n42059 );
   nor U42920 ( n42170,n40571,n42060 );
   nor U42921 ( n42168,n42172,n42173 );
   nor U42922 ( n42173,n40574,n42063 );
   nor U42923 ( n42172,n38638,n42064 );
   nand U42924 ( n42166,n42174,n42175 );
   nor U42925 ( n42175,n42176,n42177 );
   nor U42926 ( n42177,n40560,n42049 );
   nor U42927 ( n42176,n40561,n42050 );
   nor U42928 ( n42174,n42178,n42179 );
   nor U42929 ( n42179,n40564,n42053 );
   nor U42930 ( n42178,n40565,n42054 );
   nor U42931 ( n41892,n41894,n41895 );
   nand U42932 ( n41895,n42039,n42180 );
   nand U42933 ( n42180,n42181,n42182 );
   nor U42934 ( n42182,n42183,n42184 );
   nand U42935 ( n42184,n42185,n42186 );
   nor U42936 ( n42186,n42187,n42188 );
   nor U42937 ( n42188,n40741,n42049 );
   nor U42938 ( n42187,n40742,n42050 );
   nor U42939 ( n42185,n42189,n42190 );
   nor U42940 ( n42190,n40745,n42053 );
   nor U42941 ( n42189,n40746,n42054 );
   nand U42942 ( n42183,n42191,n42192 );
   nor U42943 ( n42192,n42193,n42194 );
   nor U42944 ( n42194,n40732,n42059 );
   nor U42945 ( n42193,n40733,n42060 );
   nor U42946 ( n42191,n42195,n42196 );
   nor U42947 ( n42196,n40736,n42063 );
   nor U42948 ( n42195,n38654,n42064 );
   nor U42949 ( n42181,n42197,n42198 );
   nand U42950 ( n42198,n42199,n42200 );
   nor U42951 ( n42200,n42201,n42202 );
   nor U42952 ( n42202,n40720,n42071 );
   nor U42953 ( n42201,n40721,n42072 );
   nor U42954 ( n42199,n42203,n42204 );
   nor U42955 ( n42204,n40724,n42075 );
   nor U42956 ( n42203,n40725,n42076 );
   nand U42957 ( n42197,n42205,n42206 );
   nor U42958 ( n42206,n42207,n42208 );
   nor U42959 ( n42208,n40710,n42081 );
   nor U42960 ( n42207,n40711,n42082 );
   nor U42961 ( n42205,n42209,n42210 );
   nor U42962 ( n42210,n40714,n42085 );
   nor U42963 ( n42209,n40715,n42086 );
   nand U42964 ( n41894,n41878,n41886 );
   and U42965 ( n41886,n42211,n42039 );
   nand U42966 ( n42211,n42212,n42213 );
   nor U42967 ( n42213,n42214,n42215 );
   nand U42968 ( n42215,n42216,n42217 );
   nor U42969 ( n42217,n42218,n42219 );
   nor U42970 ( n42219,n40661,n42081 );
   nor U42971 ( n42218,n40662,n42082 );
   nor U42972 ( n42216,n42220,n42221 );
   nor U42973 ( n42221,n40665,n42085 );
   nor U42974 ( n42220,n40666,n42086 );
   nand U42975 ( n42214,n42222,n42223 );
   nor U42976 ( n42223,n42224,n42225 );
   nor U42977 ( n42225,n40671,n42071 );
   nor U42978 ( n42224,n40672,n42072 );
   nor U42979 ( n42222,n42226,n42227 );
   nor U42980 ( n42227,n40675,n42075 );
   nor U42981 ( n42226,n40676,n42076 );
   nor U42982 ( n42212,n42228,n42229 );
   nand U42983 ( n42229,n42230,n42231 );
   nor U42984 ( n42231,n42232,n42233 );
   nor U42985 ( n42233,n40683,n42059 );
   nor U42986 ( n42232,n40684,n42060 );
   nor U42987 ( n42230,n42234,n42235 );
   nor U42988 ( n42235,n40687,n42063 );
   nor U42989 ( n42234,n38669,n42064 );
   nand U42990 ( n42228,n42236,n42237 );
   nor U42991 ( n42237,n42238,n42239 );
   nor U42992 ( n42239,n40692,n42049 );
   nor U42993 ( n42238,n40693,n42050 );
   nor U42994 ( n42236,n42240,n42241 );
   nor U42995 ( n42241,n40696,n42053 );
   nor U42996 ( n42240,n40697,n42054 );
   nor U42997 ( n41878,n41880,n41879 );
   nand U42998 ( n41879,n42039,n42242 );
   nand U42999 ( n42242,n42243,n42244 );
   nor U43000 ( n42244,n42245,n42246 );
   nand U43001 ( n42246,n42247,n42248 );
   nor U43002 ( n42248,n42249,n42250 );
   nor U43003 ( n42250,n40643,n42049 );
   nor U43004 ( n42249,n40644,n42050 );
   nor U43005 ( n42247,n42251,n42252 );
   nor U43006 ( n42252,n40647,n42053 );
   nor U43007 ( n42251,n40648,n42054 );
   nand U43008 ( n42245,n42253,n42254 );
   nor U43009 ( n42254,n42255,n42256 );
   nor U43010 ( n42256,n40634,n42059 );
   nor U43011 ( n42255,n40635,n42060 );
   nor U43012 ( n42253,n42257,n42258 );
   nor U43013 ( n42258,n40638,n42063 );
   nor U43014 ( n42257,n38693,n42064 );
   nor U43015 ( n42243,n42259,n42260 );
   nand U43016 ( n42260,n42261,n42262 );
   nor U43017 ( n42262,n42263,n42264 );
   nor U43018 ( n42264,n40622,n42071 );
   nor U43019 ( n42263,n40623,n42072 );
   nor U43020 ( n42261,n42265,n42266 );
   nor U43021 ( n42266,n40626,n42075 );
   nor U43022 ( n42265,n40627,n42076 );
   nand U43023 ( n42259,n42267,n42268 );
   nor U43024 ( n42268,n42269,n42270 );
   nor U43025 ( n42270,n40612,n42081 );
   nor U43026 ( n42269,n40613,n42082 );
   nor U43027 ( n42267,n42271,n42272 );
   nor U43028 ( n42272,n40616,n42085 );
   nor U43029 ( n42271,n40617,n42086 );
   not U43030 ( n42039,n42273 );
   nand U43031 ( n41880,n41871,n41870 );
   nor U43032 ( n41871,n41850,n41861 );
   nand U43033 ( n41850,n42274,n41842 );
   nor U43034 ( n41842,n41836,n41835 );
   nand U43035 ( n41835,n41798,n42275 );
   nand U43036 ( n41836,n42276,n41829 );
   not U43037 ( n42276,n41818 );
   nand U43038 ( n41818,n42277,n41812 );
   and U43039 ( n41812,n41804,n41805 );
   and U43040 ( n41805,n41796,p2_instqueue_reg_0__6_ );
   nor U43041 ( n41804,n41862,n38572 );
   nor U43042 ( n42277,n41821,n41822 );
   nand U43043 ( n41822,n41798,n42278 );
   nand U43044 ( n41821,n41798,n42279 );
   nor U43045 ( n42274,n41853,n41854 );
   nand U43046 ( n41854,n41798,n42280 );
   nand U43047 ( n41853,n41798,n42281 );
   nand U43048 ( n41934,n41936,n41935 );
   and U43049 ( n41935,n42282,n42283 );
   nand U43050 ( n42283,n42284,n42285 );
   nand U43051 ( n42285,n41798,n42286 );
   nor U43052 ( n42282,n42273,n42287 );
   nor U43053 ( n42287,n42015,n42036 );
   nor U43054 ( n42273,n41798,n42015 );
   nor U43055 ( n41936,n42288,n42289 );
   or U43056 ( n42037,n41948,n41949 );
   nor U43057 ( n41949,n42289,n42035 );
   and U43058 ( n41948,n42290,n41798 );
   xor U43059 ( n42290,n42036,n42035 );
   not U43060 ( n42035,n42291 );
   not U43061 ( n42036,n42292 );
   nor U43062 ( n42008,n42293,n42294 );
   and U43063 ( n42294,n42295,n42015 );
   nor U43064 ( n42293,n41862,n42296 );
   xor U43065 ( n42296,n42297,n42295 );
   nand U43066 ( n42295,n42298,n42299 );
   nor U43067 ( n42299,n42300,n42301 );
   nand U43068 ( n42301,n42302,n42303 );
   nor U43069 ( n42303,n42304,n42305 );
   nor U43070 ( n42305,n40497,n42306 );
   nor U43071 ( n42304,n40462,n42307 );
   nor U43072 ( n42302,n42308,n42309 );
   nor U43073 ( n42309,n40484,n42310 );
   nor U43074 ( n42308,n40493,n42311 );
   nand U43075 ( n42300,n42312,n42313 );
   nor U43076 ( n42313,n42314,n42315 );
   nor U43077 ( n42315,n40461,n42316 );
   nor U43078 ( n42314,n38572,n42317 );
   nor U43079 ( n42312,n42318,n42319 );
   nor U43080 ( n42319,n40472,n42320 );
   nor U43081 ( n42318,n40475,n42321 );
   nor U43082 ( n42298,n42322,n42323 );
   nand U43083 ( n42323,n42324,n42325 );
   nor U43084 ( n42325,n42326,n42327 );
   nor U43085 ( n42327,n40476,n42328 );
   nor U43086 ( n42326,n40465,n42329 );
   nor U43087 ( n42324,n42330,n42331 );
   nor U43088 ( n42331,n40483,n42332 );
   nor U43089 ( n42330,n40492,n42333 );
   nand U43090 ( n42322,n42334,n42335 );
   nor U43091 ( n42335,n42336,n42337 );
   nor U43092 ( n42337,n40471,n42338 );
   nor U43093 ( n42336,n40466,n42339 );
   nor U43094 ( n42334,n42340,n42341 );
   nor U43095 ( n42341,n40496,n42342 );
   nor U43096 ( n42340,n40487,n42343 );
   nand U43097 ( n42297,n42014,n42013 );
   nand U43098 ( n42013,n42344,n42345 );
   nor U43099 ( n42345,n42346,n42347 );
   nand U43100 ( n42347,n42348,n42349 );
   nor U43101 ( n42349,n42350,n42351 );
   nor U43102 ( n42351,n40546,n42306 );
   nor U43103 ( n42350,n40511,n42307 );
   nor U43104 ( n42348,n42352,n42353 );
   nor U43105 ( n42353,n40533,n42310 );
   nor U43106 ( n42352,n40542,n42311 );
   nand U43107 ( n42346,n42354,n42355 );
   nor U43108 ( n42355,n42356,n42357 );
   nor U43109 ( n42357,n40510,n42316 );
   nor U43110 ( n42356,n38590,n42317 );
   nor U43111 ( n42354,n42358,n42359 );
   nor U43112 ( n42359,n40521,n42320 );
   nor U43113 ( n42358,n40524,n42321 );
   nor U43114 ( n42344,n42360,n42361 );
   nand U43115 ( n42361,n42362,n42363 );
   nor U43116 ( n42363,n42364,n42365 );
   nor U43117 ( n42365,n40525,n42328 );
   nor U43118 ( n42364,n40514,n42329 );
   nor U43119 ( n42362,n42366,n42367 );
   nor U43120 ( n42367,n40532,n42332 );
   nor U43121 ( n42366,n40541,n42333 );
   nand U43122 ( n42360,n42368,n42369 );
   nor U43123 ( n42369,n42370,n42371 );
   nor U43124 ( n42371,n40520,n42338 );
   nor U43125 ( n42370,n40515,n42339 );
   nor U43126 ( n42368,n42372,n42373 );
   nor U43127 ( n42373,n40545,n42342 );
   nor U43128 ( n42372,n40536,n42343 );
   and U43129 ( n42014,n42019,n42020 );
   nand U43130 ( n42020,n42374,n42375 );
   nor U43131 ( n42375,n42376,n42377 );
   nand U43132 ( n42377,n42378,n42379 );
   nor U43133 ( n42379,n42380,n42381 );
   nor U43134 ( n42381,n40764,n42306 );
   nor U43135 ( n42380,n40791,n42307 );
   nor U43136 ( n42378,n42382,n42383 );
   nor U43137 ( n42383,n40770,n42310 );
   nor U43138 ( n42382,n40760,n42311 );
   nand U43139 ( n42376,n42384,n42385 );
   nor U43140 ( n42385,n42386,n42387 );
   nor U43141 ( n42387,n40790,n42316 );
   nor U43142 ( n42386,n38606,n42317 );
   nor U43143 ( n42384,n42388,n42389 );
   nor U43144 ( n42389,n40781,n42320 );
   nor U43145 ( n42388,n40784,n42321 );
   nor U43146 ( n42374,n42390,n42391 );
   nand U43147 ( n42391,n42392,n42393 );
   nor U43148 ( n42393,n42394,n42395 );
   nor U43149 ( n42395,n40785,n42328 );
   nor U43150 ( n42394,n40794,n42329 );
   nor U43151 ( n42392,n42396,n42397 );
   nor U43152 ( n42397,n40769,n42332 );
   nor U43153 ( n42396,n40759,n42333 );
   nand U43154 ( n42390,n42398,n42399 );
   nor U43155 ( n42399,n42400,n42401 );
   nor U43156 ( n42401,n40780,n42338 );
   nor U43157 ( n42400,n40795,n42339 );
   nor U43158 ( n42398,n42402,n42403 );
   nor U43159 ( n42403,n40763,n42342 );
   nor U43160 ( n42402,n40773,n42343 );
   and U43161 ( n42019,n42404,n42027 );
   and U43162 ( n42027,n42405,n42292 );
   nor U43163 ( n42292,n42288,n42284 );
   and U43164 ( n42284,n42406,n42407 );
   nor U43165 ( n42407,n42408,n42409 );
   nand U43166 ( n42409,n42410,n42411 );
   nor U43167 ( n42411,n42412,n42413 );
   nor U43168 ( n42413,n40461,n42081 );
   nand U43169 ( n42081,n42414,n42415 );
   nor U43170 ( n42412,n40462,n42082 );
   nand U43171 ( n42082,n42414,n42416 );
   nor U43172 ( n42410,n42417,n42418 );
   nor U43173 ( n42418,n40465,n42085 );
   nand U43174 ( n42085,n42414,n42419 );
   nor U43175 ( n42417,n40466,n42086 );
   nand U43176 ( n42086,n42420,n42415 );
   nand U43177 ( n42408,n42421,n42422 );
   nor U43178 ( n42422,n42423,n42424 );
   nor U43179 ( n42424,n40471,n42071 );
   nand U43180 ( n42071,n42420,n42416 );
   nor U43181 ( n42423,n40472,n42072 );
   nand U43182 ( n42072,n42420,n42419 );
   nor U43183 ( n42421,n42425,n42426 );
   nor U43184 ( n42426,n40475,n42075 );
   nand U43185 ( n42075,n42427,n42415 );
   nor U43186 ( n42425,n40476,n42076 );
   nand U43187 ( n42076,n42427,n42416 );
   nor U43188 ( n42406,n42428,n42429 );
   nand U43189 ( n42429,n42430,n42431 );
   nor U43190 ( n42431,n42432,n42433 );
   nor U43191 ( n42433,n40483,n42059 );
   nand U43192 ( n42059,n42427,n42419 );
   nor U43193 ( n42432,n40484,n42060 );
   nand U43194 ( n42060,n42434,n42415 );
   nor U43195 ( n42430,n42435,n42436 );
   nor U43196 ( n42436,n40487,n42063 );
   nand U43197 ( n42063,n42434,n42416 );
   nor U43198 ( n42435,n38572,n42064 );
   nand U43199 ( n42064,n42434,n42419 );
   nand U43200 ( n42428,n42437,n42438 );
   nor U43201 ( n42438,n42439,n42440 );
   nor U43202 ( n42440,n40492,n42049 );
   nand U43203 ( n42049,n42414,n42441 );
   nor U43204 ( n42414,n42442,n42443 );
   nor U43205 ( n42439,n40493,n42050 );
   nand U43206 ( n42050,n42420,n42441 );
   nor U43207 ( n42420,n42443,n42444 );
   not U43208 ( n42443,n42445 );
   nor U43209 ( n42437,n42446,n42447 );
   nor U43210 ( n42447,n40496,n42053 );
   nand U43211 ( n42053,n42427,n42441 );
   nor U43212 ( n42427,n42442,n42445 );
   not U43213 ( n42442,n42444 );
   nor U43214 ( n42446,n40497,n42054 );
   nand U43215 ( n42054,n42434,n42441 );
   nor U43216 ( n42434,n42445,n42444 );
   nor U43217 ( n42444,n42448,n42449 );
   xor U43218 ( n42445,n42448,p2_instqueuerd_addr_reg_3_ );
   nor U43219 ( n42448,n37154,n42450 );
   not U43220 ( n42288,n42286 );
   nand U43221 ( n42286,n42451,n42452 );
   nor U43222 ( n42452,n42453,n42454 );
   nand U43223 ( n42454,n42455,n42456 );
   nor U43224 ( n42456,n42457,n42458 );
   nor U43225 ( n42458,n40648,n42306 );
   nor U43226 ( n42457,n40613,n42307 );
   nor U43227 ( n42455,n42459,n42460 );
   nor U43228 ( n42460,n40635,n42310 );
   nor U43229 ( n42459,n40644,n42311 );
   nand U43230 ( n42453,n42461,n42462 );
   nor U43231 ( n42462,n42463,n42464 );
   nor U43232 ( n42464,n40612,n42316 );
   nor U43233 ( n42463,n38693,n42317 );
   nor U43234 ( n42461,n42465,n42466 );
   nor U43235 ( n42466,n40623,n42320 );
   nor U43236 ( n42465,n40626,n42321 );
   nor U43237 ( n42451,n42467,n42468 );
   nand U43238 ( n42468,n42469,n42470 );
   nor U43239 ( n42470,n42471,n42472 );
   nor U43240 ( n42472,n40627,n42328 );
   nor U43241 ( n42471,n40616,n42329 );
   nor U43242 ( n42469,n42473,n42474 );
   nor U43243 ( n42474,n40634,n42332 );
   nor U43244 ( n42473,n40643,n42333 );
   nand U43245 ( n42467,n42475,n42476 );
   nor U43246 ( n42476,n42477,n42478 );
   nor U43247 ( n42478,n40622,n42338 );
   nor U43248 ( n42477,n40617,n42339 );
   nor U43249 ( n42475,n42479,n42480 );
   nor U43250 ( n42480,n40647,n42342 );
   nor U43251 ( n42479,n40638,n42343 );
   and U43252 ( n42405,n42291,n42031 );
   nand U43253 ( n42031,n42481,n42482 );
   nor U43254 ( n42482,n42483,n42484 );
   nand U43255 ( n42484,n42485,n42486 );
   nor U43256 ( n42486,n42487,n42488 );
   nor U43257 ( n42488,n40746,n42306 );
   nor U43258 ( n42487,n40711,n42307 );
   nor U43259 ( n42485,n42489,n42490 );
   nor U43260 ( n42490,n40733,n42310 );
   nor U43261 ( n42489,n40742,n42311 );
   nand U43262 ( n42483,n42491,n42492 );
   nor U43263 ( n42492,n42493,n42494 );
   nor U43264 ( n42494,n40710,n42316 );
   nor U43265 ( n42493,n38654,n42317 );
   nor U43266 ( n42491,n42495,n42496 );
   nor U43267 ( n42496,n40721,n42320 );
   nor U43268 ( n42495,n40724,n42321 );
   nor U43269 ( n42481,n42497,n42498 );
   nand U43270 ( n42498,n42499,n42500 );
   nor U43271 ( n42500,n42501,n42502 );
   nor U43272 ( n42502,n40725,n42328 );
   nor U43273 ( n42501,n40714,n42329 );
   nor U43274 ( n42499,n42503,n42504 );
   nor U43275 ( n42504,n40732,n42332 );
   nor U43276 ( n42503,n40741,n42333 );
   nand U43277 ( n42497,n42505,n42506 );
   nor U43278 ( n42506,n42507,n42508 );
   nor U43279 ( n42508,n40720,n42338 );
   nor U43280 ( n42507,n40715,n42339 );
   nor U43281 ( n42505,n42509,n42510 );
   nor U43282 ( n42510,n40745,n42342 );
   nor U43283 ( n42509,n40736,n42343 );
   nand U43284 ( n42291,n42511,n42512 );
   nor U43285 ( n42512,n42513,n42514 );
   nand U43286 ( n42514,n42515,n42516 );
   nor U43287 ( n42516,n42517,n42518 );
   nor U43288 ( n42518,n40697,n42306 );
   nor U43289 ( n42517,n40662,n42307 );
   nor U43290 ( n42515,n42519,n42520 );
   nor U43291 ( n42520,n40684,n42310 );
   nor U43292 ( n42519,n40693,n42311 );
   nand U43293 ( n42513,n42521,n42522 );
   nor U43294 ( n42522,n42523,n42524 );
   nor U43295 ( n42524,n40661,n42316 );
   nor U43296 ( n42523,n38669,n42317 );
   nor U43297 ( n42521,n42525,n42526 );
   nor U43298 ( n42526,n40672,n42320 );
   nor U43299 ( n42525,n40675,n42321 );
   nor U43300 ( n42511,n42527,n42528 );
   nand U43301 ( n42528,n42529,n42530 );
   nor U43302 ( n42530,n42531,n42532 );
   nor U43303 ( n42532,n40676,n42328 );
   nor U43304 ( n42531,n40665,n42329 );
   nor U43305 ( n42529,n42533,n42534 );
   nor U43306 ( n42534,n40683,n42332 );
   nor U43307 ( n42533,n40692,n42333 );
   nand U43308 ( n42527,n42535,n42536 );
   nor U43309 ( n42536,n42537,n42538 );
   nor U43310 ( n42538,n40671,n42338 );
   nor U43311 ( n42537,n40666,n42339 );
   nor U43312 ( n42535,n42539,n42540 );
   nor U43313 ( n42540,n40696,n42342 );
   nor U43314 ( n42539,n40687,n42343 );
   and U43315 ( n42404,n42026,n42022 );
   nand U43316 ( n42022,n42541,n42542 );
   nor U43317 ( n42542,n42543,n42544 );
   nand U43318 ( n42544,n42545,n42546 );
   nor U43319 ( n42546,n42547,n42548 );
   nor U43320 ( n42548,n40853,n42306 );
   nor U43321 ( n42547,n40811,n42307 );
   nor U43322 ( n42545,n42549,n42550 );
   nor U43323 ( n42550,n40839,n42310 );
   nor U43324 ( n42549,n40849,n42311 );
   nand U43325 ( n42543,n42551,n42552 );
   nor U43326 ( n42552,n42553,n42554 );
   nor U43327 ( n42554,n40808,n42316 );
   nor U43328 ( n42553,n38622,n42317 );
   nor U43329 ( n42551,n42555,n42556 );
   nor U43330 ( n42556,n40825,n42320 );
   nor U43331 ( n42555,n40828,n42321 );
   nor U43332 ( n42541,n42557,n42558 );
   nand U43333 ( n42558,n42559,n42560 );
   nor U43334 ( n42560,n42561,n42562 );
   nor U43335 ( n42562,n40830,n42328 );
   nor U43336 ( n42561,n40816,n42329 );
   nor U43337 ( n42559,n42563,n42564 );
   nor U43338 ( n42564,n40838,n42332 );
   nor U43339 ( n42563,n40848,n42333 );
   nand U43340 ( n42557,n42565,n42566 );
   nor U43341 ( n42566,n42567,n42568 );
   nor U43342 ( n42568,n40823,n42338 );
   nor U43343 ( n42567,n40817,n42339 );
   nor U43344 ( n42565,n42569,n42570 );
   nor U43345 ( n42570,n40852,n42342 );
   nor U43346 ( n42569,n40842,n42343 );
   nand U43347 ( n42026,n42571,n42572 );
   nor U43348 ( n42572,n42573,n42574 );
   nand U43349 ( n42574,n42575,n42576 );
   nor U43350 ( n42576,n42577,n42578 );
   nor U43351 ( n42578,n40565,n42306 );
   nand U43352 ( n42306,n42579,n42580 );
   nor U43353 ( n42577,n40592,n42307 );
   nand U43354 ( n42307,n42581,n42582 );
   nor U43355 ( n42581,p2_instqueuerd_addr_reg_2_,n42579 );
   nor U43356 ( n42575,n42583,n42584 );
   nor U43357 ( n42584,n40571,n42310 );
   nand U43358 ( n42310,n42579,n42585 );
   nor U43359 ( n42583,n40561,n42311 );
   nand U43360 ( n42311,n42580,n42586 );
   nand U43361 ( n42573,n42587,n42588 );
   nor U43362 ( n42588,n42589,n42590 );
   nor U43363 ( n42590,n40591,n42316 );
   nand U43364 ( n42316,n42591,n42586 );
   nor U43365 ( n42589,n38638,n42317 );
   nand U43366 ( n42317,n42579,n42592 );
   nor U43367 ( n42587,n42593,n42594 );
   nor U43368 ( n42594,n40582,n42320 );
   nand U43369 ( n42320,n42592,n42586 );
   nor U43370 ( n42593,n40585,n42321 );
   nand U43371 ( n42321,n42579,n42591 );
   nor U43372 ( n42571,n42595,n42596 );
   nand U43373 ( n42596,n42597,n42598 );
   nor U43374 ( n42598,n42599,n42600 );
   nor U43375 ( n42600,n40586,n42328 );
   nand U43376 ( n42328,n42601,n42579 );
   nor U43377 ( n42601,p2_instqueuerd_addr_reg_2_,n42602 );
   nor U43378 ( n42599,n40595,n42329 );
   nand U43379 ( n42329,n42449,n42586 );
   nor U43380 ( n42597,n42603,n42604 );
   nor U43381 ( n42604,n40570,n42332 );
   nand U43382 ( n42332,n42579,n42449 );
   nor U43383 ( n42603,n40560,n42333 );
   nand U43384 ( n42333,n42605,n42586 );
   nand U43385 ( n42595,n42606,n42607 );
   nor U43386 ( n42607,n42608,n42609 );
   nor U43387 ( n42609,n40581,n42338 );
   nand U43388 ( n42338,n42610,n42586 );
   nor U43389 ( n42608,n40596,n42339 );
   nand U43390 ( n42339,n42585,n42586 );
   nor U43391 ( n42606,n42611,n42612 );
   nor U43392 ( n42612,n40564,n42342 );
   nand U43393 ( n42342,n42579,n42605 );
   nor U43394 ( n42611,n40574,n42343 );
   nand U43395 ( n42343,n42579,n42610 );
   not U43396 ( n42579,n42586 );
   xor U43397 ( n42586,p2_instqueuerd_addr_reg_3_,p2_instqueuerd_addr_reg_2_ );
   nor U43398 ( n41761,n28147,n39566 );
   nor U43399 ( n42006,n42613,n42614 );
   nor U43400 ( n42614,n40191,n41764 );
   nor U43401 ( n42613,n28153,n42615 );
   nand U43402 ( n42617,p2_ebx_reg_31_,n28147 );
   nand U43403 ( n42616,n39461,n41765 );
   not U43404 ( n41765,n41764 );
   nand U43405 ( n41764,n37045,n42618 );
   nand U43406 ( n42618,n42619,n39507 );
   nand U43407 ( n42619,n37180,n37168 );
   not U43408 ( n37168,n37166 );
   not U43409 ( n37180,n37167 );
   nand U43410 ( n37167,n42620,n37134 );
   and U43411 ( n37134,n42621,n42622 );
   and U43412 ( n42621,n38617,n41567 );
   nor U43413 ( n42620,n38649,n37132 );
   nor U43414 ( n42624,n42625,n42626 );
   nand U43415 ( n42626,n42627,n42628 );
   nand U43416 ( n42628,n28355,n36670 );
   nor U43417 ( n36670,n42630,n42631 );
   and U43418 ( n42631,n42632,n42633 );
   nand U43419 ( n42627,n28093,n37116 );
   not U43420 ( n37116,n38726 );
   nand U43421 ( n42625,n42635,n42636 );
   nand U43422 ( n42636,p2_phyaddrpointer_reg_0_,n42637 );
   nand U43423 ( n42637,n42638,n42639 );
   nand U43424 ( n42635,n42640,n36729 );
   not U43425 ( n36729,n36674 );
   nand U43426 ( n36674,n42641,n42642 );
   nand U43427 ( n42642,n42643,n42644 );
   nor U43428 ( n42644,p2_state2_reg_3_,n42645 );
   nor U43429 ( n42645,n38693,n41862 );
   nor U43430 ( n42643,n36783,n38585 );
   nor U43431 ( n42623,n42646,n42647 );
   nand U43432 ( n42647,n42648,n42649 );
   nand U43433 ( n42649,n42650,n42651 );
   nand U43434 ( n42648,n28122,p2_reip_reg_0_ );
   nand U43435 ( n42646,n42653,n42654 );
   nand U43436 ( n42654,n42655,n42656 );
   nand U43437 ( n42653,n28360,p2_ebx_reg_0_ );
   nor U43438 ( n42659,n42660,n42661 );
   nand U43439 ( n42661,n42662,n42663 );
   or U43440 ( n42663,n40348,n42664 );
   nand U43441 ( n40348,n40355,n42665 );
   nand U43442 ( n42665,n42651,p2_ebx_reg_1_ );
   nand U43443 ( n42662,n42640,n36740 );
   not U43444 ( n36740,n36684 );
   xor U43445 ( n36684,n42666,n42667 );
   nand U43446 ( n42667,n42668,n42669 );
   nand U43447 ( n42660,n42670,n42671 );
   nand U43448 ( n42671,n42655,n42672 );
   xor U43449 ( n42672,n36759,n36763 );
   nand U43450 ( n42670,n42629,n36680 );
   xor U43451 ( n36680,n42673,n42674 );
   xor U43452 ( n42673,n42630,n42675 );
   nor U43453 ( n42658,n42676,n42677 );
   nand U43454 ( n42677,n42678,n42679 );
   nand U43455 ( n42679,n28122,p2_reip_reg_1_ );
   nor U43456 ( n42678,n42680,n42681 );
   nor U43457 ( n42681,n39621,n42638 );
   not U43458 ( n42638,n42682 );
   nor U43459 ( n42680,p2_phyaddrpointer_reg_1_,n42639 );
   nand U43460 ( n42676,n42683,n42684 );
   nand U43461 ( n42684,n42634,n38745 );
   nand U43462 ( n42683,n42657,p2_ebx_reg_1_ );
   nor U43463 ( n42686,n42687,n42688 );
   nand U43464 ( n42688,n42689,n42690 );
   nand U43465 ( n42690,n42640,n36752 );
   not U43466 ( n36752,n36697 );
   nand U43467 ( n36697,n42691,n42692 );
   or U43468 ( n42692,n42693,n42694 );
   nand U43469 ( n42691,n42695,n42696 );
   nand U43470 ( n42696,n42668,n42666 );
   nor U43471 ( n42695,n42697,n42698 );
   nor U43472 ( n42698,n42694,n42699 );
   not U43473 ( n42694,n42700 );
   nand U43474 ( n42689,n42634,n38766 );
   not U43475 ( n38766,n37189 );
   nand U43476 ( n42687,n42701,n42702 );
   nand U43477 ( n42702,n28355,n36694 );
   not U43478 ( n36694,n41238 );
   xor U43479 ( n41238,n42703,n42704 );
   xor U43480 ( n42703,n42705,n42706 );
   nor U43481 ( n42701,n42707,n42708 );
   nor U43482 ( n42708,n42709,n42664 );
   xor U43483 ( n42709,n40354,n42710 );
   nor U43484 ( n42707,n27898,n42712 );
   nand U43485 ( n42712,n42713,n42714 );
   nand U43486 ( n42713,n39639,n42715 );
   nand U43487 ( n42715,n36759,n36763 );
   nor U43488 ( n42685,n42716,n42717 );
   nand U43489 ( n42717,n42718,n42719 );
   nand U43490 ( n42719,n42657,p2_ebx_reg_2_ );
   nand U43491 ( n42718,n28122,p2_reip_reg_2_ );
   nand U43492 ( n42716,n42720,n42721 );
   nand U43493 ( n42721,n28340,n39639 );
   nand U43494 ( n42720,n28092,p2_phyaddrpointer_reg_2_ );
   nor U43495 ( n42724,n42725,n42726 );
   nand U43496 ( n42726,n42727,n42728 );
   nand U43497 ( n42728,n42640,n36772 );
   xor U43498 ( n36772,n42729,n42730 );
   nor U43499 ( n42729,n42731,n42732 );
   not U43500 ( n42732,n42733 );
   nor U43501 ( n42731,n42734,n42735 );
   nor U43502 ( n42734,n38638,n41862 );
   not U43503 ( n42640,n42736 );
   nand U43504 ( n42727,n42634,n40843 );
   not U43505 ( n40843,n37159 );
   nand U43506 ( n42725,n42737,n42738 );
   nand U43507 ( n42738,n42650,n40334 );
   and U43508 ( n40334,n42739,n42740 );
   nand U43509 ( n42740,n42741,n40352 );
   nor U43510 ( n42737,n42742,n42743 );
   nor U43511 ( n42743,n38795,n42744 );
   xor U43512 ( n38795,n42745,n42746 );
   xor U43513 ( n42746,n42747,n42748 );
   nor U43514 ( n42742,n42711,n42749 );
   xor U43515 ( n42749,n39660,n42750 );
   nor U43516 ( n42723,n42751,n42752 );
   nand U43517 ( n42752,n42753,n42754 );
   nand U43518 ( n42754,n42657,p2_ebx_reg_3_ );
   nand U43519 ( n42753,n42652,p2_reip_reg_3_ );
   nand U43520 ( n42751,n42755,n42756 );
   nand U43521 ( n42756,n42722,n39660 );
   nand U43522 ( n42755,n28092,p2_phyaddrpointer_reg_3_ );
   nor U43523 ( n42758,n42759,n42760 );
   nand U43524 ( n42760,n42761,n42762 );
   nand U43525 ( n42762,n28355,n38812 );
   not U43526 ( n38812,n41257 );
   xor U43527 ( n41257,n42763,n42764 );
   xor U43528 ( n42763,n42765,n42766 );
   nand U43529 ( n42761,n42634,n38813 );
   not U43530 ( n38813,n39674 );
   xor U43531 ( n39674,n42767,n42768 );
   nand U43532 ( n42759,n42769,n42770 );
   nand U43533 ( n42770,n28331,n42771 );
   xor U43534 ( n42771,n42739,n40328 );
   nor U43535 ( n42769,n27897,n42773 );
   nor U43536 ( n42773,n27898,n42774 );
   nand U43537 ( n42774,n42775,n42776 );
   nand U43538 ( n42775,n39679,n42777 );
   or U43539 ( n42777,n42714,n39660 );
   nor U43540 ( n42757,n42778,n42779 );
   nand U43541 ( n42779,n42780,n42781 );
   nand U43542 ( n42781,n42657,p2_ebx_reg_4_ );
   nand U43543 ( n42780,n42652,p2_reip_reg_4_ );
   nand U43544 ( n42778,n42782,n42783 );
   nand U43545 ( n42783,n42682,p2_phyaddrpointer_reg_4_ );
   nor U43546 ( n42782,n42784,n42785 );
   nor U43547 ( n42785,n42786,n42639 );
   nor U43548 ( n42784,n41260,n42736 );
   nand U43549 ( n41260,n42787,n42788 );
   nand U43550 ( n42788,n42789,n42790 );
   not U43551 ( n42790,n42791 );
   nor U43552 ( n42789,n42792,n42793 );
   and U43553 ( n42792,n38585,p2_instqueuerd_addr_reg_4_ );
   nor U43554 ( n42795,n42796,n42797 );
   nand U43555 ( n42797,n42798,n42799 );
   nand U43556 ( n42799,n28355,n38839 );
   not U43557 ( n38839,n41270 );
   xor U43558 ( n41270,n42800,n42801 );
   xor U43559 ( n42800,n42802,n42803 );
   nand U43560 ( n42798,n42634,n38840 );
   xor U43561 ( n38840,n42804,n42805 );
   nand U43562 ( n42805,n42768,n42806 );
   nand U43563 ( n42796,n42807,n42808 );
   nand U43564 ( n42808,n42809,n42655 );
   xor U43565 ( n42809,n42776,n39699 );
   nor U43566 ( n42807,n42772,n42810 );
   nor U43567 ( n42810,n42664,n42811 );
   nand U43568 ( n42811,n40360,n40359 );
   nand U43569 ( n40360,n42812,n42813 );
   nand U43570 ( n42813,n42814,n41793 );
   nor U43571 ( n42812,n42815,n42816 );
   nor U43572 ( n42816,n40328,n42739 );
   not U43573 ( n42739,n40329 );
   nor U43574 ( n42794,n42817,n42818 );
   nand U43575 ( n42818,n42819,n42820 );
   nand U43576 ( n42820,n42657,p2_ebx_reg_5_ );
   nand U43577 ( n42819,n28122,p2_reip_reg_5_ );
   nand U43578 ( n42817,n42821,n42822 );
   nand U43579 ( n42822,n42682,p2_phyaddrpointer_reg_5_ );
   nor U43580 ( n42821,n42823,n42824 );
   nor U43581 ( n42824,n42825,n42639 );
   nor U43582 ( n42823,n41683,n42736 );
   nand U43583 ( n42736,n42826,n39573 );
   not U43584 ( n41683,n41790 );
   nor U43585 ( n41790,n41796,n42827 );
   and U43586 ( n42827,n42828,n42787 );
   nand U43587 ( n42828,n41798,p2_instqueue_reg_0__5_ );
   nor U43588 ( n41796,n42787,n38606 );
   nand U43589 ( n42787,n42791,n42793 );
   nor U43590 ( n42793,n41862,n38622 );
   nand U43591 ( n42791,n42733,n42829 );
   nand U43592 ( n42829,n42830,n42730 );
   nand U43593 ( n42730,n42700,n42693 );
   nand U43594 ( n42693,n42831,n42832 );
   or U43595 ( n42832,n42666,n42697 );
   not U43596 ( n42697,n42669 );
   nand U43597 ( n42669,n42833,n28306 );
   nor U43598 ( n42833,n42641,n38669 );
   nand U43599 ( n42666,n42834,n42835 );
   nand U43600 ( n42835,p2_instqueuerd_addr_reg_1_,n42836 );
   nor U43601 ( n42834,n42837,n42838 );
   nor U43602 ( n42838,n37125,n40877 );
   not U43603 ( n37125,n38745 );
   xor U43604 ( n38745,n42839,n42840 );
   xor U43605 ( n42839,n42841,n42842 );
   nor U43606 ( n42837,n38117,n38704 );
   nor U43607 ( n38117,n37520,n37433 );
   nor U43608 ( n37433,n37096,p2_instqueuewr_addr_reg_0_ );
   nor U43609 ( n37520,n37336,p2_instqueuewr_addr_reg_1_ );
   nor U43610 ( n42831,n42843,n42699 );
   and U43611 ( n42699,n42844,n42845 );
   nor U43612 ( n42845,n42846,n42847 );
   not U43613 ( n42847,n42848 );
   nor U43614 ( n42846,n38116,n38704 );
   not U43615 ( n38116,n38456 );
   xor U43616 ( n38456,p2_instqueuewr_addr_reg_2_,n37346 );
   nor U43617 ( n42844,n42849,n42850 );
   nor U43618 ( n42850,n38654,n41862 );
   nor U43619 ( n42849,n40877,n37189 );
   xor U43620 ( n37189,n42851,n42852 );
   xor U43621 ( n42851,n42853,n42854 );
   not U43622 ( n42843,n42668 );
   nand U43623 ( n42668,n42641,n42855 );
   nand U43624 ( n42855,n41798,p2_instqueue_reg_0__1_ );
   and U43625 ( n42641,n42856,n42857 );
   nand U43626 ( n42857,n36628,n37336 );
   nor U43627 ( n42856,n42858,n42859 );
   nor U43628 ( n42859,n40877,n38726 );
   nand U43629 ( n38726,n42841,n42860 );
   nand U43630 ( n42860,n42861,n42862 );
   nor U43631 ( n42861,n42863,n42864 );
   and U43632 ( n42858,n42836,p2_instqueuerd_addr_reg_0_ );
   nand U43633 ( n42700,n42865,n28306 );
   nor U43634 ( n42865,n42848,n38654 );
   nand U43635 ( n42848,p2_instqueuerd_addr_reg_2_,n42836 );
   nand U43636 ( n42830,n42866,n42867 );
   nand U43637 ( n42867,n41798,p2_instqueue_reg_0__3_ );
   nand U43638 ( n42733,n42868,n41798 );
   not U43639 ( n41798,n41862 );
   nand U43640 ( n41862,n40220,n39515 );
   nor U43641 ( n42868,n42866,n38638 );
   not U43642 ( n42866,n42735 );
   nand U43643 ( n42735,n42869,n42870 );
   nand U43644 ( n42870,p2_instqueuerd_addr_reg_3_,n42836 );
   nand U43645 ( n42836,n38681,n42871 );
   nand U43646 ( n42871,n42872,n38585 );
   or U43647 ( n42872,n42873,n40220 );
   nor U43648 ( n40220,n36783,n39545 );
   nor U43649 ( n42869,n42874,n42875 );
   nor U43650 ( n42875,n37159,n40877 );
   not U43651 ( n40877,n36634 );
   nor U43652 ( n36634,n37217,p2_state2_reg_0_ );
   xor U43653 ( n37159,n42876,n42877 );
   xor U43654 ( n42876,n42878,n42879 );
   nor U43655 ( n42874,n38115,n38704 );
   not U43656 ( n38115,n37427 );
   nand U43657 ( n37427,n42880,n42881 );
   or U43658 ( n42881,n37606,n37346 );
   nor U43659 ( n42880,n37697,n38024 );
   not U43660 ( n38024,n37961 );
   nand U43661 ( n37961,n38122,n37346 );
   nor U43662 ( n37346,n37336,n37096 );
   nor U43663 ( n38122,n37607,p2_instqueuewr_addr_reg_3_ );
   nor U43664 ( n37697,n37606,p2_instqueuewr_addr_reg_2_ );
   nor U43665 ( n42883,n42884,n42885 );
   nand U43666 ( n42885,n42886,n42887 );
   nand U43667 ( n42887,n42634,n38859 );
   not U43668 ( n38859,n39713 );
   nand U43669 ( n39713,n42888,n42889 );
   or U43670 ( n42888,n42890,n42891 );
   nand U43671 ( n42886,n28355,n38858 );
   not U43672 ( n38858,n41281 );
   xor U43673 ( n41281,n42892,n42893 );
   xor U43674 ( n42892,n42894,n42895 );
   nand U43675 ( n42884,n42896,n42897 );
   nand U43676 ( n42897,n42650,n42898 );
   xor U43677 ( n42898,n42899,n40318 );
   nor U43678 ( n42896,n27897,n42900 );
   nor U43679 ( n42900,n27898,n42901 );
   nand U43680 ( n42901,n42902,n42903 );
   nand U43681 ( n42902,n39718,n42904 );
   nand U43682 ( n42904,n42905,n42825 );
   not U43683 ( n42825,n39699 );
   nor U43684 ( n42882,n42906,n42907 );
   nand U43685 ( n42907,n42908,n42909 );
   nand U43686 ( n42909,n42657,p2_ebx_reg_6_ );
   nand U43687 ( n42908,n28122,p2_reip_reg_6_ );
   nand U43688 ( n42906,n42910,n42911 );
   nand U43689 ( n42911,n28340,n39718 );
   nand U43690 ( n42910,n42682,p2_phyaddrpointer_reg_6_ );
   nor U43691 ( n42913,n42914,n42915 );
   nand U43692 ( n42915,n42916,n42917 );
   nand U43693 ( n42917,n42634,n38888 );
   not U43694 ( n38888,n39733 );
   xor U43695 ( n39733,n42918,n42919 );
   nand U43696 ( n42916,n28355,n38887 );
   not U43697 ( n38887,n41292 );
   xor U43698 ( n41292,n42920,n42921 );
   xor U43699 ( n42920,n42922,n42923 );
   nand U43700 ( n42914,n42924,n42925 );
   nand U43701 ( n42925,n42926,n42655 );
   xor U43702 ( n42926,n42927,n42928 );
   nor U43703 ( n42924,n27897,n42929 );
   nor U43704 ( n42929,n42664,n42930 );
   nand U43705 ( n42930,n40365,n40364 );
   nand U43706 ( n40365,n42931,n42932 );
   nand U43707 ( n42932,n42814,n41808 );
   nor U43708 ( n42931,n42933,n42934 );
   nor U43709 ( n42934,n40317,n40359 );
   nor U43710 ( n42912,n42935,n42936 );
   nand U43711 ( n42936,n42937,n42938 );
   nand U43712 ( n42938,n42657,p2_ebx_reg_7_ );
   nand U43713 ( n42937,n28122,p2_reip_reg_7_ );
   nand U43714 ( n42935,n42939,n42940 );
   nand U43715 ( n42940,n28340,n39738 );
   nand U43716 ( n42939,n42682,p2_phyaddrpointer_reg_7_ );
   nor U43717 ( n42942,n42943,n42944 );
   nand U43718 ( n42944,n42945,n42946 );
   nand U43719 ( n42946,n42634,n42947 );
   not U43720 ( n42947,n38908 );
   nand U43721 ( n38908,n42948,n42949 );
   nand U43722 ( n42948,n42950,n42951 );
   nand U43723 ( n42951,n42919,n42952 );
   nand U43724 ( n42945,n28355,n38907 );
   not U43725 ( n38907,n41299 );
   nand U43726 ( n41299,n42953,n42954 );
   or U43727 ( n42953,n42955,n42956 );
   nand U43728 ( n42943,n42957,n42958 );
   nand U43729 ( n42958,n42959,n28331 );
   xor U43730 ( n42959,n40364,n40306 );
   nor U43731 ( n42957,n27897,n42960 );
   nor U43732 ( n42960,n42711,n42961 );
   nand U43733 ( n42961,n42962,n42963 );
   nand U43734 ( n42962,n39757,n42964 );
   nand U43735 ( n42964,n42928,n42927 );
   not U43736 ( n42927,n39738 );
   nor U43737 ( n42941,n42965,n42966 );
   nand U43738 ( n42966,n42967,n42968 );
   nand U43739 ( n42968,n42657,p2_ebx_reg_8_ );
   nand U43740 ( n42967,n28121,p2_reip_reg_8_ );
   nand U43741 ( n42965,n42969,n42970 );
   nand U43742 ( n42970,n28340,n39757 );
   nand U43743 ( n42969,n42682,p2_phyaddrpointer_reg_8_ );
   nor U43744 ( n42972,n42973,n42974 );
   nand U43745 ( n42974,n42975,n42976 );
   nand U43746 ( n42976,n42634,n38943 );
   not U43747 ( n38943,n39770 );
   xor U43748 ( n39770,n42977,n42978 );
   or U43749 ( n42975,n42744,n38938 );
   xor U43750 ( n38938,n42979,n42980 );
   nand U43751 ( n42973,n42981,n42982 );
   nand U43752 ( n42982,n42650,n40297 );
   not U43753 ( n40297,n40367 );
   nand U43754 ( n40367,n42983,n42984 );
   nand U43755 ( n42983,n42985,n42986 );
   nand U43756 ( n42986,n42987,n41825 );
   nor U43757 ( n42985,n28363,n42989 );
   nor U43758 ( n42989,n40306,n40364 );
   nor U43759 ( n42981,n27897,n42990 );
   nor U43760 ( n42990,n27898,n42991 );
   xor U43761 ( n42991,n42963,n42992 );
   nor U43762 ( n42971,n42993,n42994 );
   nand U43763 ( n42994,n42995,n42996 );
   nand U43764 ( n42996,n42657,p2_ebx_reg_9_ );
   nand U43765 ( n42995,n28121,p2_reip_reg_9_ );
   nand U43766 ( n42993,n42997,n42998 );
   nand U43767 ( n42998,n28340,n39775 );
   nand U43768 ( n42997,n42682,p2_phyaddrpointer_reg_9_ );
   nor U43769 ( n43000,n43001,n43002 );
   nand U43770 ( n43002,n43003,n43004 );
   nand U43771 ( n43004,n42634,n38962 );
   not U43772 ( n38962,n39790 );
   nand U43773 ( n39790,n43005,n43006 );
   nand U43774 ( n43005,n43007,n43008 );
   nand U43775 ( n43008,n42978,n43009 );
   nand U43776 ( n43003,n28355,n41657 );
   not U43777 ( n41657,n38957 );
   nand U43778 ( n38957,n43010,n43011 );
   nand U43779 ( n43010,n43012,n43013 );
   nand U43780 ( n43013,n42980,n43014 );
   nand U43781 ( n43001,n43015,n43016 );
   nand U43782 ( n43016,n42650,n40369 );
   xor U43783 ( n40369,n42984,n43017 );
   nor U43784 ( n43015,n27897,n43018 );
   nor U43785 ( n43018,n27898,n43019 );
   nand U43786 ( n43019,n43020,n43021 );
   nand U43787 ( n43020,n39795,n43022 );
   nand U43788 ( n43022,n43023,n42992 );
   not U43789 ( n42992,n39775 );
   nor U43790 ( n42999,n43024,n43025 );
   nand U43791 ( n43025,n43026,n43027 );
   nand U43792 ( n43027,n42657,p2_ebx_reg_10_ );
   nand U43793 ( n43026,n28122,p2_reip_reg_10_ );
   nand U43794 ( n43024,n43028,n43029 );
   nand U43795 ( n43029,n28340,n39795 );
   nand U43796 ( n43028,n42682,p2_phyaddrpointer_reg_10_ );
   nor U43797 ( n43031,n43032,n43033 );
   nand U43798 ( n43033,n43034,n43035 );
   nand U43799 ( n43035,n42634,n38991 );
   not U43800 ( n38991,n39809 );
   xor U43801 ( n39809,n43036,n43037 );
   nand U43802 ( n43034,n28355,n41646 );
   not U43803 ( n41646,n38986 );
   xor U43804 ( n38986,n43038,n43039 );
   nand U43805 ( n43032,n43040,n43041 );
   nand U43806 ( n43041,n42650,n40293 );
   not U43807 ( n40293,n40372 );
   nand U43808 ( n40372,n43042,n43043 );
   nand U43809 ( n43042,n43044,n43045 );
   nand U43810 ( n43045,n42987,n41839 );
   nor U43811 ( n43044,n28362,n43046 );
   nor U43812 ( n43046,n43017,n42984 );
   nor U43813 ( n43040,n42772,n43047 );
   nor U43814 ( n43047,n42711,n43048 );
   xor U43815 ( n43048,n43021,n43049 );
   nor U43816 ( n43030,n43050,n43051 );
   nand U43817 ( n43051,n43052,n43053 );
   nand U43818 ( n43053,n42657,p2_ebx_reg_11_ );
   nand U43819 ( n43052,n28121,p2_reip_reg_11_ );
   nand U43820 ( n43050,n43054,n43055 );
   nand U43821 ( n43055,n28340,n39814 );
   nand U43822 ( n43054,n42682,p2_phyaddrpointer_reg_11_ );
   nor U43823 ( n43057,n43058,n43059 );
   nand U43824 ( n43059,n43060,n43061 );
   nand U43825 ( n43061,n42650,n40289 );
   xor U43826 ( n40289,n43062,n43043 );
   nand U43827 ( n43060,n28355,n39003 );
   not U43828 ( n39003,n41316 );
   nand U43829 ( n41316,n43063,n43064 );
   nand U43830 ( n43063,n43065,n43066 );
   nand U43831 ( n43066,n43039,n43067 );
   nand U43832 ( n43058,n43068,n43069 );
   nand U43833 ( n43069,n42634,n39004 );
   not U43834 ( n39004,n39831 );
   nand U43835 ( n39831,n43070,n43071 );
   nand U43836 ( n43070,n43072,n43073 );
   nand U43837 ( n43073,n43037,n43074 );
   nor U43838 ( n43068,n42772,n43075 );
   nor U43839 ( n43075,n42711,n43076 );
   nand U43840 ( n43076,n43077,n43078 );
   nand U43841 ( n43077,n39836,n43079 );
   nand U43842 ( n43079,n43080,n43049 );
   not U43843 ( n43049,n39814 );
   nor U43844 ( n43056,n43081,n43082 );
   nand U43845 ( n43082,n43083,n43084 );
   nand U43846 ( n43084,n42657,p2_ebx_reg_12_ );
   nand U43847 ( n43083,n28121,p2_reip_reg_12_ );
   nand U43848 ( n43081,n43085,n43086 );
   nand U43849 ( n43086,n28340,n39836 );
   nand U43850 ( n43085,n42682,p2_phyaddrpointer_reg_12_ );
   nor U43851 ( n43088,n43089,n43090 );
   nand U43852 ( n43090,n43091,n43092 );
   nand U43853 ( n43092,n42650,n40286 );
   and U43854 ( n40286,n43093,n43094 );
   nand U43855 ( n43093,n43095,n43096 );
   nand U43856 ( n43096,n42987,n41857 );
   nor U43857 ( n43095,n28363,n43097 );
   nor U43858 ( n43097,n43062,n43043 );
   not U43859 ( n43043,n43098 );
   nand U43860 ( n43091,n28355,n39033 );
   not U43861 ( n39033,n41321 );
   xor U43862 ( n41321,n43099,n43100 );
   nand U43863 ( n43089,n43101,n43102 );
   nand U43864 ( n43102,n42634,n43103 );
   not U43865 ( n43103,n39034 );
   xor U43866 ( n39034,n43104,n43105 );
   nor U43867 ( n43101,n42772,n43106 );
   nor U43868 ( n43106,n27898,n43107 );
   xor U43869 ( n43107,n43078,n43108 );
   nor U43870 ( n43087,n43109,n43110 );
   nand U43871 ( n43110,n43111,n43112 );
   nand U43872 ( n43112,n42657,p2_ebx_reg_13_ );
   nand U43873 ( n43111,n42652,p2_reip_reg_13_ );
   nand U43874 ( n43109,n43113,n43114 );
   nand U43875 ( n43114,n28340,n39859 );
   nand U43876 ( n43113,n42682,p2_phyaddrpointer_reg_13_ );
   nor U43877 ( n43116,n43117,n43118 );
   nand U43878 ( n43118,n43119,n43120 );
   nand U43879 ( n43120,n42650,n40282 );
   xor U43880 ( n40282,n43094,n43121 );
   nand U43881 ( n43119,n28355,n39052 );
   not U43882 ( n39052,n41326 );
   nand U43883 ( n41326,n43122,n43123 );
   nand U43884 ( n43122,n43124,n43125 );
   nand U43885 ( n43125,n43100,n43126 );
   nand U43886 ( n43117,n43127,n43128 );
   nand U43887 ( n43128,n42634,n43129 );
   not U43888 ( n43129,n39053 );
   nand U43889 ( n39053,n43130,n43131 );
   nand U43890 ( n43130,n43132,n43133 );
   nand U43891 ( n43133,n43105,n43134 );
   nor U43892 ( n43127,n42772,n43135 );
   nor U43893 ( n43135,n42711,n43136 );
   nand U43894 ( n43136,n43137,n43138 );
   nand U43895 ( n43137,n39879,n43139 );
   nand U43896 ( n43139,n43140,n43108 );
   not U43897 ( n43108,n39859 );
   nor U43898 ( n43115,n43141,n43142 );
   nand U43899 ( n43142,n43143,n43144 );
   nand U43900 ( n43144,n42657,p2_ebx_reg_14_ );
   nand U43901 ( n43143,n28121,p2_reip_reg_14_ );
   nand U43902 ( n43141,n43145,n43146 );
   nand U43903 ( n43146,n28340,n39879 );
   nand U43904 ( n43145,n42682,p2_phyaddrpointer_reg_14_ );
   nor U43905 ( n43148,n43149,n43150 );
   nand U43906 ( n43150,n43151,n43152 );
   nand U43907 ( n43152,n28331,n40279 );
   and U43908 ( n40279,n43153,n43154 );
   nand U43909 ( n43153,n43155,n43156 );
   nand U43910 ( n43156,n42987,n41874 );
   nor U43911 ( n43155,n42988,n43157 );
   nor U43912 ( n43157,n43121,n43094 );
   nand U43913 ( n43151,n28355,n39080 );
   not U43914 ( n39080,n41331 );
   xor U43915 ( n41331,n43158,n43159 );
   nand U43916 ( n43149,n43160,n43161 );
   nand U43917 ( n43161,n42634,n39081 );
   not U43918 ( n39081,n39894 );
   xor U43919 ( n39894,n43162,n43163 );
   nor U43920 ( n43160,n42772,n43164 );
   nor U43921 ( n43164,n42711,n43165 );
   xor U43922 ( n43165,n43138,n43166 );
   nor U43923 ( n43147,n43167,n43168 );
   nand U43924 ( n43168,n43169,n43170 );
   nand U43925 ( n43170,n42657,p2_ebx_reg_15_ );
   nand U43926 ( n43169,n42652,p2_reip_reg_15_ );
   nand U43927 ( n43167,n43171,n43172 );
   nand U43928 ( n43172,n28340,n39899 );
   nand U43929 ( n43171,n42682,p2_phyaddrpointer_reg_15_ );
   nor U43930 ( n43174,n43175,n43176 );
   nand U43931 ( n43176,n43177,n43178 );
   nand U43932 ( n43178,n42650,n40275 );
   xor U43933 ( n40275,n43179,n43154 );
   nand U43934 ( n43177,n28355,n39100 );
   not U43935 ( n39100,n41628 );
   nand U43936 ( n41628,n43180,n43181 );
   nand U43937 ( n43180,n43182,n43183 );
   nand U43938 ( n43183,n43159,n43184 );
   nand U43939 ( n43175,n43185,n43186 );
   nand U43940 ( n43186,n28093,n43187 );
   not U43941 ( n43187,n39101 );
   nand U43942 ( n39101,n43188,n43189 );
   nand U43943 ( n43188,n43190,n43191 );
   nand U43944 ( n43191,n43163,n43192 );
   nor U43945 ( n43185,n42772,n43193 );
   nor U43946 ( n43193,n42711,n43194 );
   nand U43947 ( n43194,n43195,n43196 );
   nand U43948 ( n43195,n39924,n43197 );
   nand U43949 ( n43197,n43198,n43166 );
   not U43950 ( n43166,n39899 );
   nor U43951 ( n43173,n43199,n43200 );
   nand U43952 ( n43200,n43201,n43202 );
   nand U43953 ( n43202,n28360,p2_ebx_reg_16_ );
   nand U43954 ( n43201,n42652,p2_reip_reg_16_ );
   nand U43955 ( n43199,n43203,n43204 );
   nand U43956 ( n43204,n42722,n39924 );
   nand U43957 ( n43203,n42682,p2_phyaddrpointer_reg_16_ );
   nor U43958 ( n43206,n43207,n43208 );
   nand U43959 ( n43208,n43209,n43210 );
   nand U43960 ( n43210,n42650,n40272 );
   and U43961 ( n40272,n43211,n43212 );
   nand U43962 ( n43211,n43213,n43214 );
   nand U43963 ( n43214,n42987,n41889 );
   nor U43964 ( n43213,n28362,n43215 );
   nor U43965 ( n43215,n43179,n43154 );
   not U43966 ( n43154,n43216 );
   nand U43967 ( n43209,n42629,n39129 );
   not U43968 ( n39129,n41619 );
   xor U43969 ( n41619,n43217,n43218 );
   nand U43970 ( n43207,n43219,n43220 );
   nand U43971 ( n43220,n28093,n43221 );
   not U43972 ( n43221,n39130 );
   xor U43973 ( n39130,n43222,n43223 );
   nor U43974 ( n43219,n42772,n43224 );
   nor U43975 ( n43224,n42711,n43225 );
   xor U43976 ( n43225,n43196,n43226 );
   nor U43977 ( n43205,n43227,n43228 );
   nand U43978 ( n43228,n43229,n43230 );
   nand U43979 ( n43230,n28360,p2_ebx_reg_17_ );
   nand U43980 ( n43229,n28121,p2_reip_reg_17_ );
   nand U43981 ( n43227,n43231,n43232 );
   nand U43982 ( n43232,n42722,n39941 );
   nand U43983 ( n43231,n42682,p2_phyaddrpointer_reg_17_ );
   nor U43984 ( n43234,n43235,n43236 );
   nand U43985 ( n43236,n43237,n43238 );
   nand U43986 ( n43238,n42650,n40263 );
   xor U43987 ( n40263,n43212,n43239 );
   nand U43988 ( n43237,n42629,n39148 );
   not U43989 ( n39148,n41615 );
   nand U43990 ( n41615,n43240,n43241 );
   nand U43991 ( n43240,n43242,n43243 );
   nand U43992 ( n43243,n43218,n43244 );
   nand U43993 ( n43235,n43245,n43246 );
   nand U43994 ( n43246,n28093,n43247 );
   not U43995 ( n43247,n39149 );
   nand U43996 ( n39149,n43248,n43249 );
   nand U43997 ( n43248,n43250,n43251 );
   nand U43998 ( n43251,n43223,n43252 );
   nor U43999 ( n43245,n42772,n43253 );
   nor U44000 ( n43253,n42711,n43254 );
   nand U44001 ( n43254,n43255,n43256 );
   nand U44002 ( n43255,n39959,n43257 );
   nand U44003 ( n43257,n43258,n43226 );
   not U44004 ( n43226,n39941 );
   nor U44005 ( n43233,n43259,n43260 );
   nand U44006 ( n43260,n43261,n43262 );
   nand U44007 ( n43262,n28360,p2_ebx_reg_18_ );
   nand U44008 ( n43261,n42652,p2_reip_reg_18_ );
   nand U44009 ( n43259,n43263,n43264 );
   nand U44010 ( n43264,n42722,n39959 );
   nand U44011 ( n43263,n42682,p2_phyaddrpointer_reg_18_ );
   nor U44012 ( n43266,n43267,n43268 );
   nand U44013 ( n43268,n43269,n43270 );
   nand U44014 ( n43270,n28093,n43271 );
   not U44015 ( n43271,n39178 );
   xor U44016 ( n39178,n43272,n43273 );
   nand U44017 ( n43269,n42629,n39177 );
   not U44018 ( n39177,n41610 );
   xor U44019 ( n41610,n43274,n43275 );
   nand U44020 ( n43267,n43276,n43277 );
   nand U44021 ( n43277,n43278,n42655 );
   xor U44022 ( n43278,n39980,n43256 );
   nor U44023 ( n43276,n27897,n43279 );
   nor U44024 ( n43279,n42664,n43280 );
   nand U44025 ( n43280,n40266,n43281 );
   nand U44026 ( n40266,n43282,n43283 );
   nand U44027 ( n43283,n42987,n41904 );
   nor U44028 ( n43282,n28363,n43284 );
   nor U44029 ( n43284,n43239,n43212 );
   nor U44030 ( n42772,n36616,n42652 );
   nor U44031 ( n43265,n43285,n43286 );
   nand U44032 ( n43286,n43287,n43288 );
   nand U44033 ( n43288,n28360,p2_ebx_reg_19_ );
   nand U44034 ( n43287,n28122,p2_reip_reg_19_ );
   nand U44035 ( n43285,n43289,n43290 );
   nand U44036 ( n43290,n42722,n39980 );
   nand U44037 ( n43289,n28092,p2_phyaddrpointer_reg_19_ );
   nor U44038 ( n43292,n43293,n43294 );
   nand U44039 ( n43294,n43295,n43296 );
   nand U44040 ( n43296,n28093,n43297 );
   not U44041 ( n43297,n39197 );
   nand U44042 ( n39197,n43298,n43299 );
   nand U44043 ( n43298,n43300,n43301 );
   nand U44044 ( n43301,n43273,n43302 );
   nand U44045 ( n43295,n42629,n39196 );
   not U44046 ( n39196,n41606 );
   nand U44047 ( n41606,n43303,n43304 );
   nand U44048 ( n43303,n43305,n43306 );
   nand U44049 ( n43306,n43275,n43307 );
   nand U44050 ( n43293,n43308,n43309 );
   nand U44051 ( n43309,n43310,n42655 );
   nor U44052 ( n43310,n43311,n43312 );
   nor U44053 ( n43312,n43313,n43314 );
   nor U44054 ( n43313,n39980,n43256 );
   nand U44055 ( n43308,n40379,n28331 );
   xor U44056 ( n40379,n43315,n43281 );
   nor U44057 ( n43291,n43316,n43317 );
   nand U44058 ( n43317,n43318,n43319 );
   nand U44059 ( n43319,n28360,p2_ebx_reg_20_ );
   nand U44060 ( n43318,n28121,p2_reip_reg_20_ );
   nand U44061 ( n43316,n43320,n43321 );
   nand U44062 ( n43321,n42722,n39999 );
   nand U44063 ( n43320,n28092,p2_phyaddrpointer_reg_20_ );
   nor U44064 ( n43323,n43324,n43325 );
   nand U44065 ( n43325,n43326,n43327 );
   nand U44066 ( n43327,n28093,n43328 );
   not U44067 ( n43328,n39224 );
   xor U44068 ( n39224,n43329,n43330 );
   nand U44069 ( n43326,n42629,n39223 );
   not U44070 ( n39223,n41601 );
   xor U44071 ( n41601,n43331,n43332 );
   nand U44072 ( n43324,n43333,n43334 );
   nand U44073 ( n43334,n43335,n28331 );
   nor U44074 ( n43335,n40384,n40385 );
   not U44075 ( n40385,n40382 );
   nand U44076 ( n40382,n43336,n43337 );
   nand U44077 ( n43337,n42987,n41919 );
   nor U44078 ( n43336,n42988,n43338 );
   nor U44079 ( n43338,n43315,n43281 );
   not U44080 ( n43281,n40267 );
   nand U44081 ( n43333,n43339,n42655 );
   xor U44082 ( n43339,n40015,n43340 );
   nor U44083 ( n43322,n43341,n43342 );
   nand U44084 ( n43342,n43343,n43344 );
   nand U44085 ( n43344,n28360,p2_ebx_reg_21_ );
   nand U44086 ( n43343,n42652,p2_reip_reg_21_ );
   nand U44087 ( n43341,n43345,n43346 );
   nand U44088 ( n43346,n42722,n40015 );
   nand U44089 ( n43345,n28092,p2_phyaddrpointer_reg_21_ );
   nor U44090 ( n43348,n43349,n43350 );
   nand U44091 ( n43350,n43351,n43352 );
   nand U44092 ( n43352,n28093,n39242 );
   not U44093 ( n39242,n40038 );
   nand U44094 ( n40038,n43353,n43354 );
   nand U44095 ( n43353,n43355,n43356 );
   nand U44096 ( n43356,n43330,n43357 );
   nand U44097 ( n43351,n42629,n39241 );
   not U44098 ( n39241,n41597 );
   nand U44099 ( n41597,n43358,n43359 );
   nand U44100 ( n43358,n43360,n43361 );
   nand U44101 ( n43361,n43332,n43362 );
   nand U44102 ( n43349,n43363,n43364 );
   nand U44103 ( n43364,n43365,n42655 );
   nor U44104 ( n43365,n43366,n43367 );
   nor U44105 ( n43367,n43368,n43369 );
   nor U44106 ( n43368,n40015,n43340 );
   not U44107 ( n43340,n43311 );
   nand U44108 ( n43363,n40386,n28331 );
   xor U44109 ( n40386,n43370,n43371 );
   nor U44110 ( n43347,n43372,n43373 );
   nand U44111 ( n43373,n43374,n43375 );
   nand U44112 ( n43375,n28360,p2_ebx_reg_22_ );
   nand U44113 ( n43374,n28121,p2_reip_reg_22_ );
   nand U44114 ( n43372,n43376,n43377 );
   nand U44115 ( n43377,n42722,n40043 );
   nand U44116 ( n43376,n28092,p2_phyaddrpointer_reg_22_ );
   nor U44117 ( n43379,n43380,n43381 );
   nand U44118 ( n43381,n43382,n43383 );
   nand U44119 ( n43383,n42629,n39272 );
   not U44120 ( n39272,n41592 );
   xor U44121 ( n41592,n43384,n43385 );
   nand U44122 ( n43382,n28093,n43386 );
   not U44123 ( n43386,n39273 );
   xor U44124 ( n39273,n43387,n43388 );
   nand U44125 ( n43380,n43389,n43390 );
   nand U44126 ( n43390,n43391,n28331 );
   nor U44127 ( n43391,n40391,n40392 );
   not U44128 ( n40392,n40389 );
   nand U44129 ( n40389,n43392,n43393 );
   nand U44130 ( n43393,n42987,n41939 );
   nor U44131 ( n43392,n42988,n43394 );
   nor U44132 ( n43394,n43371,n43370 );
   nand U44133 ( n43389,n43395,n42655 );
   xor U44134 ( n43395,n40061,n43396 );
   nor U44135 ( n43378,n43397,n43398 );
   nand U44136 ( n43398,n43399,n43400 );
   nand U44137 ( n43400,n28360,p2_ebx_reg_23_ );
   nand U44138 ( n43399,n28122,p2_reip_reg_23_ );
   nand U44139 ( n43397,n43401,n43402 );
   nand U44140 ( n43402,n42722,n40061 );
   nand U44141 ( n43401,n28092,p2_phyaddrpointer_reg_23_ );
   nor U44142 ( n43404,n43405,n43406 );
   nand U44143 ( n43406,n43407,n43408 );
   nand U44144 ( n43408,n42629,n39291 );
   not U44145 ( n39291,n41589 );
   nand U44146 ( n41589,n43409,n43410 );
   nand U44147 ( n43409,n43411,n43412 );
   nand U44148 ( n43412,n43385,n43413 );
   nand U44149 ( n43407,n28093,n43414 );
   not U44150 ( n43414,n39292 );
   nand U44151 ( n39292,n43415,n43416 );
   nand U44152 ( n43415,n43417,n43418 );
   nand U44153 ( n43418,n43388,n43419 );
   nand U44154 ( n43405,n43420,n43421 );
   nand U44155 ( n43421,n43422,n42655 );
   nor U44156 ( n43422,n43423,n43424 );
   nor U44157 ( n43424,n43425,n43426 );
   nor U44158 ( n43425,n40061,n43396 );
   nand U44159 ( n43420,n40393,n28331 );
   xor U44160 ( n40393,n43427,n43428 );
   nor U44161 ( n43403,n43429,n43430 );
   nand U44162 ( n43430,n43431,n43432 );
   nand U44163 ( n43432,n28360,p2_ebx_reg_24_ );
   nand U44164 ( n43431,n28122,p2_reip_reg_24_ );
   nand U44165 ( n43429,n43433,n43434 );
   nand U44166 ( n43434,n42722,n40086 );
   nand U44167 ( n43433,n28092,p2_phyaddrpointer_reg_24_ );
   nor U44168 ( n43436,n43437,n43438 );
   nand U44169 ( n43438,n43439,n43440 );
   nand U44170 ( n43440,n28093,n39320 );
   not U44171 ( n39320,n40098 );
   xor U44172 ( n40098,n43441,n43442 );
   nand U44173 ( n43439,n42629,n39319 );
   not U44174 ( n39319,n41584 );
   xor U44175 ( n41584,n43443,n43444 );
   nand U44176 ( n43437,n43445,n43446 );
   nand U44177 ( n43446,n43447,n28331 );
   and U44178 ( n43447,n43448,n40243 );
   nand U44179 ( n40243,n43449,n43450 );
   nand U44180 ( n43450,n42987,n41963 );
   nor U44181 ( n43449,n28362,n43451 );
   nor U44182 ( n43451,n43427,n43428 );
   nand U44183 ( n43445,n43452,n42655 );
   xor U44184 ( n43452,n40103,n43453 );
   nor U44185 ( n43435,n43454,n43455 );
   nand U44186 ( n43455,n43456,n43457 );
   nand U44187 ( n43457,n28360,p2_ebx_reg_25_ );
   nand U44188 ( n43456,n28121,p2_reip_reg_25_ );
   nand U44189 ( n43454,n43458,n43459 );
   nand U44190 ( n43459,n42722,n40103 );
   nand U44191 ( n43458,n28092,p2_phyaddrpointer_reg_25_ );
   nor U44192 ( n43461,n43462,n43463 );
   nand U44193 ( n43463,n43464,n43465 );
   nand U44194 ( n43465,n42650,n40237 );
   not U44195 ( n40237,n40234 );
   xor U44196 ( n40234,n40244,n43466 );
   nand U44197 ( n43464,n42629,n39339 );
   not U44198 ( n39339,n41581 );
   nand U44199 ( n41581,n43467,n43468 );
   nand U44200 ( n43467,n43469,n43470 );
   nand U44201 ( n43470,n43444,n43471 );
   nand U44202 ( n43462,n43472,n43473 );
   nand U44203 ( n43473,n43474,n42655 );
   nor U44204 ( n43474,n43475,n43476 );
   nor U44205 ( n43476,n43477,n43478 );
   nor U44206 ( n43477,n40103,n43453 );
   nand U44207 ( n43472,n28093,n43479 );
   not U44208 ( n43479,n39340 );
   nand U44209 ( n39340,n43480,n43481 );
   nand U44210 ( n43480,n43482,n43483 );
   nand U44211 ( n43483,n43442,n43484 );
   nor U44212 ( n43460,n43485,n43486 );
   nand U44213 ( n43486,n43487,n43488 );
   nand U44214 ( n43488,n28360,p2_ebx_reg_26_ );
   nand U44215 ( n43487,n28122,p2_reip_reg_26_ );
   nand U44216 ( n43485,n43489,n43490 );
   nand U44217 ( n43490,n42722,n40128 );
   nand U44218 ( n43489,n28092,p2_phyaddrpointer_reg_26_ );
   nor U44219 ( n43492,n43493,n43494 );
   nand U44220 ( n43494,n43495,n43496 );
   nand U44221 ( n43496,n42629,n39368 );
   not U44222 ( n39368,n41576 );
   xor U44223 ( n41576,n43497,n43498 );
   nand U44224 ( n43495,n28093,n43499 );
   not U44225 ( n43499,n39369 );
   xor U44226 ( n39369,n43500,n43501 );
   nand U44227 ( n43493,n43502,n43503 );
   nand U44228 ( n43503,n43504,n42655 );
   xor U44229 ( n43504,n40144,n43505 );
   nand U44230 ( n43502,n42650,n40232 );
   and U44231 ( n40232,n43506,n43507 );
   nand U44232 ( n43506,n43508,n43509 );
   nand U44233 ( n43509,n42987,n41986 );
   nor U44234 ( n43508,n28363,n43510 );
   nor U44235 ( n43510,n43466,n43448 );
   nor U44236 ( n43491,n43511,n43512 );
   nand U44237 ( n43512,n43513,n43514 );
   nand U44238 ( n43514,n28360,p2_ebx_reg_27_ );
   nand U44239 ( n43513,n42652,p2_reip_reg_27_ );
   nand U44240 ( n43511,n43515,n43516 );
   nand U44241 ( n43516,n42722,n40144 );
   nand U44242 ( n43515,n28092,p2_phyaddrpointer_reg_27_ );
   nor U44243 ( n43518,n43519,n43520 );
   nand U44244 ( n43520,n43521,n43522 );
   nand U44245 ( n43522,n42650,n40228 );
   xor U44246 ( n40228,n43523,n43507 );
   nand U44247 ( n43521,n42629,n39386 );
   not U44248 ( n39386,n41573 );
   nand U44249 ( n41573,n43524,n43525 );
   nand U44250 ( n43524,n43526,n43527 );
   nand U44251 ( n43527,n43498,n43528 );
   nand U44252 ( n43519,n43529,n43530 );
   nand U44253 ( n43530,n43531,n42655 );
   nor U44254 ( n43531,n43532,n43533 );
   nor U44255 ( n43533,n43534,n43535 );
   nor U44256 ( n43534,n40144,n43505 );
   nand U44257 ( n43529,n28093,n39387 );
   not U44258 ( n39387,n40159 );
   nand U44259 ( n40159,n43536,n43537 );
   nand U44260 ( n43536,n43538,n43539 );
   nand U44261 ( n43539,n43501,n43540 );
   nor U44262 ( n43517,n43541,n43542 );
   nand U44263 ( n43542,n43543,n43544 );
   nand U44264 ( n43544,n28360,p2_ebx_reg_28_ );
   nand U44265 ( n43543,n42652,p2_reip_reg_28_ );
   nand U44266 ( n43541,n43545,n43546 );
   nand U44267 ( n43546,n42722,n40164 );
   nand U44268 ( n43545,n28092,p2_phyaddrpointer_reg_28_ );
   nor U44269 ( n43548,n43549,n43550 );
   nand U44270 ( n43550,n43551,n43552 );
   nand U44271 ( n43552,n42650,n40225 );
   nor U44272 ( n40225,n43553,n43554 );
   and U44273 ( n43553,n43555,n43556 );
   nand U44274 ( n43556,n28274,n42005 );
   nor U44275 ( n43555,n42988,n43557 );
   nor U44276 ( n43557,n43523,n43507 );
   nand U44277 ( n43551,n42629,n39406 );
   xor U44278 ( n39406,n43558,n43525 );
   nand U44279 ( n43549,n43559,n43560 );
   nand U44280 ( n43560,n43561,n42655 );
   nor U44281 ( n43561,n43562,n43563 );
   nor U44282 ( n43563,n43532,n43564 );
   nand U44283 ( n43559,n28093,n43565 );
   not U44284 ( n43565,n39407 );
   xor U44285 ( n39407,n43566,n43567 );
   nor U44286 ( n43547,n43568,n43569 );
   nand U44287 ( n43569,n43570,n43571 );
   nand U44288 ( n43571,n28360,p2_ebx_reg_29_ );
   nand U44289 ( n43570,n28121,p2_reip_reg_29_ );
   nand U44290 ( n43568,n43572,n43573 );
   nand U44291 ( n43573,n42722,n40183 );
   nand U44292 ( n43572,n28092,p2_phyaddrpointer_reg_29_ );
   nor U44293 ( n43575,n43576,n43577 );
   nand U44294 ( n43577,n43578,n43579 );
   nand U44295 ( n43579,n42650,n40218 );
   and U44296 ( n40218,n43580,n40401 );
   nand U44297 ( n43580,n43581,n43582 );
   nand U44298 ( n43582,n42987,n42615 );
   nor U44299 ( n43581,n28362,n43554 );
   not U44300 ( n42650,n42664 );
   nand U44301 ( n43578,n42629,n39432 );
   and U44302 ( n39432,n43583,n43584 );
   nand U44303 ( n43583,n43585,n43586 );
   nor U44304 ( n43586,n43587,n43588 );
   nor U44305 ( n43585,n43589,n43590 );
   nor U44306 ( n43590,n43558,n43525 );
   nand U44307 ( n43576,n43591,n43592 );
   nand U44308 ( n43592,n43593,n42655 );
   not U44309 ( n42655,n42711 );
   xor U44310 ( n43593,n40201,n43594 );
   nand U44311 ( n43591,n28093,n39424 );
   not U44312 ( n39424,n40191 );
   nand U44313 ( n40191,n43595,n43596 );
   nand U44314 ( n43595,n43597,n43598 );
   nor U44315 ( n43598,n43599,n43600 );
   nor U44316 ( n43597,n43601,n43602 );
   nor U44317 ( n43601,n43566,n43537 );
   nor U44318 ( n43574,n43603,n43604 );
   nand U44319 ( n43604,n43605,n43606 );
   nand U44320 ( n43606,n28360,p2_ebx_reg_30_ );
   nand U44321 ( n43605,n42652,p2_reip_reg_30_ );
   nand U44322 ( n43603,n43607,n43608 );
   nand U44323 ( n43608,n28340,n40201 );
   not U44324 ( n42722,n42639 );
   nand U44325 ( n42639,n43609,p2_state2_reg_1_ );
   nor U44326 ( n43609,n42652,n36764 );
   nand U44327 ( n43607,n28092,p2_phyaddrpointer_reg_30_ );
   nor U44328 ( n43611,n43612,n43613 );
   nand U44329 ( n43613,n43614,n43615 );
   nand U44330 ( n43615,n28093,n39461 );
   xor U44331 ( n39461,n43616,n43596 );
   nand U44332 ( n43596,n43617,n43567 );
   not U44333 ( n43567,n43537 );
   nand U44334 ( n43537,n43618,n43501 );
   not U44335 ( n43501,n43481 );
   nand U44336 ( n43481,n43619,n43442 );
   not U44337 ( n43442,n43416 );
   nand U44338 ( n43416,n43620,n43388 );
   not U44339 ( n43388,n43354 );
   nand U44340 ( n43354,n43621,n43330 );
   not U44341 ( n43330,n43299 );
   nand U44342 ( n43299,n43622,n43273 );
   not U44343 ( n43273,n43249 );
   nand U44344 ( n43249,n43623,n43223 );
   not U44345 ( n43223,n43189 );
   nand U44346 ( n43189,n43624,n43163 );
   not U44347 ( n43163,n43131 );
   nand U44348 ( n43131,n43625,n43105 );
   not U44349 ( n43105,n43071 );
   nand U44350 ( n43071,n43626,n43037 );
   not U44351 ( n43037,n43006 );
   nand U44352 ( n43006,n43627,n42978 );
   not U44353 ( n42978,n42949 );
   nand U44354 ( n42949,n43628,n42919 );
   not U44355 ( n42919,n42889 );
   nand U44356 ( n42889,n42891,n42890 );
   nand U44357 ( n42890,n43629,n43630 );
   nor U44358 ( n43630,n43631,n43632 );
   nor U44359 ( n43632,n28389,n41801 );
   nor U44360 ( n43631,n28410,n38877 );
   not U44361 ( n38877,p2_instaddrpointer_reg_6_ );
   nor U44362 ( n43629,n43635,n43636 );
   nor U44363 ( n43636,n28181,n39719 );
   nor U44364 ( n43635,n28384,n36935 );
   and U44365 ( n42891,n43638,n42768 );
   and U44366 ( n42768,n43639,n43640 );
   nand U44367 ( n43640,n42879,n43641 );
   or U44368 ( n43641,n42877,n42878 );
   and U44369 ( n42879,n43642,n43643 );
   nand U44370 ( n43643,p2_instqueuerd_addr_reg_3_,n43644 );
   nand U44371 ( n43642,n37216,p2_instqueuewr_addr_reg_3_ );
   nand U44372 ( n43639,n42878,n42877 );
   nand U44373 ( n42877,n43645,n43646 );
   nand U44374 ( n43646,n42854,n43647 );
   nand U44375 ( n43647,n42852,n42853 );
   and U44376 ( n42854,n43648,n43649 );
   nand U44377 ( n43649,n43650,n42842 );
   nand U44378 ( n42842,n43651,n43652 );
   nor U44379 ( n43652,n43653,n43654 );
   nor U44380 ( n43654,n37096,n43655 );
   nor U44381 ( n43653,n43656,n37120 );
   nor U44382 ( n43651,n43657,n43658 );
   nor U44383 ( n43657,n41756,n41037 );
   nand U44384 ( n43650,n42840,n42841 );
   or U44385 ( n43648,n42841,n42840 );
   and U44386 ( n42840,n43659,n43660 );
   nor U44387 ( n43660,n43661,n43662 );
   nor U44388 ( n43662,n41771,n28390 );
   nor U44389 ( n43661,n28409,n36758 );
   nor U44390 ( n43659,n43663,n43664 );
   nor U44391 ( n43664,n28178,n39621 );
   nor U44392 ( n43663,n28383,n36961 );
   nand U44393 ( n42841,n42864,n43665 );
   nand U44394 ( n43665,n43666,n42862 );
   nor U44395 ( n42862,n43667,n43668 );
   and U44396 ( n43668,n41750,n36650 );
   nor U44397 ( n43666,n42863,n43669 );
   nor U44398 ( n43669,n37336,n43655 );
   nor U44399 ( n42863,n37114,n43656 );
   nand U44400 ( n42864,n43670,n43671 );
   nor U44401 ( n43671,n43672,n43673 );
   nand U44402 ( n43673,n43674,n43675 );
   nand U44403 ( n43675,p2_reip_reg_0_,n43676 );
   nand U44404 ( n43674,p2_ebx_reg_0_,n43677 );
   nand U44405 ( n43672,n43678,n43679 );
   nand U44406 ( n43679,p2_instaddrpointer_reg_0_,n43680 );
   nor U44407 ( n43678,n43681,n43682 );
   not U44408 ( n43681,n43683 );
   nor U44409 ( n43670,n43684,n43685 );
   nand U44410 ( n43685,n43686,n43687 );
   nand U44411 ( n43687,n43688,p2_state2_reg_0_ );
   nor U44412 ( n43688,n39528,n43689 );
   nor U44413 ( n43689,n39573,n43690 );
   nor U44414 ( n39528,n36646,n41567 );
   nand U44415 ( n43684,n43655,n43691 );
   nand U44416 ( n43691,p2_phyaddrpointer_reg_0_,p2_state2_reg_1_ );
   not U44417 ( n43655,n37216 );
   nor U44418 ( n37216,p2_state2_reg_1_,p2_state2_reg_0_ );
   or U44419 ( n43645,n42852,n42853 );
   nand U44420 ( n42853,n43692,n43693 );
   nor U44421 ( n43693,n43694,n43695 );
   nor U44422 ( n43695,n28409,n38786 );
   not U44423 ( n38786,p2_instaddrpointer_reg_2_ );
   nor U44424 ( n43694,n43637,n36955 );
   nor U44425 ( n43692,n43696,n43697 );
   nor U44426 ( n43697,n28181,n39641 );
   nor U44427 ( n43696,n28389,n41776 );
   nand U44428 ( n42852,n43698,n43699 );
   nand U44429 ( n43699,p2_instqueuewr_addr_reg_2_,n36783 );
   nor U44430 ( n43698,p2_state2_reg_1_,n43700 );
   nor U44431 ( n43700,n43656,n37154 );
   not U44432 ( n43656,n43644 );
   nand U44433 ( n43644,n43701,n43702 );
   nor U44434 ( n43702,n43682,n43703 );
   nand U44435 ( n43703,n43683,n36655 );
   nand U44436 ( n43683,n43704,n39573 );
   nor U44437 ( n43704,n40863,n39519 );
   and U44438 ( n39519,n43705,n43706 );
   nor U44439 ( n43706,n43707,n43708 );
   nor U44440 ( n43708,n38649,n43709 );
   nor U44441 ( n43709,n43710,n43711 );
   nor U44442 ( n43711,n39515,n42814 );
   nor U44443 ( n43710,n38617,n38585 );
   nor U44444 ( n43707,n37113,n43712 );
   nor U44445 ( n43705,n39566,n43713 );
   nor U44446 ( n43713,n41567,n37130 );
   and U44447 ( n43682,n43714,n36644 );
   nor U44448 ( n43714,n43715,n36646 );
   nor U44449 ( n43715,n39558,n43716 );
   nand U44450 ( n43716,n37195,n38633 );
   nand U44451 ( n39558,n41332,n43717 );
   nor U44452 ( n41332,n41567,n39566 );
   nor U44453 ( n43701,n43718,n43719 );
   nand U44454 ( n43719,n43720,n43686 );
   nand U44455 ( n43686,n36644,n43721 );
   nand U44456 ( n43721,n37113,n39506 );
   not U44457 ( n39506,n37192 );
   nand U44458 ( n43720,n36650,n43690 );
   nand U44459 ( n43690,n43722,n43723 );
   nand U44460 ( n43723,n37130,n43724 );
   or U44461 ( n43722,n39520,n37130 );
   nor U44462 ( n39520,n43725,n39559 );
   nand U44463 ( n39559,n43717,n43726 );
   nand U44464 ( n43726,n41567,n37195 );
   nand U44465 ( n43717,n42814,n38585 );
   or U44466 ( n43725,n39566,n39553 );
   nor U44467 ( n39553,n41567,n37195 );
   nor U44468 ( n43718,n42814,n42289 );
   and U44469 ( n42878,n43727,n43728 );
   nor U44470 ( n43728,n43729,n43730 );
   nor U44471 ( n43730,n43634,n38805 );
   not U44472 ( n38805,p2_instaddrpointer_reg_3_ );
   nor U44473 ( n43729,n43637,n36950 );
   nor U44474 ( n43727,n43731,n43732 );
   nor U44475 ( n43732,n28180,n39661 );
   nor U44476 ( n43731,n43633,n41781 );
   not U44477 ( n41781,p2_ebx_reg_3_ );
   nor U44478 ( n43638,n42767,n42804 );
   and U44479 ( n42804,n43733,n43734 );
   nor U44480 ( n43734,n43735,n43736 );
   nor U44481 ( n43736,n28390,n41793 );
   not U44482 ( n41793,p2_ebx_reg_5_ );
   nor U44483 ( n43735,n28409,n38851 );
   not U44484 ( n38851,p2_instaddrpointer_reg_5_ );
   nor U44485 ( n43733,n43737,n43738 );
   nor U44486 ( n43738,n28180,n39700 );
   nor U44487 ( n43737,n28383,n36940 );
   not U44488 ( n42767,n42806 );
   nand U44489 ( n42806,n43739,n43740 );
   nor U44490 ( n43740,n43741,n43742 );
   nor U44491 ( n43742,n28410,n38830 );
   not U44492 ( n38830,p2_instaddrpointer_reg_4_ );
   nor U44493 ( n43741,n28384,n36945 );
   nor U44494 ( n43739,n43743,n43744 );
   nor U44495 ( n43744,n28178,n39680 );
   nor U44496 ( n43743,n28389,n41787 );
   nor U44497 ( n43628,n42918,n42950 );
   and U44498 ( n42950,n43745,n43746 );
   nor U44499 ( n43746,n43747,n43748 );
   nor U44500 ( n43748,n28390,n41815 );
   nor U44501 ( n43747,n43634,n38925 );
   nor U44502 ( n43745,n43749,n43750 );
   nor U44503 ( n43750,n28179,n39758 );
   nor U44504 ( n43749,n43637,n36925 );
   not U44505 ( n42918,n42952 );
   nand U44506 ( n42952,n43751,n43752 );
   nor U44507 ( n43752,n43753,n43754 );
   nor U44508 ( n43754,n28389,n41808 );
   not U44509 ( n41808,p2_ebx_reg_7_ );
   nor U44510 ( n43753,n43634,n38899 );
   not U44511 ( n38899,p2_instaddrpointer_reg_7_ );
   nor U44512 ( n43751,n43755,n43756 );
   nor U44513 ( n43756,n28179,n39739 );
   nor U44514 ( n43755,n43637,n36930 );
   nor U44515 ( n43627,n42977,n43007 );
   and U44516 ( n43007,n43757,n43758 );
   nor U44517 ( n43758,n43759,n43760 );
   nor U44518 ( n43760,n43633,n41832 );
   nor U44519 ( n43759,n28409,n38974 );
   nor U44520 ( n43757,n43761,n43762 );
   nor U44521 ( n43762,n28181,n39796 );
   nor U44522 ( n43761,n28383,n36915 );
   not U44523 ( n42977,n43009 );
   nand U44524 ( n43009,n43763,n43764 );
   nor U44525 ( n43764,n43765,n43766 );
   nor U44526 ( n43766,n28390,n41825 );
   nor U44527 ( n43765,n28410,n38948 );
   nor U44528 ( n43763,n43767,n43768 );
   nor U44529 ( n43768,n28181,n39776 );
   nor U44530 ( n43767,n28384,n36920 );
   nor U44531 ( n43626,n43036,n43072 );
   and U44532 ( n43072,n43769,n43770 );
   nor U44533 ( n43770,n43771,n43772 );
   nor U44534 ( n43772,n28389,n41846 );
   nor U44535 ( n43771,n43634,n39022 );
   nor U44536 ( n43769,n43773,n43774 );
   nor U44537 ( n43774,n28178,n39837 );
   nor U44538 ( n43773,n43637,n36905 );
   not U44539 ( n43036,n43074 );
   nand U44540 ( n43074,n43775,n43776 );
   nor U44541 ( n43776,n43777,n43778 );
   nor U44542 ( n43778,n43633,n41839 );
   nor U44543 ( n43777,n28409,n38996 );
   nor U44544 ( n43775,n43779,n43780 );
   nor U44545 ( n43780,n28179,n39815 );
   nor U44546 ( n43779,n28383,n36910 );
   nor U44547 ( n43625,n43104,n43132 );
   and U44548 ( n43132,n43781,n43782 );
   nor U44549 ( n43782,n43783,n43784 );
   nor U44550 ( n43784,n28389,n41865 );
   nor U44551 ( n43783,n28410,n39070 );
   nor U44552 ( n43781,n43785,n43786 );
   nor U44553 ( n43786,n28179,n39880 );
   nor U44554 ( n43785,n28384,n36895 );
   not U44555 ( n43104,n43134 );
   nand U44556 ( n43134,n43787,n43788 );
   nor U44557 ( n43788,n43789,n43790 );
   nor U44558 ( n43790,n28390,n41857 );
   nor U44559 ( n43789,n28410,n39043 );
   nor U44560 ( n43787,n43791,n43792 );
   nor U44561 ( n43792,n28180,n39860 );
   nor U44562 ( n43791,n28383,n36900 );
   nor U44563 ( n43624,n43162,n43190 );
   and U44564 ( n43190,n43793,n43794 );
   nor U44565 ( n43794,n43795,n43796 );
   nor U44566 ( n43796,n28390,n41883 );
   nor U44567 ( n43795,n28409,n39118 );
   nor U44568 ( n43793,n43797,n43798 );
   nor U44569 ( n43798,n28180,n39925 );
   nor U44570 ( n43797,n43637,n36885 );
   not U44571 ( n43162,n43192 );
   nand U44572 ( n43192,n43799,n43800 );
   nor U44573 ( n43800,n43801,n43802 );
   nor U44574 ( n43802,n28390,n41874 );
   nor U44575 ( n43801,n28410,n39092 );
   nor U44576 ( n43799,n43803,n43804 );
   nor U44577 ( n43804,n28178,n39900 );
   nor U44578 ( n43803,n28384,n36890 );
   nor U44579 ( n43623,n43222,n43250 );
   and U44580 ( n43250,n43805,n43806 );
   nor U44581 ( n43806,n43807,n43808 );
   nor U44582 ( n43808,n43633,n41898 );
   nor U44583 ( n43807,n43634,n39166 );
   nor U44584 ( n43805,n43809,n43810 );
   nor U44585 ( n43810,n28179,n39960 );
   nor U44586 ( n43809,n28383,n36875 );
   not U44587 ( n43222,n43252 );
   nand U44588 ( n43252,n43811,n43812 );
   nor U44589 ( n43812,n43813,n43814 );
   nor U44590 ( n43814,n28389,n41889 );
   nor U44591 ( n43813,n43634,n39140 );
   nor U44592 ( n43811,n43815,n43816 );
   nor U44593 ( n43816,n28181,n39942 );
   nor U44594 ( n43815,n43637,n36880 );
   nor U44595 ( n43622,n43272,n43300 );
   and U44596 ( n43300,n43817,n43818 );
   nor U44597 ( n43818,n43819,n43820 );
   nor U44598 ( n43820,n43633,n41913 );
   nor U44599 ( n43819,n28410,n39212 );
   nor U44600 ( n43817,n43821,n43822 );
   nor U44601 ( n43822,n28181,n40000 );
   nor U44602 ( n43821,n28384,n36865 );
   not U44603 ( n43272,n43302 );
   nand U44604 ( n43302,n43823,n43824 );
   nor U44605 ( n43824,n43825,n43826 );
   nor U44606 ( n43826,n28390,n41904 );
   nor U44607 ( n43825,n28409,n39188 );
   nor U44608 ( n43823,n43827,n43828 );
   nor U44609 ( n43828,n28178,n39981 );
   nor U44610 ( n43827,n43637,n36870 );
   nor U44611 ( n43621,n43329,n43355 );
   and U44612 ( n43355,n43829,n43830 );
   nor U44613 ( n43830,n43831,n43832 );
   nor U44614 ( n43832,n43633,n41928 );
   nor U44615 ( n43831,n43634,n39261 );
   nor U44616 ( n43829,n43833,n43834 );
   nor U44617 ( n43834,n28178,n40044 );
   nor U44618 ( n43833,n28383,n36855 );
   not U44619 ( n43329,n43357 );
   nand U44620 ( n43357,n43835,n43836 );
   nor U44621 ( n43836,n43837,n43838 );
   nor U44622 ( n43838,n28389,n41919 );
   nor U44623 ( n43837,n28410,n39234 );
   nor U44624 ( n43835,n43839,n43840 );
   nor U44625 ( n43840,n28180,n40016 );
   nor U44626 ( n43839,n28384,n36860 );
   nor U44627 ( n43620,n43387,n43417 );
   and U44628 ( n43417,n43841,n43842 );
   nor U44629 ( n43842,n43843,n43844 );
   nor U44630 ( n43844,n43633,n41952 );
   nor U44631 ( n43843,n43634,n39309 );
   nor U44632 ( n43841,n43845,n43846 );
   nor U44633 ( n43846,n28180,n40087 );
   nor U44634 ( n43845,n43637,n36845 );
   not U44635 ( n43387,n43419 );
   nand U44636 ( n43419,n43847,n43848 );
   nor U44637 ( n43848,n43849,n43850 );
   nor U44638 ( n43850,n28390,n41939 );
   nor U44639 ( n43849,n28409,n39283 );
   nor U44640 ( n43847,n43851,n43852 );
   nor U44641 ( n43852,n28180,n40062 );
   nor U44642 ( n43851,n28383,n36850 );
   nor U44643 ( n43619,n43441,n43482 );
   and U44644 ( n43482,n43853,n43854 );
   nor U44645 ( n43854,n43855,n43856 );
   nor U44646 ( n43856,n28389,n41975 );
   nor U44647 ( n43855,n43634,n39357 );
   nor U44648 ( n43853,n43857,n43858 );
   nor U44649 ( n43858,n28179,n40129 );
   nor U44650 ( n43857,n28384,n36835 );
   not U44651 ( n43441,n43484 );
   nand U44652 ( n43484,n43859,n43860 );
   nor U44653 ( n43860,n43861,n43862 );
   nor U44654 ( n43862,n43633,n41963 );
   nor U44655 ( n43861,n28410,n39331 );
   nor U44656 ( n43859,n43863,n43864 );
   nor U44657 ( n43864,n28180,n40104 );
   nor U44658 ( n43863,n43637,n36840 );
   nor U44659 ( n43618,n43500,n43538 );
   and U44660 ( n43538,n43865,n43866 );
   nor U44661 ( n43866,n43867,n43868 );
   nor U44662 ( n43868,n28390,n41998 );
   nor U44663 ( n43867,n28409,n39396 );
   nor U44664 ( n43865,n43869,n43870 );
   nor U44665 ( n43870,n28181,n40165 );
   nor U44666 ( n43869,n28383,n36825 );
   not U44667 ( n43500,n43540 );
   nand U44668 ( n43540,n43871,n43872 );
   nor U44669 ( n43872,n43873,n43874 );
   nor U44670 ( n43874,n28389,n41986 );
   nor U44671 ( n43873,n43634,n39379 );
   nor U44672 ( n43871,n43875,n43876 );
   nor U44673 ( n43876,n28179,n40145 );
   nor U44674 ( n43875,n28384,n36830 );
   nor U44675 ( n43617,n43566,n43877 );
   nor U44676 ( n43877,n43602,n43878 );
   or U44677 ( n43878,n43600,n43599 );
   nor U44678 ( n43599,n39435,n28409 );
   nor U44679 ( n43600,n42615,n43633 );
   not U44680 ( n42615,p2_ebx_reg_30_ );
   nand U44681 ( n43602,n43879,n43880 );
   nand U44682 ( n43880,p2_reip_reg_30_,n43676 );
   nand U44683 ( n43879,p2_phyaddrpointer_reg_30_,p2_state2_reg_1_ );
   and U44684 ( n43566,n43881,n43882 );
   nor U44685 ( n43882,n43883,n43884 );
   nor U44686 ( n43884,n43633,n42005 );
   not U44687 ( n43633,n43677 );
   nor U44688 ( n43883,n28409,n39416 );
   nor U44689 ( n43881,n43885,n43886 );
   nor U44690 ( n43886,n28179,n40184 );
   nor U44691 ( n43885,n28383,n36820 );
   not U44692 ( n43637,n43676 );
   nor U44693 ( n43616,n43887,n43888 );
   nand U44694 ( n43888,n43889,n43890 );
   nand U44695 ( n43890,p2_reip_reg_31_,n43676 );
   nor U44696 ( n43676,n43891,n41756 );
   nand U44697 ( n43889,p2_phyaddrpointer_reg_31_,p2_state2_reg_1_ );
   nand U44698 ( n43887,n43892,n43893 );
   nand U44699 ( n43893,p2_instaddrpointer_reg_31_,n43680 );
   not U44700 ( n43680,n28410 );
   nor U44701 ( n43634,n43894,n43658 );
   nand U44702 ( n43658,n41202,n43895 );
   nand U44703 ( n43895,n43896,n43897 );
   nor U44704 ( n43897,n40863,n39515 );
   nor U44705 ( n43896,n38680,n39466 );
   or U44706 ( n43894,n43667,n43898 );
   and U44707 ( n43898,p2_state2_reg_0_,n37068 );
   nor U44708 ( n37068,n37203,n41756 );
   and U44709 ( n43667,n43899,n43900 );
   nor U44710 ( n43900,n37195,n38680 );
   not U44711 ( n37195,n38617 );
   nor U44712 ( n43899,n39466,n42289 );
   not U44713 ( n42289,n42015 );
   nor U44714 ( n42015,n38585,n40863 );
   nand U44715 ( n39466,n43901,n43902 );
   nor U44716 ( n43902,n39566,n38649 );
   nor U44717 ( n43901,n38601,n38633 );
   nand U44718 ( n43892,p2_ebx_reg_31_,n43677 );
   nor U44719 ( n43677,n39507,n36783 );
   nand U44720 ( n39507,n41750,n39455 );
   and U44721 ( n41750,n43903,n39529 );
   not U44722 ( n39529,n43724 );
   nand U44723 ( n43724,n43904,n43905 );
   nor U44724 ( n43905,n39515,n38617 );
   nor U44725 ( n43904,n38601,n38565 );
   nor U44726 ( n43903,n38649,n38633 );
   and U44727 ( n42634,n43906,n42826 );
   nor U44728 ( n43906,n37132,n43907 );
   nand U44729 ( n43614,n28092,p2_phyaddrpointer_reg_31_ );
   nor U44730 ( n42682,n38681,n28121 );
   nand U44731 ( n43612,n43908,n43909 );
   nand U44732 ( n43909,n43910,n43562 );
   not U44733 ( n43562,n43594 );
   nand U44734 ( n43594,n43532,n43564 );
   not U44735 ( n43564,n40183 );
   xor U44736 ( n40183,p2_phyaddrpointer_reg_29_,n43911 );
   and U44737 ( n43532,n43912,n43475 );
   not U44738 ( n43475,n43505 );
   nand U44739 ( n43505,n43913,n43423 );
   not U44740 ( n43423,n43453 );
   nand U44741 ( n43453,n43914,n43366 );
   not U44742 ( n43366,n43396 );
   nand U44743 ( n43396,n43915,n43311 );
   nor U44744 ( n43311,n43916,n43256 );
   nand U44745 ( n43256,n43917,n43258 );
   not U44746 ( n43258,n43196 );
   nand U44747 ( n43196,n43918,n43198 );
   not U44748 ( n43198,n43138 );
   nand U44749 ( n43138,n43919,n43140 );
   not U44750 ( n43140,n43078 );
   nand U44751 ( n43078,n43920,n43080 );
   not U44752 ( n43080,n43021 );
   nand U44753 ( n43021,n43921,n43023 );
   not U44754 ( n43023,n42963 );
   nand U44755 ( n42963,n43922,n42928 );
   not U44756 ( n42928,n42903 );
   nand U44757 ( n42903,n43923,n42905 );
   not U44758 ( n42905,n42776 );
   nand U44759 ( n42776,n43924,n42750 );
   not U44760 ( n42750,n42714 );
   nand U44761 ( n42714,n43925,n36759 );
   nand U44762 ( n36759,n43926,n43927 );
   nand U44763 ( n43927,p2_phyaddrpointer_reg_1_,n27895 );
   nand U44764 ( n43926,p2_state2_reg_0_,n36758 );
   nor U44765 ( n43925,n39639,n42656 );
   not U44766 ( n42656,n36763 );
   nand U44767 ( n36763,n43928,n43929 );
   or U44768 ( n43929,p2_phyaddrpointer_reg_0_,p2_state2_reg_0_ );
   nand U44769 ( n43928,p2_state2_reg_0_,n36762 );
   and U44770 ( n39639,n43930,n43931 );
   nand U44771 ( n43931,n39621,n39641 );
   not U44772 ( n39641,p2_phyaddrpointer_reg_2_ );
   not U44773 ( n39621,p2_phyaddrpointer_reg_1_ );
   nor U44774 ( n43924,n39679,n39660 );
   xor U44775 ( n39660,n39661,n43930 );
   not U44776 ( n39679,n42786 );
   nand U44777 ( n42786,n43932,n43933 );
   nand U44778 ( n43932,n39680,n43934 );
   or U44779 ( n43934,n43930,n39661 );
   not U44780 ( n39680,p2_phyaddrpointer_reg_4_ );
   nor U44781 ( n43923,n39718,n39699 );
   xor U44782 ( n39699,n39700,n43933 );
   and U44783 ( n39718,n43935,n43936 );
   nand U44784 ( n43935,n39719,n43937 );
   or U44785 ( n43937,n39700,n43933 );
   not U44786 ( n39719,p2_phyaddrpointer_reg_6_ );
   nor U44787 ( n43922,n39757,n39738 );
   xor U44788 ( n39738,n39739,n43936 );
   and U44789 ( n39757,n43938,n43939 );
   nand U44790 ( n43938,n39758,n43940 );
   or U44791 ( n43940,n39739,n43936 );
   not U44792 ( n39758,p2_phyaddrpointer_reg_8_ );
   nor U44793 ( n43921,n39795,n39775 );
   xor U44794 ( n39775,n39776,n43939 );
   and U44795 ( n39795,n43941,n43942 );
   nand U44796 ( n43941,n39796,n43943 );
   or U44797 ( n43943,n39776,n43939 );
   not U44798 ( n39776,p2_phyaddrpointer_reg_9_ );
   nor U44799 ( n43920,n39836,n39814 );
   xor U44800 ( n39814,n39815,n43942 );
   and U44801 ( n39836,n43944,n43945 );
   nand U44802 ( n43944,n39837,n43946 );
   or U44803 ( n43946,n39815,n43942 );
   not U44804 ( n39837,p2_phyaddrpointer_reg_12_ );
   nor U44805 ( n43919,n39879,n39859 );
   xor U44806 ( n39859,n39860,n43945 );
   and U44807 ( n39879,n43947,n43948 );
   nand U44808 ( n43947,n39880,n43949 );
   or U44809 ( n43949,n39860,n43945 );
   not U44810 ( n39880,p2_phyaddrpointer_reg_14_ );
   nor U44811 ( n43918,n39924,n39899 );
   xor U44812 ( n39899,n39900,n43948 );
   and U44813 ( n39924,n43950,n43951 );
   nand U44814 ( n43950,n39925,n43952 );
   or U44815 ( n43952,n39900,n43948 );
   not U44816 ( n39925,p2_phyaddrpointer_reg_16_ );
   nor U44817 ( n43917,n39959,n39941 );
   xor U44818 ( n39941,n39942,n43951 );
   and U44819 ( n39959,n43953,n43954 );
   nand U44820 ( n43953,n39960,n43955 );
   or U44821 ( n43955,n39942,n43951 );
   not U44822 ( n39960,p2_phyaddrpointer_reg_18_ );
   or U44823 ( n43916,n39999,n39980 );
   xor U44824 ( n39980,n39981,n43954 );
   not U44825 ( n39999,n43314 );
   nand U44826 ( n43314,n43956,n43957 );
   nand U44827 ( n43957,n43958,n40000 );
   nor U44828 ( n43915,n40043,n40015 );
   xor U44829 ( n40015,n40016,n43956 );
   not U44830 ( n40043,n43369 );
   nand U44831 ( n43369,n43959,n43960 );
   nand U44832 ( n43960,n43961,n40044 );
   nor U44833 ( n43914,n40086,n40061 );
   xor U44834 ( n40061,n40062,n43959 );
   not U44835 ( n40086,n43426 );
   nand U44836 ( n43426,n43962,n43963 );
   nand U44837 ( n43963,n43964,n40087 );
   nor U44838 ( n43913,n40128,n40103 );
   xor U44839 ( n40103,n40104,n43962 );
   not U44840 ( n40128,n43478 );
   nand U44841 ( n43478,n43965,n43966 );
   nand U44842 ( n43966,n43967,n40129 );
   nor U44843 ( n43912,n40164,n40144 );
   xor U44844 ( n40144,n40145,n43965 );
   not U44845 ( n40164,n43535 );
   nand U44846 ( n43535,n43968,n43969 );
   nand U44847 ( n43969,n43970,n40165 );
   nor U44848 ( n43910,n40201,n27898 );
   nand U44849 ( n42711,n43971,n36764 );
   not U44850 ( n36764,n36757 );
   nand U44851 ( n36757,n43972,n43973 );
   nand U44852 ( n43973,p2_state2_reg_0_,n39482 );
   not U44853 ( n39482,p2_instaddrpointer_reg_31_ );
   nand U44854 ( n43972,n43974,n27895 );
   xor U44855 ( n43974,p2_phyaddrpointer_reg_31_,n40872 );
   nor U44856 ( n43971,n28121,n28180 );
   and U44857 ( n40201,n43975,n40872 );
   nand U44858 ( n40872,n43976,p2_phyaddrpointer_reg_30_ );
   nor U44859 ( n43976,n43968,n40184 );
   not U44860 ( n40184,p2_phyaddrpointer_reg_29_ );
   not U44861 ( n43968,n43911 );
   nand U44862 ( n43975,n40202,n43977 );
   nand U44863 ( n43977,p2_phyaddrpointer_reg_29_,n43911 );
   nor U44864 ( n43911,n40165,n43970 );
   or U44865 ( n43970,n40145,n43965 );
   or U44866 ( n43965,n40129,n43967 );
   or U44867 ( n43967,n40104,n43962 );
   or U44868 ( n43962,n40087,n43964 );
   or U44869 ( n43964,n40062,n43959 );
   or U44870 ( n43959,n40044,n43961 );
   or U44871 ( n43961,n40016,n43956 );
   or U44872 ( n43956,n40000,n43958 );
   or U44873 ( n43958,n39981,n43954 );
   nand U44874 ( n43954,n43978,p2_phyaddrpointer_reg_18_ );
   nor U44875 ( n43978,n43951,n39942 );
   not U44876 ( n39942,p2_phyaddrpointer_reg_17_ );
   nand U44877 ( n43951,n43979,p2_phyaddrpointer_reg_16_ );
   nor U44878 ( n43979,n43948,n39900 );
   not U44879 ( n39900,p2_phyaddrpointer_reg_15_ );
   nand U44880 ( n43948,n43980,p2_phyaddrpointer_reg_14_ );
   nor U44881 ( n43980,n43945,n39860 );
   not U44882 ( n39860,p2_phyaddrpointer_reg_13_ );
   nand U44883 ( n43945,n43981,p2_phyaddrpointer_reg_12_ );
   nor U44884 ( n43981,n43942,n39815 );
   not U44885 ( n39815,p2_phyaddrpointer_reg_11_ );
   nand U44886 ( n43942,n43982,p2_phyaddrpointer_reg_9_ );
   nor U44887 ( n43982,n43939,n39796 );
   not U44888 ( n39796,p2_phyaddrpointer_reg_10_ );
   nand U44889 ( n43939,n43983,p2_phyaddrpointer_reg_8_ );
   nor U44890 ( n43983,n43936,n39739 );
   not U44891 ( n39739,p2_phyaddrpointer_reg_7_ );
   nand U44892 ( n43936,n43984,p2_phyaddrpointer_reg_6_ );
   nor U44893 ( n43984,n43933,n39700 );
   not U44894 ( n39700,p2_phyaddrpointer_reg_5_ );
   nand U44895 ( n43933,n43985,p2_phyaddrpointer_reg_4_ );
   nor U44896 ( n43985,n39661,n43930 );
   nand U44897 ( n43930,p2_phyaddrpointer_reg_2_,p2_phyaddrpointer_reg_1_ );
   not U44898 ( n39661,p2_phyaddrpointer_reg_3_ );
   not U44899 ( n39981,p2_phyaddrpointer_reg_19_ );
   not U44900 ( n40000,p2_phyaddrpointer_reg_20_ );
   not U44901 ( n40016,p2_phyaddrpointer_reg_21_ );
   not U44902 ( n40044,p2_phyaddrpointer_reg_22_ );
   not U44903 ( n40062,p2_phyaddrpointer_reg_23_ );
   not U44904 ( n40087,p2_phyaddrpointer_reg_24_ );
   not U44905 ( n40104,p2_phyaddrpointer_reg_25_ );
   not U44906 ( n40129,p2_phyaddrpointer_reg_26_ );
   not U44907 ( n40145,p2_phyaddrpointer_reg_27_ );
   not U44908 ( n40165,p2_phyaddrpointer_reg_28_ );
   not U44909 ( n40202,p2_phyaddrpointer_reg_30_ );
   or U44910 ( n43908,n42664,n40401 );
   nand U44911 ( n40401,n43554,n43986 );
   nand U44912 ( n43986,p2_ebx_reg_30_,n40399 );
   nor U44913 ( n43554,n43987,n43507 );
   nand U44914 ( n43507,n43988,n40244 );
   not U44915 ( n40244,n43448 );
   nand U44916 ( n43448,n43989,n40391 );
   not U44917 ( n40391,n43428 );
   nand U44918 ( n43428,n43990,n40384 );
   not U44919 ( n40384,n43370 );
   nand U44920 ( n43370,n43991,n40267 );
   nor U44921 ( n40267,n43992,n43212 );
   nand U44922 ( n43212,n43993,n43216 );
   nor U44923 ( n43216,n43994,n43094 );
   nand U44924 ( n43094,n43995,n43098 );
   nor U44925 ( n43098,n43996,n42984 );
   nand U44926 ( n42984,n43997,n40307 );
   not U44927 ( n40307,n40364 );
   nand U44928 ( n40364,n43998,n40318 );
   not U44929 ( n40318,n40359 );
   nand U44930 ( n40359,n43999,n40329 );
   nor U44931 ( n40329,n40352,n42741 );
   nand U44932 ( n42741,n44000,n44001 );
   nand U44933 ( n44001,n44002,n28239 );
   nand U44934 ( n44000,p2_ebx_reg_3_,n42814 );
   or U44935 ( n40352,n40355,n40354 );
   and U44936 ( n40354,n44003,n44004 );
   nand U44937 ( n44004,n42814,n41776 );
   not U44938 ( n41776,p2_ebx_reg_2_ );
   nand U44939 ( n44003,n44005,n28239 );
   not U44940 ( n40355,n42710 );
   nor U44941 ( n42710,n44006,n42651 );
   nor U44942 ( n42651,n41766,n38601 );
   not U44943 ( n41766,p2_ebx_reg_0_ );
   or U44944 ( n44006,n44007,n44008 );
   nor U44945 ( n44008,n41771,n38601 );
   not U44946 ( n41771,p2_ebx_reg_1_ );
   nor U44947 ( n44007,n42814,n44009 );
   nor U44948 ( n43999,n44010,n40328 );
   and U44949 ( n40328,n44011,n44012 );
   nand U44950 ( n44012,n42814,n41787 );
   not U44951 ( n41787,p2_ebx_reg_4_ );
   nand U44952 ( n44011,n44013,n28239 );
   nor U44953 ( n44010,n42815,n44014 );
   nor U44954 ( n44014,p2_ebx_reg_5_,n38601 );
   and U44955 ( n42815,n44015,n44016 );
   or U44956 ( n44016,n40749,n37132 );
   nor U44957 ( n43998,n44017,n40317 );
   not U44958 ( n40317,n42899 );
   nand U44959 ( n42899,n44018,n44019 );
   nand U44960 ( n44019,n42814,n41801 );
   not U44961 ( n41801,p2_ebx_reg_6_ );
   nand U44962 ( n44018,n44020,n28239 );
   nor U44963 ( n44017,n42933,n44021 );
   nor U44964 ( n44021,p2_ebx_reg_7_,n38601 );
   and U44965 ( n42933,n44015,n40229 );
   nor U44966 ( n44015,n44022,n42814 );
   nor U44967 ( n43997,n40306,n44023 );
   nor U44968 ( n44023,n28363,n41825 );
   not U44969 ( n41825,p2_ebx_reg_9_ );
   and U44970 ( n40306,n40399,n44024 );
   nand U44971 ( n44024,n42987,n41815 );
   not U44972 ( n41815,p2_ebx_reg_8_ );
   or U44973 ( n43996,n43017,n44025 );
   nor U44974 ( n44025,n28363,n41839 );
   not U44975 ( n41839,p2_ebx_reg_11_ );
   and U44976 ( n43017,n40399,n44026 );
   nand U44977 ( n44026,n42987,n41832 );
   not U44978 ( n41832,p2_ebx_reg_10_ );
   nor U44979 ( n43995,n43062,n44027 );
   nor U44980 ( n44027,n28362,n41857 );
   not U44981 ( n41857,p2_ebx_reg_13_ );
   and U44982 ( n43062,n40399,n44028 );
   nand U44983 ( n44028,n42987,n41846 );
   not U44984 ( n41846,p2_ebx_reg_12_ );
   or U44985 ( n43994,n43121,n44029 );
   nor U44986 ( n44029,n42988,n41874 );
   not U44987 ( n41874,p2_ebx_reg_15_ );
   and U44988 ( n43121,n40399,n44030 );
   nand U44989 ( n44030,n42987,n41865 );
   not U44990 ( n41865,p2_ebx_reg_14_ );
   nor U44991 ( n43993,n43179,n44031 );
   nor U44992 ( n44031,n28363,n41889 );
   not U44993 ( n41889,p2_ebx_reg_17_ );
   and U44994 ( n43179,n40399,n44032 );
   nand U44995 ( n44032,n42987,n41883 );
   not U44996 ( n41883,p2_ebx_reg_16_ );
   or U44997 ( n43992,n43239,n44033 );
   nor U44998 ( n44033,n28362,n41904 );
   not U44999 ( n41904,p2_ebx_reg_19_ );
   and U45000 ( n43239,n40399,n44034 );
   nand U45001 ( n44034,n28274,n41898 );
   not U45002 ( n41898,p2_ebx_reg_18_ );
   nor U45003 ( n43991,n43315,n44035 );
   nor U45004 ( n44035,n42988,n41919 );
   not U45005 ( n41919,p2_ebx_reg_21_ );
   and U45006 ( n43315,n40399,n44036 );
   nand U45007 ( n44036,n28274,n41913 );
   not U45008 ( n41913,p2_ebx_reg_20_ );
   nor U45009 ( n43990,n43371,n44037 );
   nor U45010 ( n44037,n28363,n41939 );
   not U45011 ( n41939,p2_ebx_reg_23_ );
   and U45012 ( n43371,n40399,n44038 );
   nand U45013 ( n44038,n28274,n41928 );
   not U45014 ( n41928,p2_ebx_reg_22_ );
   nor U45015 ( n43989,n43427,n44039 );
   nor U45016 ( n44039,n28362,n41963 );
   not U45017 ( n41963,p2_ebx_reg_25_ );
   and U45018 ( n43427,n40399,n44040 );
   nand U45019 ( n44040,n28274,n41952 );
   not U45020 ( n41952,p2_ebx_reg_24_ );
   nor U45021 ( n43988,n43466,n44041 );
   nor U45022 ( n44041,n42988,n41986 );
   not U45023 ( n41986,p2_ebx_reg_27_ );
   and U45024 ( n43466,n40399,n44042 );
   nand U45025 ( n44042,n28274,n41975 );
   not U45026 ( n41975,p2_ebx_reg_26_ );
   or U45027 ( n43987,n43523,n44043 );
   nor U45028 ( n44043,n28362,n42005 );
   not U45029 ( n42005,p2_ebx_reg_29_ );
   not U45030 ( n42988,n40399 );
   and U45031 ( n43523,n40399,n44044 );
   nand U45032 ( n44044,n28274,n41998 );
   not U45033 ( n41998,p2_ebx_reg_28_ );
   nand U45034 ( n40399,n38601,n28274 );
   nand U45035 ( n42987,n44022,n28239 );
   not U45036 ( n44022,n44045 );
   nand U45037 ( n42664,n44046,n44047 );
   nor U45038 ( n44047,n44048,n37132 );
   and U45039 ( n44046,p2_ebx_reg_31_,n42826 );
   nor U45040 ( n43610,n44049,n44050 );
   nand U45041 ( n44050,n44051,n44052 );
   nand U45042 ( n44052,n28355,n41758 );
   xor U45043 ( n41758,n44053,n43584 );
   nand U45044 ( n43584,n44054,n44055 );
   not U45045 ( n44055,n43525 );
   nand U45046 ( n43525,n44056,n43498 );
   not U45047 ( n43498,n43468 );
   nand U45048 ( n43468,n44057,n43444 );
   not U45049 ( n43444,n43410 );
   nand U45050 ( n43410,n44058,n43385 );
   not U45051 ( n43385,n43359 );
   nand U45052 ( n43359,n44059,n43332 );
   not U45053 ( n43332,n43304 );
   nand U45054 ( n43304,n44060,n43275 );
   not U45055 ( n43275,n43241 );
   nand U45056 ( n43241,n44061,n43218 );
   not U45057 ( n43218,n43181 );
   nand U45058 ( n43181,n44062,n43159 );
   not U45059 ( n43159,n43123 );
   nand U45060 ( n43123,n44063,n43100 );
   not U45061 ( n43100,n43064 );
   nand U45062 ( n43064,n44064,n43039 );
   not U45063 ( n43039,n43011 );
   nand U45064 ( n43011,n44065,n42980 );
   not U45065 ( n42980,n42954 );
   nand U45066 ( n42954,n42956,n42955 );
   nand U45067 ( n42955,n44066,n44067 );
   nor U45068 ( n44067,n44068,n44069 );
   nor U45069 ( n44069,n28369,n38925 );
   not U45070 ( n38925,p2_instaddrpointer_reg_8_ );
   and U45071 ( n44068,n42278,n44071 );
   nand U45072 ( n42278,n44072,n44073 );
   nor U45073 ( n44073,n44074,n44075 );
   nand U45074 ( n44075,n44076,n44077 );
   nor U45075 ( n44077,n44078,n44079 );
   nor U45076 ( n44079,n38693,n44080 );
   nor U45077 ( n44078,n40634,n44081 );
   nor U45078 ( n44076,n44082,n44083 );
   nor U45079 ( n44083,n40623,n44084 );
   nor U45080 ( n44082,n40616,n44085 );
   nand U45081 ( n44074,n44086,n44087 );
   nor U45082 ( n44087,n44088,n44089 );
   nor U45083 ( n44089,n40644,n44090 );
   nor U45084 ( n44088,n40613,n44091 );
   nor U45085 ( n44086,n44092,n44093 );
   nor U45086 ( n44093,n40612,n44094 );
   nor U45087 ( n44092,n40643,n44095 );
   nor U45088 ( n44072,n44096,n44097 );
   nand U45089 ( n44097,n44098,n44099 );
   nor U45090 ( n44099,n44100,n44101 );
   nor U45091 ( n44101,n40626,n44102 );
   nor U45092 ( n44100,n40647,n44103 );
   nor U45093 ( n44098,n44104,n44105 );
   nor U45094 ( n44105,n40622,n44106 );
   nor U45095 ( n44104,n40617,n44107 );
   nand U45096 ( n44096,n44108,n44109 );
   nor U45097 ( n44109,n44110,n44111 );
   nor U45098 ( n44111,n40638,n44112 );
   nor U45099 ( n44110,n40635,n44113 );
   nor U45100 ( n44108,n44114,n44115 );
   nor U45101 ( n44115,n40648,n44116 );
   nor U45102 ( n44114,n40627,n44117 );
   nor U45103 ( n44066,n44118,n44119 );
   nor U45104 ( n44119,n44120,n40924 );
   not U45105 ( n40924,p2_eax_reg_8_ );
   nor U45106 ( n44118,n44121,n36925 );
   not U45107 ( n36925,p2_reip_reg_8_ );
   and U45108 ( n42956,n44122,n44123 );
   nand U45109 ( n44123,n44124,n42923 );
   nand U45110 ( n42923,n44125,n44126 );
   nand U45111 ( n44126,n42895,n44127 );
   or U45112 ( n44127,n42893,n42894 );
   and U45113 ( n42895,n44128,n44129 );
   nand U45114 ( n44129,p2_instaddrpointer_reg_6_,n44130 );
   nor U45115 ( n44128,n44131,n44132 );
   nor U45116 ( n44132,n28149,n36935 );
   not U45117 ( n36935,p2_reip_reg_6_ );
   nor U45118 ( n44131,n44120,n40934 );
   not U45119 ( n40934,p2_eax_reg_6_ );
   nand U45120 ( n44125,n42893,n42894 );
   nand U45121 ( n42894,n44071,n40500 );
   nand U45122 ( n42893,n44133,n44134 );
   nand U45123 ( n44134,n44135,n42803 );
   nand U45124 ( n42803,n44136,n44137 );
   nand U45125 ( n44137,n42766,n44138 );
   or U45126 ( n44138,n42764,n42765 );
   and U45127 ( n42766,n44139,n44140 );
   nand U45128 ( n44140,p2_instaddrpointer_reg_4_,n44130 );
   nor U45129 ( n44139,n44141,n44142 );
   nor U45130 ( n44142,n28150,n36945 );
   not U45131 ( n36945,p2_reip_reg_4_ );
   nor U45132 ( n44141,n44120,n40944 );
   not U45133 ( n40944,p2_eax_reg_4_ );
   nand U45134 ( n44136,n42764,n42765 );
   nand U45135 ( n42765,n44071,n40798 );
   nand U45136 ( n42764,n44143,n44144 );
   nand U45137 ( n44144,n42747,n44145 );
   nand U45138 ( n44145,n42745,n42748 );
   and U45139 ( n42747,n44146,n44147 );
   nand U45140 ( n44147,n44071,n40550 );
   nand U45141 ( n44146,p2_state2_reg_3_,p2_instqueuewr_addr_reg_3_ );
   or U45142 ( n44143,n42748,n42745 );
   and U45143 ( n42745,n44148,n44149 );
   nand U45144 ( n44149,n42705,n44150 );
   nand U45145 ( n44150,n42704,n42706 );
   and U45146 ( n42705,n44151,n44152 );
   nand U45147 ( n44152,n42630,n44153 );
   or U45148 ( n44153,n42674,n42675 );
   nor U45149 ( n42630,n42633,n42632 );
   and U45150 ( n42632,n44154,n44155 );
   nor U45151 ( n44155,n44156,n44157 );
   nor U45152 ( n44154,n44158,n44159 );
   and U45153 ( n44159,n40602,n44071 );
   nor U45154 ( n44158,n37336,n38681 );
   not U45155 ( n37336,p2_instqueuewr_addr_reg_0_ );
   and U45156 ( n42633,n44160,n44161 );
   nor U45157 ( n44161,p2_state2_reg_3_,n44162 );
   nor U45158 ( n44162,n28368,n36762 );
   not U45159 ( n36762,p2_instaddrpointer_reg_0_ );
   nor U45160 ( n44160,n44163,n44164 );
   nor U45161 ( n44164,n28330,n40964 );
   not U45162 ( n40964,p2_eax_reg_0_ );
   nor U45163 ( n44163,n39602,n28149 );
   nand U45164 ( n44151,n42674,n42675 );
   nand U45165 ( n42675,n44165,n44166 );
   nor U45166 ( n44166,n44167,n44168 );
   nor U45167 ( n44168,n41567,n44169 );
   nor U45168 ( n44165,n44170,n44171 );
   nor U45169 ( n44171,n37096,n38681 );
   and U45170 ( n44170,n40651,n44071 );
   nand U45171 ( n42674,n44172,n44173 );
   nand U45172 ( n44173,p2_eax_reg_1_,n44156 );
   nor U45173 ( n44172,n44174,n44175 );
   nor U45174 ( n44175,n44121,n36961 );
   nor U45175 ( n44174,n44070,n36758 );
   not U45176 ( n36758,p2_instaddrpointer_reg_1_ );
   or U45177 ( n44148,n42704,n42706 );
   nand U45178 ( n42706,n44176,n44177 );
   nand U45179 ( n44177,p2_instaddrpointer_reg_2_,n44130 );
   nor U45180 ( n44176,n44178,n44179 );
   nor U45181 ( n44179,n28149,n36955 );
   not U45182 ( n36955,p2_reip_reg_2_ );
   nor U45183 ( n44178,n44120,n40954 );
   not U45184 ( n40954,p2_eax_reg_2_ );
   nand U45185 ( n42704,n44180,n44181 );
   nand U45186 ( n44181,p2_state2_reg_3_,p2_instqueuewr_addr_reg_2_ );
   nor U45187 ( n44180,n44157,n44182 );
   and U45188 ( n44182,n40700,n44071 );
   nand U45189 ( n42748,n44183,n44184 );
   nand U45190 ( n44184,p2_instaddrpointer_reg_3_,n44130 );
   nor U45191 ( n44183,n44185,n44186 );
   nor U45192 ( n44186,n44121,n36950 );
   not U45193 ( n36950,p2_reip_reg_3_ );
   nor U45194 ( n44185,n44120,n40949 );
   not U45195 ( n40949,p2_eax_reg_3_ );
   nand U45196 ( n44135,n42801,n42802 );
   or U45197 ( n44133,n42802,n42801 );
   and U45198 ( n42801,n44071,n40749 );
   nand U45199 ( n40749,n44187,n44188 );
   nor U45200 ( n44188,n44189,n44190 );
   nand U45201 ( n44190,n44191,n44192 );
   nor U45202 ( n44192,n44193,n44194 );
   nor U45203 ( n44194,n40773,n44195 );
   nor U45204 ( n44193,n40770,n44196 );
   nor U45205 ( n44191,n44197,n44198 );
   nor U45206 ( n44198,n40764,n44199 );
   nor U45207 ( n44197,n40785,n44200 );
   nand U45208 ( n44189,n44201,n44202 );
   nor U45209 ( n44202,n44203,n44204 );
   nor U45210 ( n44204,n40784,n44205 );
   nor U45211 ( n44203,n40763,n44206 );
   nor U45212 ( n44201,n44207,n44208 );
   nor U45213 ( n44208,n40790,n44209 );
   nor U45214 ( n44207,n40791,n44210 );
   nor U45215 ( n44187,n44211,n44212 );
   nand U45216 ( n44212,n44213,n44214 );
   nor U45217 ( n44214,n44215,n44216 );
   nor U45218 ( n44216,n40794,n44217 );
   nor U45219 ( n44215,n40795,n44218 );
   nor U45220 ( n44213,n44219,n44220 );
   nor U45221 ( n44220,n40780,n44221 );
   nor U45222 ( n44219,n40781,n44222 );
   nand U45223 ( n44211,n44223,n44224 );
   nor U45224 ( n44224,n44225,n44226 );
   nor U45225 ( n44226,n38606,n44227 );
   nor U45226 ( n44225,n40759,n44228 );
   nor U45227 ( n44223,n44229,n44230 );
   nor U45228 ( n44230,n40769,n44231 );
   nor U45229 ( n44229,n40760,n44232 );
   nand U45230 ( n42802,n44233,n44234 );
   nand U45231 ( n44234,p2_instaddrpointer_reg_5_,n44130 );
   nor U45232 ( n44233,n44235,n44236 );
   nor U45233 ( n44236,n28150,n36940 );
   not U45234 ( n36940,p2_reip_reg_5_ );
   nor U45235 ( n44235,n44120,n40939 );
   not U45236 ( n40939,p2_eax_reg_5_ );
   nand U45237 ( n44124,n42921,n42922 );
   or U45238 ( n44122,n42922,n42921 );
   nor U45239 ( n42921,n44237,n28370 );
   not U45240 ( n40219,n40229 );
   nand U45241 ( n40229,n44238,n44239 );
   nor U45242 ( n44239,n44240,n44241 );
   nand U45243 ( n44241,n44242,n44243 );
   nor U45244 ( n44243,n44244,n44245 );
   nor U45245 ( n44245,n40487,n44195 );
   nor U45246 ( n44244,n40484,n44196 );
   nor U45247 ( n44242,n44246,n44247 );
   nor U45248 ( n44247,n40497,n44199 );
   nor U45249 ( n44246,n40476,n44200 );
   nand U45250 ( n44240,n44248,n44249 );
   nor U45251 ( n44249,n44250,n44251 );
   nor U45252 ( n44251,n40475,n44205 );
   nor U45253 ( n44250,n40496,n44206 );
   nor U45254 ( n44248,n44252,n44253 );
   nor U45255 ( n44253,n40461,n44209 );
   nor U45256 ( n44252,n40462,n44210 );
   nor U45257 ( n44238,n44254,n44255 );
   nand U45258 ( n44255,n44256,n44257 );
   nor U45259 ( n44257,n44258,n44259 );
   nor U45260 ( n44259,n40465,n44217 );
   nor U45261 ( n44258,n40466,n44218 );
   nor U45262 ( n44256,n44260,n44261 );
   nor U45263 ( n44261,n40471,n44221 );
   nor U45264 ( n44260,n40472,n44222 );
   nand U45265 ( n44254,n44262,n44263 );
   nor U45266 ( n44263,n44264,n44265 );
   nor U45267 ( n44265,n38572,n44227 );
   nor U45268 ( n44264,n40492,n44228 );
   nor U45269 ( n44262,n44266,n44267 );
   nor U45270 ( n44267,n40483,n44231 );
   nor U45271 ( n44266,n40493,n44232 );
   nand U45272 ( n42922,n44268,n44269 );
   nand U45273 ( n44269,p2_instaddrpointer_reg_7_,n44130 );
   nor U45274 ( n44268,n44270,n44271 );
   nor U45275 ( n44271,n28150,n36930 );
   not U45276 ( n36930,p2_reip_reg_7_ );
   nor U45277 ( n44270,n44120,n40929 );
   not U45278 ( n40929,p2_eax_reg_7_ );
   nor U45279 ( n44065,n42979,n43012 );
   and U45280 ( n43012,n44272,n44273 );
   nor U45281 ( n44273,n44274,n44275 );
   nor U45282 ( n44275,n28369,n38974 );
   not U45283 ( n38974,p2_instaddrpointer_reg_10_ );
   and U45284 ( n44274,n41829,n44071 );
   nand U45285 ( n41829,n44276,n44277 );
   nor U45286 ( n44277,n44278,n44279 );
   nand U45287 ( n44279,n44280,n44281 );
   nor U45288 ( n44281,n44282,n44283 );
   nor U45289 ( n44283,n40736,n44112 );
   nor U45290 ( n44282,n40733,n44113 );
   nor U45291 ( n44280,n44284,n44285 );
   nor U45292 ( n44285,n40746,n44116 );
   nor U45293 ( n44284,n40725,n44117 );
   nand U45294 ( n44278,n44286,n44287 );
   nor U45295 ( n44287,n44288,n44289 );
   nor U45296 ( n44289,n40724,n44102 );
   nor U45297 ( n44288,n40745,n44103 );
   nor U45298 ( n44286,n44290,n44291 );
   nor U45299 ( n44291,n40720,n44106 );
   nor U45300 ( n44290,n40715,n44107 );
   nor U45301 ( n44276,n44292,n44293 );
   nand U45302 ( n44293,n44294,n44295 );
   nor U45303 ( n44295,n44296,n44297 );
   nor U45304 ( n44297,n40742,n44090 );
   nor U45305 ( n44296,n40711,n44091 );
   nor U45306 ( n44294,n44298,n44299 );
   nor U45307 ( n44299,n40710,n44094 );
   nor U45308 ( n44298,n40741,n44095 );
   nand U45309 ( n44292,n44300,n44301 );
   nor U45310 ( n44301,n44302,n44303 );
   nor U45311 ( n44303,n38654,n44080 );
   nor U45312 ( n44302,n40732,n44081 );
   nor U45313 ( n44300,n44304,n44305 );
   nor U45314 ( n44305,n40721,n44084 );
   nor U45315 ( n44304,n40714,n44085 );
   nor U45316 ( n44272,n44306,n44307 );
   nor U45317 ( n44307,n44120,n40914 );
   not U45318 ( n40914,p2_eax_reg_10_ );
   nor U45319 ( n44306,n44121,n36915 );
   not U45320 ( n36915,p2_reip_reg_10_ );
   not U45321 ( n42979,n43014 );
   nand U45322 ( n43014,n44308,n44309 );
   nor U45323 ( n44309,n44310,n44311 );
   nor U45324 ( n44311,n28369,n38948 );
   not U45325 ( n38948,p2_instaddrpointer_reg_9_ );
   and U45326 ( n44310,n42279,n44071 );
   nand U45327 ( n42279,n44312,n44313 );
   nor U45328 ( n44313,n44314,n44315 );
   nand U45329 ( n44315,n44316,n44317 );
   nor U45330 ( n44317,n44318,n44319 );
   nor U45331 ( n44319,n40687,n44112 );
   nor U45332 ( n44318,n40684,n44113 );
   nor U45333 ( n44316,n44320,n44321 );
   nor U45334 ( n44321,n40697,n44116 );
   nor U45335 ( n44320,n40676,n44117 );
   nand U45336 ( n44314,n44322,n44323 );
   nor U45337 ( n44323,n44324,n44325 );
   nor U45338 ( n44325,n40675,n44102 );
   nor U45339 ( n44324,n40696,n44103 );
   nor U45340 ( n44322,n44326,n44327 );
   nor U45341 ( n44327,n40671,n44106 );
   nor U45342 ( n44326,n40666,n44107 );
   nor U45343 ( n44312,n44328,n44329 );
   nand U45344 ( n44329,n44330,n44331 );
   nor U45345 ( n44331,n44332,n44333 );
   nor U45346 ( n44333,n40693,n44090 );
   nor U45347 ( n44332,n40662,n44091 );
   nor U45348 ( n44330,n44334,n44335 );
   nor U45349 ( n44335,n40661,n44094 );
   nor U45350 ( n44334,n40692,n44095 );
   nand U45351 ( n44328,n44336,n44337 );
   nor U45352 ( n44337,n44338,n44339 );
   nor U45353 ( n44339,n38669,n44080 );
   nor U45354 ( n44338,n40683,n44081 );
   nor U45355 ( n44336,n44340,n44341 );
   nor U45356 ( n44341,n40672,n44084 );
   nor U45357 ( n44340,n40665,n44085 );
   nor U45358 ( n44308,n44342,n44343 );
   nor U45359 ( n44343,n44120,n40919 );
   not U45360 ( n40919,p2_eax_reg_9_ );
   nor U45361 ( n44342,n28149,n36920 );
   not U45362 ( n36920,p2_reip_reg_9_ );
   nor U45363 ( n44064,n43038,n43065 );
   and U45364 ( n43065,n44344,n44345 );
   nor U45365 ( n44345,n44346,n44347 );
   nor U45366 ( n44347,n44070,n39022 );
   not U45367 ( n39022,p2_instaddrpointer_reg_12_ );
   and U45368 ( n44346,n42280,n44071 );
   nand U45369 ( n42280,n44348,n44349 );
   nor U45370 ( n44349,n44350,n44351 );
   nand U45371 ( n44351,n44352,n44353 );
   nor U45372 ( n44353,n44354,n44355 );
   nor U45373 ( n44355,n38622,n44080 );
   nor U45374 ( n44354,n40838,n44081 );
   nor U45375 ( n44352,n44356,n44357 );
   nor U45376 ( n44357,n40825,n44084 );
   nor U45377 ( n44356,n40816,n44085 );
   nand U45378 ( n44350,n44358,n44359 );
   nor U45379 ( n44359,n44360,n44361 );
   nor U45380 ( n44361,n40849,n44090 );
   nor U45381 ( n44360,n40811,n44091 );
   nor U45382 ( n44358,n44362,n44363 );
   nor U45383 ( n44363,n40808,n44094 );
   nor U45384 ( n44362,n40848,n44095 );
   nor U45385 ( n44348,n44364,n44365 );
   nand U45386 ( n44365,n44366,n44367 );
   nor U45387 ( n44367,n44368,n44369 );
   nor U45388 ( n44369,n40828,n44102 );
   nor U45389 ( n44368,n40852,n44103 );
   nor U45390 ( n44366,n44370,n44371 );
   nor U45391 ( n44371,n40823,n44106 );
   nor U45392 ( n44370,n40817,n44107 );
   nand U45393 ( n44364,n44372,n44373 );
   nor U45394 ( n44373,n44374,n44375 );
   nor U45395 ( n44375,n40842,n44112 );
   nor U45396 ( n44374,n40839,n44113 );
   nor U45397 ( n44372,n44376,n44377 );
   nor U45398 ( n44377,n40853,n44116 );
   nor U45399 ( n44376,n40830,n44117 );
   nor U45400 ( n44344,n44378,n44379 );
   nor U45401 ( n44379,n28330,n40904 );
   not U45402 ( n40904,p2_eax_reg_12_ );
   nor U45403 ( n44378,n28150,n36905 );
   not U45404 ( n36905,p2_reip_reg_12_ );
   not U45405 ( n43038,n43067 );
   nand U45406 ( n43067,n44380,n44381 );
   nor U45407 ( n44381,n44382,n44383 );
   nor U45408 ( n44383,n44070,n38996 );
   not U45409 ( n38996,p2_instaddrpointer_reg_11_ );
   and U45410 ( n44382,n42275,n44071 );
   nand U45411 ( n42275,n44384,n44385 );
   nor U45412 ( n44385,n44386,n44387 );
   nand U45413 ( n44387,n44388,n44389 );
   nor U45414 ( n44389,n44390,n44391 );
   nor U45415 ( n44391,n40574,n44112 );
   nor U45416 ( n44390,n40571,n44113 );
   nor U45417 ( n44388,n44392,n44393 );
   nor U45418 ( n44393,n40565,n44116 );
   nor U45419 ( n44392,n40586,n44117 );
   nand U45420 ( n44386,n44394,n44395 );
   nor U45421 ( n44395,n44396,n44397 );
   nor U45422 ( n44397,n40585,n44102 );
   nor U45423 ( n44396,n40564,n44103 );
   nor U45424 ( n44394,n44398,n44399 );
   nor U45425 ( n44399,n40581,n44106 );
   nor U45426 ( n44398,n40596,n44107 );
   nor U45427 ( n44384,n44400,n44401 );
   nand U45428 ( n44401,n44402,n44403 );
   nor U45429 ( n44403,n44404,n44405 );
   nor U45430 ( n44405,n40561,n44090 );
   nor U45431 ( n44404,n40592,n44091 );
   nor U45432 ( n44402,n44406,n44407 );
   nor U45433 ( n44407,n40591,n44094 );
   nor U45434 ( n44406,n40560,n44095 );
   nand U45435 ( n44400,n44408,n44409 );
   nor U45436 ( n44409,n44410,n44411 );
   nor U45437 ( n44411,n38638,n44080 );
   nor U45438 ( n44410,n40570,n44081 );
   nor U45439 ( n44408,n44412,n44413 );
   nor U45440 ( n44413,n40582,n44084 );
   nor U45441 ( n44412,n40595,n44085 );
   nor U45442 ( n44380,n44414,n44415 );
   nor U45443 ( n44415,n28330,n40909 );
   not U45444 ( n40909,p2_eax_reg_11_ );
   nor U45445 ( n44414,n28150,n36910 );
   not U45446 ( n36910,p2_reip_reg_11_ );
   nor U45447 ( n44063,n43099,n43124 );
   and U45448 ( n43124,n44416,n44417 );
   nor U45449 ( n44417,n44418,n44419 );
   nor U45450 ( n44419,n28369,n39070 );
   not U45451 ( n39070,p2_instaddrpointer_reg_14_ );
   nor U45452 ( n44418,n41861,n44237 );
   and U45453 ( n41861,n44420,n44421 );
   nor U45454 ( n44421,n44422,n44423 );
   nand U45455 ( n44423,n44424,n44425 );
   nor U45456 ( n44425,n44426,n44427 );
   nor U45457 ( n44427,n40536,n44112 );
   nor U45458 ( n44426,n40533,n44113 );
   nor U45459 ( n44424,n44428,n44429 );
   nor U45460 ( n44429,n40546,n44116 );
   nor U45461 ( n44428,n40525,n44117 );
   nand U45462 ( n44422,n44430,n44431 );
   nor U45463 ( n44431,n44432,n44433 );
   nor U45464 ( n44433,n40524,n44102 );
   nor U45465 ( n44432,n40545,n44103 );
   nor U45466 ( n44430,n44434,n44435 );
   nor U45467 ( n44435,n40520,n44106 );
   nor U45468 ( n44434,n40515,n44107 );
   nor U45469 ( n44420,n44436,n44437 );
   nand U45470 ( n44437,n44438,n44439 );
   nor U45471 ( n44439,n44440,n44441 );
   nor U45472 ( n44441,n40542,n44090 );
   nor U45473 ( n44440,n40511,n44091 );
   nor U45474 ( n44438,n44442,n44443 );
   nor U45475 ( n44443,n40510,n44094 );
   nor U45476 ( n44442,n40541,n44095 );
   nand U45477 ( n44436,n44444,n44445 );
   nor U45478 ( n44445,n44446,n44447 );
   nor U45479 ( n44447,n38590,n44080 );
   nor U45480 ( n44446,n40532,n44081 );
   nor U45481 ( n44444,n44448,n44449 );
   nor U45482 ( n44449,n40521,n44084 );
   nor U45483 ( n44448,n40514,n44085 );
   nor U45484 ( n44416,n44450,n44451 );
   nor U45485 ( n44451,n28330,n40894 );
   not U45486 ( n40894,p2_eax_reg_14_ );
   nor U45487 ( n44450,n28149,n36895 );
   not U45488 ( n36895,p2_reip_reg_14_ );
   not U45489 ( n43099,n43126 );
   nand U45490 ( n43126,n44452,n44453 );
   nor U45491 ( n44453,n44454,n44455 );
   nor U45492 ( n44455,n28368,n39043 );
   not U45493 ( n39043,p2_instaddrpointer_reg_13_ );
   and U45494 ( n44454,n42281,n44071 );
   nand U45495 ( n42281,n44456,n44457 );
   nor U45496 ( n44457,n44458,n44459 );
   nand U45497 ( n44459,n44460,n44461 );
   nor U45498 ( n44461,n44462,n44463 );
   nor U45499 ( n44463,n40773,n44112 );
   nor U45500 ( n44462,n40770,n44113 );
   nor U45501 ( n44460,n44464,n44465 );
   nor U45502 ( n44465,n40764,n44116 );
   nor U45503 ( n44464,n40785,n44117 );
   nand U45504 ( n44458,n44466,n44467 );
   nor U45505 ( n44467,n44468,n44469 );
   nor U45506 ( n44469,n40784,n44102 );
   nor U45507 ( n44468,n40763,n44103 );
   nor U45508 ( n44466,n44470,n44471 );
   nor U45509 ( n44471,n40780,n44106 );
   nor U45510 ( n44470,n40795,n44107 );
   nor U45511 ( n44456,n44472,n44473 );
   nand U45512 ( n44473,n44474,n44475 );
   nor U45513 ( n44475,n44476,n44477 );
   nor U45514 ( n44477,n40760,n44090 );
   nor U45515 ( n44476,n40791,n44091 );
   nor U45516 ( n44474,n44478,n44479 );
   nor U45517 ( n44479,n40790,n44094 );
   nor U45518 ( n44478,n40759,n44095 );
   nand U45519 ( n44472,n44480,n44481 );
   nor U45520 ( n44481,n44482,n44483 );
   nor U45521 ( n44483,n38606,n44080 );
   nor U45522 ( n44482,n40769,n44081 );
   nor U45523 ( n44480,n44484,n44485 );
   nor U45524 ( n44485,n40781,n44084 );
   nor U45525 ( n44484,n40794,n44085 );
   nor U45526 ( n44452,n44486,n44487 );
   nor U45527 ( n44487,n28330,n40899 );
   not U45528 ( n40899,p2_eax_reg_13_ );
   nor U45529 ( n44486,n28150,n36900 );
   not U45530 ( n36900,p2_reip_reg_13_ );
   nor U45531 ( n44062,n43158,n43182 );
   and U45532 ( n43182,n44488,n44489 );
   nand U45533 ( n44489,p2_eax_reg_16_,n44156 );
   nor U45534 ( n44488,n44490,n44491 );
   nor U45535 ( n44491,n44121,n36885 );
   not U45536 ( n36885,p2_reip_reg_16_ );
   nor U45537 ( n44490,n44070,n39118 );
   not U45538 ( n39118,p2_instaddrpointer_reg_16_ );
   not U45539 ( n43158,n43184 );
   nand U45540 ( n43184,n44492,n44493 );
   nor U45541 ( n44493,n44494,n44495 );
   nor U45542 ( n44495,n28368,n39092 );
   not U45543 ( n39092,p2_instaddrpointer_reg_15_ );
   and U45544 ( n44494,n41870,n44071 );
   not U45545 ( n44071,n44237 );
   nand U45546 ( n44237,n44496,n27896 );
   nor U45547 ( n44496,p2_state2_reg_3_,n42814 );
   nand U45548 ( n41870,n44497,n44498 );
   nor U45549 ( n44498,n44499,n44500 );
   nand U45550 ( n44500,n44501,n44502 );
   nor U45551 ( n44502,n44503,n44504 );
   nor U45552 ( n44504,n40487,n44112 );
   nand U45553 ( n44112,n44505,n44506 );
   nor U45554 ( n44503,n40484,n44113 );
   nand U45555 ( n44113,n44505,n42450 );
   nor U45556 ( n44501,n44507,n44508 );
   nor U45557 ( n44508,n40497,n44116 );
   nand U45558 ( n44116,n44505,n42582 );
   nor U45559 ( n44507,n40476,n44117 );
   nand U45560 ( n44117,n44509,n44506 );
   nand U45561 ( n44499,n44510,n44511 );
   nor U45562 ( n44511,n44512,n44513 );
   nor U45563 ( n44513,n40475,n44102 );
   nand U45564 ( n44102,n44509,n42450 );
   nor U45565 ( n44512,n40496,n44103 );
   nand U45566 ( n44103,n44509,n42582 );
   nor U45567 ( n44510,n44514,n44515 );
   nor U45568 ( n44515,n40471,n44106 );
   nand U45569 ( n44106,n44516,n44506 );
   nor U45570 ( n44514,n40466,n44107 );
   nand U45571 ( n44107,n44516,n42450 );
   nor U45572 ( n44497,n44517,n44518 );
   nand U45573 ( n44518,n44519,n44520 );
   nor U45574 ( n44520,n44521,n44522 );
   nor U45575 ( n44522,n40493,n44090 );
   nand U45576 ( n44090,n44516,n42582 );
   nor U45577 ( n44521,n40462,n44091 );
   nand U45578 ( n44091,n44523,n44506 );
   nor U45579 ( n44519,n44524,n44525 );
   nor U45580 ( n44525,n40461,n44094 );
   nand U45581 ( n44094,n44523,n42450 );
   nor U45582 ( n44524,n40492,n44095 );
   nand U45583 ( n44095,n44523,n42582 );
   nand U45584 ( n44517,n44526,n44527 );
   nor U45585 ( n44527,n44528,n44529 );
   nor U45586 ( n44529,n38572,n44080 );
   nand U45587 ( n44080,n44505,n44530 );
   nor U45588 ( n44505,n44531,n44532 );
   nor U45589 ( n44528,n40483,n44081 );
   nand U45590 ( n44081,n44509,n44530 );
   nor U45591 ( n44509,n44531,n37186 );
   nor U45592 ( n44526,n44533,n44534 );
   nor U45593 ( n44534,n40472,n44084 );
   nand U45594 ( n44084,n44516,n44530 );
   nor U45595 ( n44516,n37158,n44532 );
   not U45596 ( n44532,n37186 );
   nor U45597 ( n44533,n40465,n44085 );
   nand U45598 ( n44085,n44523,n44530 );
   nor U45599 ( n44523,n37186,n37158 );
   not U45600 ( n37158,n44531 );
   xor U45601 ( n44531,n37139,n36779 );
   nand U45602 ( n37186,n36779,n44535 );
   nand U45603 ( n44535,n37120,n37154 );
   nor U45604 ( n44492,n44536,n44537 );
   nor U45605 ( n44537,n28330,n40887 );
   not U45606 ( n40887,p2_eax_reg_15_ );
   nor U45607 ( n44536,n28149,n36890 );
   not U45608 ( n36890,p2_reip_reg_15_ );
   nor U45609 ( n44061,n43217,n43242 );
   and U45610 ( n43242,n44538,n44539 );
   nand U45611 ( n44539,p2_eax_reg_18_,n44156 );
   nor U45612 ( n44538,n44540,n44541 );
   nor U45613 ( n44541,n44121,n36875 );
   not U45614 ( n36875,p2_reip_reg_18_ );
   nor U45615 ( n44540,n28368,n39166 );
   not U45616 ( n39166,p2_instaddrpointer_reg_18_ );
   not U45617 ( n43217,n43244 );
   nand U45618 ( n43244,n44542,n44543 );
   nand U45619 ( n44543,p2_eax_reg_17_,n44156 );
   nor U45620 ( n44542,n44544,n44545 );
   nor U45621 ( n44545,n28150,n36880 );
   not U45622 ( n36880,p2_reip_reg_17_ );
   nor U45623 ( n44544,n28369,n39140 );
   not U45624 ( n39140,p2_instaddrpointer_reg_17_ );
   nor U45625 ( n44060,n43274,n43305 );
   and U45626 ( n43305,n44546,n44547 );
   nand U45627 ( n44547,p2_eax_reg_20_,n44156 );
   nor U45628 ( n44546,n44548,n44549 );
   nor U45629 ( n44549,n28149,n36865 );
   not U45630 ( n36865,p2_reip_reg_20_ );
   nor U45631 ( n44548,n44070,n39212 );
   not U45632 ( n39212,p2_instaddrpointer_reg_20_ );
   not U45633 ( n43274,n43307 );
   nand U45634 ( n43307,n44550,n44551 );
   nand U45635 ( n44551,p2_eax_reg_19_,n44156 );
   nor U45636 ( n44550,n44552,n44553 );
   nor U45637 ( n44553,n44121,n36870 );
   not U45638 ( n36870,p2_reip_reg_19_ );
   nor U45639 ( n44552,n28368,n39188 );
   not U45640 ( n39188,p2_instaddrpointer_reg_19_ );
   nor U45641 ( n44059,n43331,n43360 );
   and U45642 ( n43360,n44554,n44555 );
   nand U45643 ( n44555,p2_eax_reg_22_,n44156 );
   nor U45644 ( n44554,n44556,n44557 );
   nor U45645 ( n44557,n44121,n36855 );
   not U45646 ( n36855,p2_reip_reg_22_ );
   nor U45647 ( n44556,n28369,n39261 );
   not U45648 ( n39261,p2_instaddrpointer_reg_22_ );
   not U45649 ( n43331,n43362 );
   nand U45650 ( n43362,n44558,n44559 );
   nand U45651 ( n44559,p2_eax_reg_21_,n44156 );
   nor U45652 ( n44558,n44560,n44561 );
   nor U45653 ( n44561,n28149,n36860 );
   not U45654 ( n36860,p2_reip_reg_21_ );
   nor U45655 ( n44560,n44070,n39234 );
   not U45656 ( n39234,p2_instaddrpointer_reg_21_ );
   nor U45657 ( n44058,n43384,n43411 );
   and U45658 ( n43411,n44562,n44563 );
   nand U45659 ( n44563,p2_eax_reg_24_,n44156 );
   nor U45660 ( n44562,n44564,n44565 );
   nor U45661 ( n44565,n28150,n36845 );
   not U45662 ( n36845,p2_reip_reg_24_ );
   nor U45663 ( n44564,n28368,n39309 );
   not U45664 ( n39309,p2_instaddrpointer_reg_24_ );
   not U45665 ( n43384,n43413 );
   nand U45666 ( n43413,n44566,n44567 );
   nand U45667 ( n44567,p2_eax_reg_23_,n44156 );
   nor U45668 ( n44566,n44568,n44569 );
   nor U45669 ( n44569,n44121,n36850 );
   not U45670 ( n36850,p2_reip_reg_23_ );
   nor U45671 ( n44568,n28369,n39283 );
   not U45672 ( n39283,p2_instaddrpointer_reg_23_ );
   nor U45673 ( n44057,n43443,n43469 );
   and U45674 ( n43469,n44570,n44571 );
   nand U45675 ( n44571,p2_eax_reg_26_,n44156 );
   nor U45676 ( n44570,n44572,n44573 );
   nor U45677 ( n44573,n28149,n36835 );
   not U45678 ( n36835,p2_reip_reg_26_ );
   nor U45679 ( n44572,n44070,n39357 );
   not U45680 ( n39357,p2_instaddrpointer_reg_26_ );
   not U45681 ( n43443,n43471 );
   nand U45682 ( n43471,n44574,n44575 );
   nand U45683 ( n44575,p2_eax_reg_25_,n44156 );
   nor U45684 ( n44574,n44576,n44577 );
   nor U45685 ( n44577,n28150,n36840 );
   not U45686 ( n36840,p2_reip_reg_25_ );
   nor U45687 ( n44576,n28368,n39331 );
   not U45688 ( n39331,p2_instaddrpointer_reg_25_ );
   nor U45689 ( n44056,n43497,n43526 );
   and U45690 ( n43526,n44578,n44579 );
   nand U45691 ( n44579,p2_eax_reg_28_,n44156 );
   nor U45692 ( n44578,n44580,n44581 );
   nor U45693 ( n44581,n44121,n36825 );
   not U45694 ( n36825,p2_reip_reg_28_ );
   nor U45695 ( n44580,n28369,n39396 );
   not U45696 ( n39396,p2_instaddrpointer_reg_28_ );
   not U45697 ( n43497,n43528 );
   nand U45698 ( n43528,n44582,n44583 );
   nand U45699 ( n44583,p2_eax_reg_27_,n44156 );
   nor U45700 ( n44582,n44584,n44585 );
   nor U45701 ( n44585,n28149,n36830 );
   not U45702 ( n36830,p2_reip_reg_27_ );
   nor U45703 ( n44584,n44070,n39379 );
   not U45704 ( n39379,p2_instaddrpointer_reg_27_ );
   nor U45705 ( n44054,n43558,n44586 );
   nor U45706 ( n44586,n43589,n44587 );
   or U45707 ( n44587,n43588,n43587 );
   nor U45708 ( n43587,n40968,n28330 );
   not U45709 ( n40968,p2_eax_reg_30_ );
   nor U45710 ( n43588,n39435,n28368 );
   not U45711 ( n39435,p2_instaddrpointer_reg_30_ );
   nor U45712 ( n43589,n36815,n28150 );
   not U45713 ( n36815,p2_reip_reg_30_ );
   and U45714 ( n43558,n44588,n44589 );
   nand U45715 ( n44589,p2_eax_reg_29_,n44156 );
   nor U45716 ( n44588,n44590,n44591 );
   nor U45717 ( n44591,n28149,n36820 );
   not U45718 ( n36820,p2_reip_reg_29_ );
   nor U45719 ( n44590,n28368,n39416 );
   not U45720 ( n39416,p2_instaddrpointer_reg_29_ );
   not U45721 ( n44070,n44130 );
   nor U45722 ( n44053,n44592,n44593 );
   nand U45723 ( n44593,n44594,n44595 );
   nand U45724 ( n44595,p2_instaddrpointer_reg_31_,n44130 );
   nand U45725 ( n44130,n44596,n44597 );
   nand U45726 ( n44597,n44598,n38585 );
   nor U45727 ( n44596,n44157,n44167 );
   and U45728 ( n44167,n44599,n42814 );
   and U45729 ( n44157,n44599,n41567 );
   nor U45730 ( n41567,n38585,n42814 );
   nor U45731 ( n44599,p2_state2_reg_3_,n39545 );
   or U45732 ( n44594,n36813,n44121 );
   nand U45733 ( n44121,n44600,n44598 );
   not U45734 ( n44598,n44169 );
   nand U45735 ( n44169,n44601,n44602 );
   nor U45736 ( n44601,p2_state2_reg_3_,n39566 );
   nor U45737 ( n44600,n38601,n36646 );
   nor U45738 ( n44592,n44120,n41746 );
   not U45739 ( n41746,p2_eax_reg_31_ );
   not U45740 ( n44120,n44156 );
   nor U45741 ( n44156,n38565,p2_state2_reg_3_ );
   not U45742 ( n42629,n42744 );
   nand U45743 ( n42744,n44603,n42826 );
   nor U45744 ( n44603,n37203,n44604 );
   not U45745 ( n37203,n39557 );
   nand U45746 ( n44051,n28360,p2_ebx_reg_31_ );
   and U45747 ( n42657,n42826,n44605 );
   nand U45748 ( n44605,n44606,n44607 );
   nand U45749 ( n44607,n44608,n39455 );
   nor U45750 ( n44608,p2_ebx_reg_31_,n44048 );
   nand U45751 ( n44606,n39557,n44604 );
   not U45752 ( n44604,n37067 );
   nor U45753 ( n37067,n43907,n36647 );
   not U45754 ( n43907,n44048 );
   nor U45755 ( n44048,n37052,p2_statebs16_reg );
   nor U45756 ( n42826,n37217,n28122 );
   not U45757 ( n42652,n44609 );
   nor U45758 ( n44049,n36813,n44609 );
   nand U45759 ( n44609,n44610,n44611 );
   nor U45760 ( n44611,n37040,n44612 );
   not U45761 ( n44612,n37051 );
   nand U45762 ( n37051,n44613,n36642 );
   nor U45763 ( n36642,n36783,p2_state2_reg_2_ );
   nor U45764 ( n44613,p2_state2_reg_1_,n38681 );
   not U45765 ( n38681,p2_state2_reg_3_ );
   and U45766 ( n37040,n44614,n44615 );
   nor U45767 ( n44615,p2_statebs16_reg,p2_state2_reg_2_ );
   nor U45768 ( n44614,p2_state2_reg_0_,n28179 );
   nor U45769 ( n44610,n36629,n44616 );
   nor U45770 ( n44616,p2_state2_reg_0_,n36616 );
   not U45771 ( n36616,n39574 );
   not U45772 ( n36629,n36612 );
   nand U45773 ( n36612,n37045,n44617 );
   nand U45774 ( n44617,n44618,n44619 );
   nand U45775 ( n44619,n37213,n37215 );
   nand U45776 ( n37215,n37078,n44620 );
   nand U45777 ( n37078,n44621,n39467 );
   nand U45778 ( n44618,n37171,n37166 );
   not U45779 ( n37171,n37211 );
   nand U45780 ( n37211,n44621,n39530 );
   not U45781 ( n36813,p2_reip_reg_31_ );
   nand U45782 ( n44623,p2_byteenable_reg_3_,n44624 );
   nor U45783 ( n44622,n44625,n44626 );
   nor U45784 ( n44626,p2_reip_reg_1_,n44627 );
   nand U45785 ( n44629,p2_byteenable_reg_2_,n44624 );
   nor U45786 ( n44628,n44630,n44631 );
   nor U45787 ( n44631,n39602,n44632 );
   nor U45788 ( n44630,n44627,n44633 );
   nand U45789 ( n44633,n44634,n36961 );
   nand U45790 ( n44634,p2_datawidth_reg_0_,p2_reip_reg_0_ );
   not U45791 ( n44627,n44635 );
   nand U45792 ( n44637,p2_byteenable_reg_1_,n44624 );
   nor U45793 ( n44636,n44625,n44638 );
   and U45794 ( n44625,n44639,n44635 );
   nor U45795 ( n44635,n44624,p2_datawidth_reg_1_ );
   nor U45796 ( n44639,p2_reip_reg_0_,p2_datawidth_reg_0_ );
   not U45797 ( n44632,n44638 );
   nor U45798 ( n44638,n44624,n36961 );
   not U45799 ( n36961,p2_reip_reg_1_ );
   nor U45800 ( n44640,n44641,n44642 );
   nor U45801 ( n44642,n39602,n44624 );
   not U45802 ( n39602,p2_reip_reg_0_ );
   and U45803 ( n44641,n44624,p2_byteenable_reg_0_ );
   nand U45804 ( n44624,n44643,n44644 );
   nor U45805 ( n44644,n44645,n44646 );
   nand U45806 ( n44646,n44647,n44648 );
   nor U45807 ( n44648,n44649,n44650 );
   nand U45808 ( n44650,n37026,n37027 );
   not U45809 ( n37027,p2_datawidth_reg_29_ );
   not U45810 ( n37026,p2_datawidth_reg_28_ );
   nand U45811 ( n44649,n37000,n37028 );
   not U45812 ( n37028,p2_datawidth_reg_30_ );
   not U45813 ( n37000,p2_datawidth_reg_2_ );
   nor U45814 ( n44647,n44651,n44652 );
   nand U45815 ( n44652,n37022,n37023 );
   not U45816 ( n37023,p2_datawidth_reg_25_ );
   not U45817 ( n37022,p2_datawidth_reg_24_ );
   nand U45818 ( n44651,n37024,n37025 );
   not U45819 ( n37025,p2_datawidth_reg_27_ );
   not U45820 ( n37024,p2_datawidth_reg_26_ );
   nand U45821 ( n44645,n44653,n44654 );
   nor U45822 ( n44654,n44655,n44656 );
   nand U45823 ( n44656,n37004,n37005 );
   not U45824 ( n37005,p2_datawidth_reg_7_ );
   not U45825 ( n37004,p2_datawidth_reg_6_ );
   nand U45826 ( n44655,n37006,n37007 );
   not U45827 ( n37007,p2_datawidth_reg_9_ );
   not U45828 ( n37006,p2_datawidth_reg_8_ );
   nor U45829 ( n44653,n44657,n44658 );
   nand U45830 ( n44658,n37029,n37001 );
   not U45831 ( n37001,p2_datawidth_reg_3_ );
   not U45832 ( n37029,p2_datawidth_reg_31_ );
   nand U45833 ( n44657,n37002,n37003 );
   not U45834 ( n37003,p2_datawidth_reg_5_ );
   not U45835 ( n37002,p2_datawidth_reg_4_ );
   nor U45836 ( n44643,n44659,n44660 );
   nand U45837 ( n44660,n44661,n44662 );
   nor U45838 ( n44662,n44663,n44664 );
   nand U45839 ( n44664,n37010,n37011 );
   not U45840 ( n37011,p2_datawidth_reg_13_ );
   not U45841 ( n37010,p2_datawidth_reg_12_ );
   nand U45842 ( n44663,n37012,n37013 );
   not U45843 ( n37013,p2_datawidth_reg_15_ );
   not U45844 ( n37012,p2_datawidth_reg_14_ );
   nor U45845 ( n44661,n44665,n44666 );
   nand U45846 ( n44666,n37008,n37009 );
   not U45847 ( n37009,p2_datawidth_reg_11_ );
   not U45848 ( n37008,p2_datawidth_reg_10_ );
   and U45849 ( n44665,p2_datawidth_reg_1_,p2_datawidth_reg_0_ );
   nand U45850 ( n44659,n44667,n44668 );
   nor U45851 ( n44668,n44669,n44670 );
   nand U45852 ( n44670,n37018,n37019 );
   not U45853 ( n37019,p2_datawidth_reg_21_ );
   not U45854 ( n37018,p2_datawidth_reg_20_ );
   nand U45855 ( n44669,n37020,n37021 );
   not U45856 ( n37021,p2_datawidth_reg_23_ );
   not U45857 ( n37020,p2_datawidth_reg_22_ );
   nor U45858 ( n44667,n44671,n44672 );
   nand U45859 ( n44672,n37014,n37015 );
   not U45860 ( n37015,p2_datawidth_reg_17_ );
   not U45861 ( n37014,p2_datawidth_reg_16_ );
   nand U45862 ( n44671,n37016,n37017 );
   not U45863 ( n37017,p2_datawidth_reg_19_ );
   not U45864 ( n37016,p2_datawidth_reg_18_ );
   nand U45865 ( n44674,n44675,n37192 );
   nor U45866 ( n37192,n44676,n44677 );
   nand U45867 ( n44676,n38585,n28239 );
   nor U45868 ( n44675,n44678,n41036 );
   nor U45869 ( n44678,n44679,n44680 );
   nor U45870 ( n44680,n37201,n43891 );
   not U45871 ( n43891,n36650 );
   nand U45872 ( n37201,n44681,n44682 );
   nand U45873 ( n44682,p2_state2_reg_1_,n44683 );
   nand U45874 ( n44683,n44684,n44685 );
   nand U45875 ( n44685,n44686,p2_instqueuerd_addr_reg_3_ );
   nor U45876 ( n44686,p2_flush_reg,n44687 );
   nor U45877 ( n44687,n44688,n44689 );
   nor U45878 ( n44689,n37114,n44690 );
   nor U45879 ( n44688,n37120,n44691 );
   nand U45880 ( n44684,p2_instqueuerd_addr_reg_4_,n38712 );
   not U45881 ( n38712,p2_flush_reg );
   nand U45882 ( n44681,n44692,n28181 );
   nand U45883 ( n44692,n44693,n44694 );
   nand U45884 ( n44694,n44695,n44696 );
   not U45885 ( n44696,n44697 );
   nor U45886 ( n44695,n44698,n44699 );
   and U45887 ( n44698,n44691,n44690 );
   nand U45888 ( n44690,n44700,n44701 );
   nand U45889 ( n44701,n44702,n28180 );
   nand U45890 ( n44691,n44700,n44703 );
   nand U45891 ( n44703,n44704,n28179 );
   and U45892 ( n44700,n44705,n44706 );
   nand U45893 ( n44706,p2_state2_reg_1_,n37154 );
   nand U45894 ( n44705,n44707,n28178 );
   nor U45895 ( n44679,n37205,n44708 );
   nand U45896 ( n44708,n36644,n27896 );
   nand U45897 ( n37205,n44020,n44709 );
   nand U45898 ( n44709,n44710,n44013 );
   nor U45899 ( n44710,n44711,n44002 );
   not U45900 ( n44002,n44712 );
   nor U45901 ( n44711,n44713,n44005 );
   nor U45902 ( n44713,n40345,n44714 );
   not U45903 ( n44020,n44715 );
   nand U45904 ( n44673,p2_flush_reg,n36660 );
   not U45905 ( n36660,n36658 );
   nor U45906 ( n36658,n36787,n37075 );
   and U45907 ( n37075,n44716,n44717 );
   nor U45908 ( n44716,n44718,n44719 );
   nor U45909 ( n44719,n36615,n37052 );
   nor U45910 ( n36615,n39455,n39467 );
   and U45911 ( n44718,n39527,n37170 );
   nor U45912 ( n37170,n36647,n37052 );
   not U45913 ( n37052,n36635 );
   nand U45914 ( n36635,ready21_reg,ready12_reg );
   nand U45915 ( n36647,n44602,n36972 );
   and U45916 ( n44602,n36795,n44720 );
   nand U45917 ( n44720,p2_state_reg_2_,p2_state_reg_1_ );
   not U45918 ( n36795,n36799 );
   not U45919 ( n39527,n37194 );
   not U45920 ( n36787,n37045 );
   nor U45921 ( n44721,n44723,n44724 );
   nor U45922 ( n44724,n36648,n28167 );
   not U45923 ( n36648,p2_statebs16_reg );
   nor U45924 ( n44723,n28163,n28898 );
   nand U45925 ( n44722,n36799,n36972 );
   nor U45926 ( n36799,p2_state_reg_1_,p2_state_reg_2_ );
   nor U45927 ( n44725,n44726,n44727 );
   and U45928 ( n44727,n36619,p2_d_c_n_reg );
   nor U45929 ( n44726,p2_codefetch_reg,n36619 );
   not U45930 ( n36619,n36620 );
   nor U45931 ( n36620,n36973,p2_state_reg_0_ );
   nand U45932 ( n44729,p2_codefetch_reg,n44730 );
   nand U45933 ( n44730,n44717,n37045 );
   and U45934 ( n44717,n44731,n37187 );
   nand U45935 ( n37187,n44732,n44620 );
   nand U45936 ( n44620,n39456,n38680 );
   nand U45937 ( n44732,n44621,n39573 );
   nor U45938 ( n44621,n37113,n39569 );
   nor U45939 ( n44731,n44733,n44734 );
   nor U45940 ( n44734,n39505,n37166 );
   not U45941 ( n39505,n39530 );
   nor U45942 ( n44733,n39530,n37213 );
   nand U45943 ( n44728,n39574,p2_state2_reg_0_ );
   nand U45944 ( n44735,p2_ads_n_reg,p2_state_reg_0_ );
   nand U45945 ( n44736,n44737,p2_state_reg_0_ );
   nor U45946 ( n44737,p2_state_reg_2_,n36973 );
   nand U45947 ( n36987,n36972,n36973 );
   not U45948 ( n36973,p2_state_reg_1_ );
   not U45949 ( n36972,p2_state_reg_0_ );
   nand U45950 ( n44739,p2_memoryfetch_reg,n44740 );
   nand U45951 ( n44740,n44741,n44742 );
   nor U45952 ( n44742,n44743,n44744 );
   nor U45953 ( n44744,n39545,n37166 );
   nand U45954 ( n37166,n44745,n44746 );
   nand U45955 ( n44746,n44747,n44748 );
   not U45956 ( n44748,n44693 );
   nor U45957 ( n44747,n44749,n41037 );
   nor U45958 ( n44749,n44750,n44751 );
   nand U45959 ( n44745,n44750,n44751 );
   nand U45960 ( n44751,n44715,n36651 );
   nand U45961 ( n44715,n44045,n44752 );
   or U45962 ( n44752,n40500,n37132 );
   nand U45963 ( n40500,n44753,n44754 );
   nor U45964 ( n44754,n44755,n44756 );
   nand U45965 ( n44756,n44757,n44758 );
   nor U45966 ( n44758,n44759,n44760 );
   nor U45967 ( n44760,n40536,n44195 );
   nor U45968 ( n44759,n40533,n44196 );
   nor U45969 ( n44757,n44761,n44762 );
   nor U45970 ( n44762,n40546,n44199 );
   nor U45971 ( n44761,n40525,n44200 );
   nand U45972 ( n44755,n44763,n44764 );
   nor U45973 ( n44764,n44765,n44766 );
   nor U45974 ( n44766,n40524,n44205 );
   nor U45975 ( n44765,n40545,n44206 );
   nor U45976 ( n44763,n44767,n44768 );
   nor U45977 ( n44768,n40510,n44209 );
   nor U45978 ( n44767,n40511,n44210 );
   nor U45979 ( n44753,n44769,n44770 );
   nand U45980 ( n44770,n44771,n44772 );
   nor U45981 ( n44772,n44773,n44774 );
   nor U45982 ( n44774,n40514,n44217 );
   nor U45983 ( n44773,n40515,n44218 );
   nor U45984 ( n44771,n44775,n44776 );
   nor U45985 ( n44776,n40520,n44221 );
   nor U45986 ( n44775,n40521,n44222 );
   nand U45987 ( n44769,n44777,n44778 );
   nor U45988 ( n44778,n44779,n44780 );
   nor U45989 ( n44780,n38590,n44227 );
   nor U45990 ( n44779,n40541,n44228 );
   nor U45991 ( n44777,n44781,n44782 );
   nor U45992 ( n44782,n40532,n44231 );
   nor U45993 ( n44781,n40542,n44232 );
   nand U45994 ( n44045,n44783,n44784 );
   nand U45995 ( n44784,n44785,n44786 );
   or U45996 ( n44785,n44787,n44788 );
   nand U45997 ( n44783,n44788,n44787 );
   and U45998 ( n44750,n44789,n44790 );
   nand U45999 ( n44790,n44791,n44792 );
   nand U46000 ( n44791,n44793,n36651 );
   nand U46001 ( n44789,n44794,n44795 );
   nand U46002 ( n44795,n44796,n36651 );
   nand U46003 ( n44796,n44797,n44712 );
   xor U46004 ( n44712,n44798,n44799 );
   nand U46005 ( n44799,n44800,n44801 );
   xor U46006 ( n44798,n44802,n44803 );
   or U46007 ( n44797,n44792,n44013 );
   not U46008 ( n44013,n44793 );
   xor U46009 ( n44793,n44804,n44788 );
   and U46010 ( n44788,n44805,n44806 );
   nand U46011 ( n44806,n39455,n40798 );
   nand U46012 ( n40798,n44807,n44808 );
   nor U46013 ( n44808,n44809,n44810 );
   nand U46014 ( n44810,n44811,n44812 );
   nor U46015 ( n44812,n44813,n44814 );
   nor U46016 ( n44814,n40842,n44195 );
   nor U46017 ( n44813,n40839,n44196 );
   nor U46018 ( n44811,n44815,n44816 );
   nor U46019 ( n44816,n40853,n44199 );
   nor U46020 ( n44815,n40830,n44200 );
   nand U46021 ( n44809,n44817,n44818 );
   nor U46022 ( n44818,n44819,n44820 );
   nor U46023 ( n44820,n40828,n44205 );
   nor U46024 ( n44819,n40852,n44206 );
   nor U46025 ( n44817,n44821,n44822 );
   nor U46026 ( n44822,n40808,n44209 );
   nor U46027 ( n44821,n40811,n44210 );
   nor U46028 ( n44807,n44823,n44824 );
   nand U46029 ( n44824,n44825,n44826 );
   nor U46030 ( n44826,n44827,n44828 );
   nor U46031 ( n44828,n40816,n44217 );
   nor U46032 ( n44827,n40817,n44218 );
   nor U46033 ( n44825,n44829,n44830 );
   nor U46034 ( n44830,n40823,n44221 );
   nor U46035 ( n44829,n40825,n44222 );
   nand U46036 ( n44823,n44831,n44832 );
   nor U46037 ( n44832,n44833,n44834 );
   nor U46038 ( n44834,n38622,n44227 );
   nor U46039 ( n44833,n40848,n44228 );
   nor U46040 ( n44831,n44835,n44836 );
   nor U46041 ( n44836,n40838,n44231 );
   nor U46042 ( n44835,n40849,n44232 );
   nand U46043 ( n44805,p2_instqueuerd_addr_reg_4_,n44837 );
   xor U46044 ( n44804,n44787,n44786 );
   nand U46045 ( n44786,n44838,n37132 );
   nand U46046 ( n44838,p2_instqueuewr_addr_reg_4_,n44837 );
   nand U46047 ( n44787,n44839,n44840 );
   nand U46048 ( n44840,n44803,n44841 );
   nor U46049 ( n44839,n44842,n44843 );
   nor U46050 ( n44843,n44802,n44844 );
   nor U46051 ( n44844,n44841,n44803 );
   not U46052 ( n44802,n44845 );
   nor U46053 ( n44842,n44846,n44801 );
   nand U46054 ( n44801,n44847,n44848 );
   nor U46055 ( n44846,n44803,n44845 );
   nand U46056 ( n44845,n37132,n44849 );
   nand U46057 ( n44849,p2_instqueuewr_addr_reg_3_,n44837 );
   and U46058 ( n44803,n44850,n44851 );
   nand U46059 ( n44851,n39455,n40550 );
   nand U46060 ( n40550,n44852,n44853 );
   nor U46061 ( n44853,n44854,n44855 );
   nand U46062 ( n44855,n44856,n44857 );
   nor U46063 ( n44857,n44858,n44859 );
   nor U46064 ( n44859,n40574,n44195 );
   nor U46065 ( n44858,n40571,n44196 );
   nor U46066 ( n44856,n44860,n44861 );
   nor U46067 ( n44861,n40565,n44199 );
   nor U46068 ( n44860,n40586,n44200 );
   nand U46069 ( n44854,n44862,n44863 );
   nor U46070 ( n44863,n44864,n44865 );
   nor U46071 ( n44865,n40585,n44205 );
   nor U46072 ( n44864,n40564,n44206 );
   nor U46073 ( n44862,n44866,n44867 );
   nor U46074 ( n44867,n40591,n44209 );
   nor U46075 ( n44866,n40592,n44210 );
   nor U46076 ( n44852,n44868,n44869 );
   nand U46077 ( n44869,n44870,n44871 );
   nor U46078 ( n44871,n44872,n44873 );
   nor U46079 ( n44873,n40595,n44217 );
   nor U46080 ( n44872,n40596,n44218 );
   nor U46081 ( n44870,n44874,n44875 );
   nor U46082 ( n44875,n40581,n44221 );
   nor U46083 ( n44874,n40582,n44222 );
   nand U46084 ( n44868,n44876,n44877 );
   nor U46085 ( n44877,n44878,n44879 );
   nor U46086 ( n44879,n38638,n44227 );
   nor U46087 ( n44878,n40560,n44228 );
   nor U46088 ( n44876,n44880,n44881 );
   nor U46089 ( n44881,n40570,n44231 );
   nor U46090 ( n44880,n40561,n44232 );
   nand U46091 ( n44850,p2_instqueuerd_addr_reg_3_,n44837 );
   nand U46092 ( n44792,n44882,n44883 );
   nand U46093 ( n44883,n36644,n44697 );
   nand U46094 ( n44882,p2_instqueuerd_addr_reg_4_,n27895 );
   nand U46095 ( n44794,n44884,n44885 );
   nand U46096 ( n44885,n44886,n44005 );
   not U46097 ( n44005,n44887 );
   nor U46098 ( n44886,n40863,n38680 );
   nor U46099 ( n44884,n44888,n44889 );
   nor U46100 ( n44889,n44890,n44891 );
   nand U46101 ( n44891,n44892,n44893 );
   nand U46102 ( n44893,n44894,n44895 );
   nand U46103 ( n44892,n44896,n44897 );
   nand U46104 ( n44897,n44707,n36644 );
   nor U46105 ( n44896,n42873,n44898 );
   nor U46106 ( n44898,n38680,n44887 );
   nand U46107 ( n44887,n44899,n44900 );
   nand U46108 ( n44900,n44901,n44848 );
   nand U46109 ( n44901,n44800,n44847 );
   nand U46110 ( n44847,n44902,n44903 );
   not U46111 ( n44800,n44841 );
   nor U46112 ( n44841,n44903,n44902 );
   nand U46113 ( n44899,n44904,n44905 );
   xor U46114 ( n44905,n44903,n44902 );
   and U46115 ( n44902,n44906,n37132 );
   nand U46116 ( n44906,p2_instqueuewr_addr_reg_2_,n44837 );
   nand U46117 ( n44903,n44907,n44908 );
   nand U46118 ( n44908,n39455,n40700 );
   nand U46119 ( n40700,n44909,n44910 );
   nor U46120 ( n44910,n44911,n44912 );
   nand U46121 ( n44912,n44913,n44914 );
   nor U46122 ( n44914,n44915,n44916 );
   nor U46123 ( n44916,n40736,n44195 );
   nor U46124 ( n44915,n40733,n44196 );
   nor U46125 ( n44913,n44917,n44918 );
   nor U46126 ( n44918,n40746,n44199 );
   nor U46127 ( n44917,n40725,n44200 );
   nand U46128 ( n44911,n44919,n44920 );
   nor U46129 ( n44920,n44921,n44922 );
   nor U46130 ( n44922,n40724,n44205 );
   nor U46131 ( n44921,n40745,n44206 );
   nor U46132 ( n44919,n44923,n44924 );
   nor U46133 ( n44924,n40710,n44209 );
   nor U46134 ( n44923,n40711,n44210 );
   nor U46135 ( n44909,n44925,n44926 );
   nand U46136 ( n44926,n44927,n44928 );
   nor U46137 ( n44928,n44929,n44930 );
   nor U46138 ( n44930,n40714,n44217 );
   nor U46139 ( n44929,n40715,n44218 );
   nor U46140 ( n44927,n44931,n44932 );
   nor U46141 ( n44932,n40720,n44221 );
   nor U46142 ( n44931,n40721,n44222 );
   nand U46143 ( n44925,n44933,n44934 );
   nor U46144 ( n44934,n44935,n44936 );
   nor U46145 ( n44936,n38654,n44227 );
   nor U46146 ( n44935,n40741,n44228 );
   nor U46147 ( n44933,n44937,n44938 );
   nor U46148 ( n44938,n40732,n44231 );
   nor U46149 ( n44937,n40742,n44232 );
   nand U46150 ( n44907,p2_instqueuerd_addr_reg_2_,n44837 );
   not U46151 ( n44904,n44848 );
   nand U46152 ( n44848,n44939,n44940 );
   nand U46153 ( n44940,n44941,n44942 );
   nand U46154 ( n44941,n44943,n44944 );
   or U46155 ( n44939,n44944,n44943 );
   nor U46156 ( n44890,n44945,n44946 );
   nor U46157 ( n44946,n44947,n44948 );
   nor U46158 ( n44948,n44949,n42873 );
   and U46159 ( n44949,n44702,n36644 );
   nand U46160 ( n44702,n44950,n44951 );
   nand U46161 ( n44951,p2_instqueuewr_addr_reg_0_,n37114 );
   nor U46162 ( n44947,n36650,n44952 );
   nor U46163 ( n44952,n38680,n40345 );
   nand U46164 ( n40345,n44953,n44954 );
   nand U46165 ( n44954,n44955,p2_instqueuewr_addr_reg_0_ );
   and U46166 ( n44955,n37114,n44837 );
   nor U46167 ( n44953,n44956,n44957 );
   nor U46168 ( n44957,n37132,n40602 );
   nand U46169 ( n40602,n44958,n44959 );
   nor U46170 ( n44959,n44960,n44961 );
   nand U46171 ( n44961,n44962,n44963 );
   nor U46172 ( n44963,n44964,n44965 );
   nor U46173 ( n44965,n40638,n44195 );
   nor U46174 ( n44964,n40635,n44196 );
   nor U46175 ( n44962,n44966,n44967 );
   nor U46176 ( n44967,n40648,n44199 );
   nor U46177 ( n44966,n40627,n44200 );
   nand U46178 ( n44960,n44968,n44969 );
   nor U46179 ( n44969,n44970,n44971 );
   nor U46180 ( n44971,n40626,n44205 );
   nor U46181 ( n44970,n40647,n44206 );
   nor U46182 ( n44968,n44972,n44973 );
   nor U46183 ( n44973,n40612,n44209 );
   nor U46184 ( n44972,n40613,n44210 );
   nor U46185 ( n44958,n44974,n44975 );
   nand U46186 ( n44975,n44976,n44977 );
   nor U46187 ( n44977,n44978,n44979 );
   nor U46188 ( n44979,n40616,n44217 );
   nor U46189 ( n44978,n40617,n44218 );
   nor U46190 ( n44976,n44980,n44981 );
   nor U46191 ( n44981,n40622,n44221 );
   nor U46192 ( n44980,n40623,n44222 );
   nand U46193 ( n44974,n44982,n44983 );
   nor U46194 ( n44983,n44984,n44985 );
   nor U46195 ( n44985,n38693,n44227 );
   nor U46196 ( n44984,n40643,n44228 );
   nor U46197 ( n44982,n44986,n44987 );
   nor U46198 ( n44987,n40634,n44231 );
   nor U46199 ( n44986,n40644,n44232 );
   not U46200 ( n37132,n39455 );
   not U46201 ( n44956,n44942 );
   nor U46202 ( n36650,n41037,n39545 );
   not U46203 ( n41037,n36644 );
   nor U46204 ( n44945,n44895,n44894 );
   nor U46205 ( n44894,n44988,n44009 );
   not U46206 ( n44009,n44714 );
   xor U46207 ( n44714,n44989,n44943 );
   nor U46208 ( n44943,p2_instqueuewr_addr_reg_1_,n39455 );
   xor U46209 ( n44989,n44944,n44942 );
   nand U46210 ( n44942,n44990,n44837 );
   nand U46211 ( n44944,n44991,n44992 );
   nand U46212 ( n44992,n39455,n40651 );
   nand U46213 ( n40651,n44993,n44994 );
   nor U46214 ( n44994,n44995,n44996 );
   nand U46215 ( n44996,n44997,n44998 );
   nor U46216 ( n44998,n44999,n45000 );
   nor U46217 ( n45000,n40687,n44195 );
   nand U46218 ( n44195,n45001,n42441 );
   nor U46219 ( n44999,n40684,n44196 );
   nand U46220 ( n44196,n45001,n42419 );
   nor U46221 ( n44997,n45002,n45003 );
   nor U46222 ( n45003,n40697,n44199 );
   nand U46223 ( n44199,n45001,n42416 );
   nor U46224 ( n45002,n40676,n44200 );
   nand U46225 ( n44200,n42441,n45004 );
   nand U46226 ( n44995,n45005,n45006 );
   nor U46227 ( n45006,n45007,n45008 );
   nor U46228 ( n45008,n40675,n44205 );
   nand U46229 ( n44205,n42419,n45004 );
   nor U46230 ( n45007,n40696,n44206 );
   nand U46231 ( n44206,n42416,n45004 );
   nor U46232 ( n45005,n45009,n45010 );
   nor U46233 ( n45010,n40661,n44209 );
   nand U46234 ( n44209,n45011,n42419 );
   nor U46235 ( n45009,n40662,n44210 );
   nand U46236 ( n44210,n42441,n45011 );
   nor U46237 ( n44993,n45012,n45013 );
   nand U46238 ( n45013,n45014,n45015 );
   nor U46239 ( n45015,n45016,n45017 );
   nor U46240 ( n45017,n40665,n44217 );
   nand U46241 ( n44217,n42415,n45011 );
   nor U46242 ( n45016,n40666,n44218 );
   nand U46243 ( n44218,n45018,n42419 );
   nor U46244 ( n42419,n37126,n37114 );
   nor U46245 ( n45014,n45019,n45020 );
   nor U46246 ( n45020,n40671,n44221 );
   nand U46247 ( n44221,n45018,n42441 );
   nor U46248 ( n42441,n45021,p2_instqueuerd_addr_reg_0_ );
   nor U46249 ( n45019,n40672,n44222 );
   nand U46250 ( n44222,n45018,n42415 );
   nand U46251 ( n45012,n45022,n45023 );
   nor U46252 ( n45023,n45024,n45025 );
   nor U46253 ( n45025,n38669,n44227 );
   nand U46254 ( n44227,n42415,n45001 );
   nor U46255 ( n45001,n37178,n45026 );
   nor U46256 ( n45024,n40692,n44228 );
   nand U46257 ( n44228,n45011,n42416 );
   nor U46258 ( n45011,n37150,n37181 );
   nor U46259 ( n45022,n45027,n45028 );
   nor U46260 ( n45028,n40683,n44231 );
   nand U46261 ( n44231,n42415,n45004 );
   nor U46262 ( n45004,n45026,n37181 );
   not U46263 ( n45026,n37150 );
   nor U46264 ( n42415,n37114,n45021 );
   nor U46265 ( n45027,n40693,n44232 );
   nand U46266 ( n44232,n45018,n42416 );
   nor U46267 ( n42416,n37126,p2_instqueuerd_addr_reg_0_ );
   not U46268 ( n37126,n45021 );
   nor U46269 ( n45021,n44506,n42450 );
   nor U46270 ( n45018,n37178,n37150 );
   nand U46271 ( n37150,n45029,n45030 );
   or U46272 ( n45030,n42580,p2_instqueuerd_addr_reg_3_ );
   not U46273 ( n37178,n37181 );
   nor U46274 ( n37181,n45031,n42605 );
   nor U46275 ( n45031,n37154,n44506 );
   nor U46276 ( n39455,n39545,n39573 );
   nand U46277 ( n44991,p2_instqueuerd_addr_reg_1_,n44837 );
   nand U46278 ( n44837,n37194,n37136 );
   not U46279 ( n37136,n39467 );
   nor U46280 ( n39467,n28234,n28280 );
   nor U46281 ( n37194,n39530,n39557 );
   nor U46282 ( n39557,n36646,n39573 );
   not U46283 ( n44988,n36651 );
   nand U46284 ( n36651,n40863,n36655 );
   not U46285 ( n40863,n42873 );
   nor U46286 ( n42873,n36646,n36783 );
   and U46287 ( n44895,n36655,n45032 );
   nand U46288 ( n45032,n36644,n44704 );
   nand U46289 ( n36655,n39530,p2_state2_reg_0_ );
   nor U46290 ( n39530,n38680,n39545 );
   and U46291 ( n44888,n36644,n44699 );
   nor U46292 ( n36644,n36783,n39573 );
   not U46293 ( n39573,n38680 );
   not U46294 ( n39545,n36646 );
   nor U46295 ( n44743,n37213,n36646 );
   nand U46296 ( n36646,n45033,n45034 );
   nor U46297 ( n45034,n45035,n45036 );
   nand U46298 ( n45036,n45037,n45038 );
   nor U46299 ( n45038,n45039,n45040 );
   nor U46300 ( n45040,n45029,n40692 );
   not U46301 ( n40692,p2_instqueue_reg_15__1_ );
   nor U46302 ( n45039,n45041,n40671 );
   not U46303 ( n40671,p2_instqueue_reg_9__1_ );
   nor U46304 ( n45037,n45042,n45043 );
   nor U46305 ( n45043,n45044,n40675 );
   not U46306 ( n40675,p2_instqueue_reg_6__1_ );
   nor U46307 ( n45042,n45045,n40696 );
   not U46308 ( n40696,p2_instqueue_reg_7__1_ );
   nand U46309 ( n45035,n45046,n45047 );
   nor U46310 ( n45047,n45048,n45049 );
   nor U46311 ( n45049,n45050,n40665 );
   not U46312 ( n40665,p2_instqueue_reg_12__1_ );
   nor U46313 ( n45048,n45051,n40666 );
   not U46314 ( n40666,p2_instqueue_reg_10__1_ );
   nor U46315 ( n45046,n45052,n45053 );
   nor U46316 ( n45053,n45054,n40683 );
   not U46317 ( n40683,p2_instqueue_reg_4__1_ );
   nor U46318 ( n45052,n45055,n40684 );
   not U46319 ( n40684,p2_instqueue_reg_2__1_ );
   nor U46320 ( n45033,n45056,n45057 );
   nand U46321 ( n45057,n45058,n45059 );
   nor U46322 ( n45059,n45060,n45061 );
   nor U46323 ( n45061,n45062,n40687 );
   not U46324 ( n40687,p2_instqueue_reg_1__1_ );
   nor U46325 ( n45060,n45063,n40672 );
   not U46326 ( n40672,p2_instqueue_reg_8__1_ );
   nor U46327 ( n45058,n45064,n45065 );
   nor U46328 ( n45065,n45066,n38669 );
   not U46329 ( n38669,p2_instqueue_reg_0__1_ );
   nor U46330 ( n45064,n45067,n40693 );
   not U46331 ( n40693,p2_instqueue_reg_11__1_ );
   nand U46332 ( n45056,n45068,n45069 );
   nor U46333 ( n45069,n45070,n45071 );
   nor U46334 ( n45071,n45072,n40676 );
   not U46335 ( n40676,p2_instqueue_reg_5__1_ );
   nor U46336 ( n45070,n45073,n40661 );
   not U46337 ( n40661,p2_instqueue_reg_14__1_ );
   nor U46338 ( n45068,n45074,n45075 );
   nor U46339 ( n45075,n45076,n40697 );
   not U46340 ( n40697,p2_instqueue_reg_3__1_ );
   nor U46341 ( n45074,n45077,n40662 );
   not U46342 ( n40662,p2_instqueue_reg_13__1_ );
   nor U46343 ( n44741,n41036,n41202 );
   nand U46344 ( n41202,n45078,n45079 );
   nor U46345 ( n45079,n37113,n36783 );
   not U46346 ( n37113,n38649 );
   nor U46347 ( n45078,n38680,n39569 );
   nand U46348 ( n39569,n45080,n41715 );
   nor U46349 ( n41715,n39515,n39566 );
   and U46350 ( n45080,n43712,n37130 );
   nor U46351 ( n43712,n38617,n42814 );
   not U46352 ( n42814,n38601 );
   nor U46353 ( n44738,n39574,n45081 );
   nor U46354 ( n45081,n39549,n45082 );
   nand U46355 ( n45082,n37045,n38680 );
   nand U46356 ( n38680,n45083,n45084 );
   nor U46357 ( n45084,n45085,n45086 );
   nand U46358 ( n45086,n45087,n45088 );
   nor U46359 ( n45088,n45089,n45090 );
   nor U46360 ( n45090,n45029,n40643 );
   not U46361 ( n40643,p2_instqueue_reg_15__0_ );
   nor U46362 ( n45089,n45041,n40622 );
   not U46363 ( n40622,p2_instqueue_reg_9__0_ );
   nor U46364 ( n45087,n45091,n45092 );
   nor U46365 ( n45092,n45044,n40626 );
   not U46366 ( n40626,p2_instqueue_reg_6__0_ );
   nor U46367 ( n45091,n45045,n40647 );
   not U46368 ( n40647,p2_instqueue_reg_7__0_ );
   nand U46369 ( n45085,n45093,n45094 );
   nor U46370 ( n45094,n45095,n45096 );
   nor U46371 ( n45096,n45050,n40616 );
   not U46372 ( n40616,p2_instqueue_reg_12__0_ );
   nor U46373 ( n45095,n45051,n40617 );
   not U46374 ( n40617,p2_instqueue_reg_10__0_ );
   nor U46375 ( n45093,n45097,n45098 );
   nor U46376 ( n45098,n45054,n40634 );
   not U46377 ( n40634,p2_instqueue_reg_4__0_ );
   nor U46378 ( n45097,n45055,n40635 );
   not U46379 ( n40635,p2_instqueue_reg_2__0_ );
   nor U46380 ( n45083,n45099,n45100 );
   nand U46381 ( n45100,n45101,n45102 );
   nor U46382 ( n45102,n45103,n45104 );
   nor U46383 ( n45104,n45062,n40638 );
   not U46384 ( n40638,p2_instqueue_reg_1__0_ );
   nor U46385 ( n45103,n45063,n40623 );
   not U46386 ( n40623,p2_instqueue_reg_8__0_ );
   nor U46387 ( n45101,n45105,n45106 );
   nor U46388 ( n45106,n45066,n38693 );
   not U46389 ( n38693,p2_instqueue_reg_0__0_ );
   nor U46390 ( n45105,n45067,n40644 );
   not U46391 ( n40644,p2_instqueue_reg_11__0_ );
   nand U46392 ( n45099,n45107,n45108 );
   nor U46393 ( n45108,n45109,n45110 );
   nor U46394 ( n45110,n45072,n40627 );
   not U46395 ( n40627,p2_instqueue_reg_5__0_ );
   nor U46396 ( n45109,n45073,n40612 );
   not U46397 ( n40612,p2_instqueue_reg_14__0_ );
   nor U46398 ( n45107,n45111,n45112 );
   nor U46399 ( n45112,n45076,n40648 );
   not U46400 ( n40648,p2_instqueue_reg_3__0_ );
   nor U46401 ( n45111,n45077,n40613 );
   not U46402 ( n40613,p2_instqueue_reg_13__0_ );
   nor U46403 ( n37045,n36783,n41036 );
   not U46404 ( n41036,n37035 );
   nor U46405 ( n37035,n37217,p2_state2_reg_1_ );
   not U46406 ( n37217,p2_state2_reg_2_ );
   not U46407 ( n36783,p2_state2_reg_0_ );
   nand U46408 ( n39549,n37213,n39456 );
   not U46409 ( n39456,n41756 );
   nand U46410 ( n41756,n45113,n39515 );
   not U46411 ( n39515,n38585 );
   nand U46412 ( n38585,n45114,n45115 );
   nor U46413 ( n45115,n45116,n45117 );
   nand U46414 ( n45117,n45118,n45119 );
   nor U46415 ( n45119,n45120,n45121 );
   nor U46416 ( n45121,n45029,n40541 );
   not U46417 ( n40541,p2_instqueue_reg_15__6_ );
   nor U46418 ( n45120,n45041,n40520 );
   not U46419 ( n40520,p2_instqueue_reg_9__6_ );
   nor U46420 ( n45118,n45122,n45123 );
   nor U46421 ( n45123,n45044,n40524 );
   not U46422 ( n40524,p2_instqueue_reg_6__6_ );
   nor U46423 ( n45122,n45045,n40545 );
   not U46424 ( n40545,p2_instqueue_reg_7__6_ );
   nand U46425 ( n45116,n45124,n45125 );
   nor U46426 ( n45125,n45126,n45127 );
   nor U46427 ( n45127,n45050,n40514 );
   not U46428 ( n40514,p2_instqueue_reg_12__6_ );
   nor U46429 ( n45126,n45051,n40515 );
   not U46430 ( n40515,p2_instqueue_reg_10__6_ );
   nor U46431 ( n45124,n45128,n45129 );
   nor U46432 ( n45129,n45054,n40532 );
   not U46433 ( n40532,p2_instqueue_reg_4__6_ );
   nor U46434 ( n45128,n45055,n40533 );
   not U46435 ( n40533,p2_instqueue_reg_2__6_ );
   nor U46436 ( n45114,n45130,n45131 );
   nand U46437 ( n45131,n45132,n45133 );
   nor U46438 ( n45133,n45134,n45135 );
   nor U46439 ( n45135,n45062,n40536 );
   not U46440 ( n40536,p2_instqueue_reg_1__6_ );
   nor U46441 ( n45134,n45063,n40521 );
   not U46442 ( n40521,p2_instqueue_reg_8__6_ );
   nor U46443 ( n45132,n45136,n45137 );
   nor U46444 ( n45137,n45066,n38590 );
   not U46445 ( n38590,p2_instqueue_reg_0__6_ );
   nor U46446 ( n45136,n45067,n40542 );
   not U46447 ( n40542,p2_instqueue_reg_11__6_ );
   nand U46448 ( n45130,n45138,n45139 );
   nor U46449 ( n45139,n45140,n45141 );
   nor U46450 ( n45141,n45072,n40525 );
   not U46451 ( n40525,p2_instqueue_reg_5__6_ );
   nor U46452 ( n45140,n45073,n40510 );
   not U46453 ( n40510,p2_instqueue_reg_14__6_ );
   nor U46454 ( n45138,n45142,n45143 );
   nor U46455 ( n45143,n45076,n40546 );
   not U46456 ( n40546,p2_instqueue_reg_3__6_ );
   nor U46457 ( n45142,n45077,n40511 );
   not U46458 ( n40511,p2_instqueue_reg_13__6_ );
   nor U46459 ( n45113,n44677,n38601 );
   nand U46460 ( n38601,n45144,n45145 );
   nor U46461 ( n45145,n45146,n45147 );
   nand U46462 ( n45147,n45148,n45149 );
   nor U46463 ( n45149,n45150,n45151 );
   nor U46464 ( n45151,n45029,n40759 );
   not U46465 ( n40759,p2_instqueue_reg_15__5_ );
   nor U46466 ( n45150,n45041,n40780 );
   not U46467 ( n40780,p2_instqueue_reg_9__5_ );
   nor U46468 ( n45148,n45152,n45153 );
   nor U46469 ( n45153,n45044,n40784 );
   not U46470 ( n40784,p2_instqueue_reg_6__5_ );
   nor U46471 ( n45152,n45045,n40763 );
   not U46472 ( n40763,p2_instqueue_reg_7__5_ );
   nand U46473 ( n45146,n45154,n45155 );
   nor U46474 ( n45155,n45156,n45157 );
   nor U46475 ( n45157,n45050,n40794 );
   not U46476 ( n40794,p2_instqueue_reg_12__5_ );
   nor U46477 ( n45156,n45051,n40795 );
   not U46478 ( n40795,p2_instqueue_reg_10__5_ );
   nor U46479 ( n45154,n45158,n45159 );
   nor U46480 ( n45159,n45054,n40769 );
   not U46481 ( n40769,p2_instqueue_reg_4__5_ );
   nor U46482 ( n45158,n45055,n40770 );
   not U46483 ( n40770,p2_instqueue_reg_2__5_ );
   nor U46484 ( n45144,n45160,n45161 );
   nand U46485 ( n45161,n45162,n45163 );
   nor U46486 ( n45163,n45164,n45165 );
   nor U46487 ( n45165,n45062,n40773 );
   not U46488 ( n40773,p2_instqueue_reg_1__5_ );
   nor U46489 ( n45164,n45063,n40781 );
   not U46490 ( n40781,p2_instqueue_reg_8__5_ );
   nor U46491 ( n45162,n45166,n45167 );
   nor U46492 ( n45167,n45066,n38606 );
   not U46493 ( n38606,p2_instqueue_reg_0__5_ );
   nor U46494 ( n45166,n45067,n40760 );
   not U46495 ( n40760,p2_instqueue_reg_11__5_ );
   nand U46496 ( n45160,n45168,n45169 );
   nor U46497 ( n45169,n45170,n45171 );
   nor U46498 ( n45171,n45072,n40785 );
   not U46499 ( n40785,p2_instqueue_reg_5__5_ );
   nor U46500 ( n45170,n45073,n40790 );
   not U46501 ( n40790,p2_instqueue_reg_14__5_ );
   nor U46502 ( n45168,n45172,n45173 );
   nor U46503 ( n45173,n45076,n40764 );
   not U46504 ( n40764,p2_instqueue_reg_3__5_ );
   nor U46505 ( n45172,n45077,n40791 );
   not U46506 ( n40791,p2_instqueue_reg_13__5_ );
   nand U46507 ( n44677,n45174,n42622 );
   nor U46508 ( n42622,n37130,n39566 );
   not U46509 ( n39566,n38565 );
   nand U46510 ( n38565,n45175,n45176 );
   nor U46511 ( n45176,n45177,n45178 );
   nand U46512 ( n45178,n45179,n45180 );
   nor U46513 ( n45180,n45181,n45182 );
   nor U46514 ( n45182,n45029,n40492 );
   not U46515 ( n40492,p2_instqueue_reg_15__7_ );
   nor U46516 ( n45181,n45041,n40471 );
   not U46517 ( n40471,p2_instqueue_reg_9__7_ );
   nor U46518 ( n45179,n45183,n45184 );
   nor U46519 ( n45184,n45044,n40475 );
   not U46520 ( n40475,p2_instqueue_reg_6__7_ );
   nor U46521 ( n45183,n45045,n40496 );
   not U46522 ( n40496,p2_instqueue_reg_7__7_ );
   nand U46523 ( n45177,n45185,n45186 );
   nor U46524 ( n45186,n45187,n45188 );
   nor U46525 ( n45188,n45050,n40465 );
   not U46526 ( n40465,p2_instqueue_reg_12__7_ );
   nor U46527 ( n45187,n45051,n40466 );
   not U46528 ( n40466,p2_instqueue_reg_10__7_ );
   nor U46529 ( n45185,n45189,n45190 );
   nor U46530 ( n45190,n45054,n40483 );
   not U46531 ( n40483,p2_instqueue_reg_4__7_ );
   nor U46532 ( n45189,n45055,n40484 );
   not U46533 ( n40484,p2_instqueue_reg_2__7_ );
   nor U46534 ( n45175,n45191,n45192 );
   nand U46535 ( n45192,n45193,n45194 );
   nor U46536 ( n45194,n45195,n45196 );
   nor U46537 ( n45196,n45062,n40487 );
   not U46538 ( n40487,p2_instqueue_reg_1__7_ );
   nor U46539 ( n45195,n45063,n40472 );
   not U46540 ( n40472,p2_instqueue_reg_8__7_ );
   nor U46541 ( n45193,n45197,n45198 );
   nor U46542 ( n45198,n45066,n38572 );
   not U46543 ( n38572,p2_instqueue_reg_0__7_ );
   nor U46544 ( n45197,n45067,n40493 );
   not U46545 ( n40493,p2_instqueue_reg_11__7_ );
   nand U46546 ( n45191,n45199,n45200 );
   nor U46547 ( n45200,n45201,n45202 );
   nor U46548 ( n45202,n45072,n40476 );
   not U46549 ( n40476,p2_instqueue_reg_5__7_ );
   nor U46550 ( n45201,n45073,n40461 );
   not U46551 ( n40461,p2_instqueue_reg_14__7_ );
   nor U46552 ( n45199,n45203,n45204 );
   nor U46553 ( n45204,n45076,n40497 );
   not U46554 ( n40497,p2_instqueue_reg_3__7_ );
   nor U46555 ( n45203,n45077,n40462 );
   not U46556 ( n40462,p2_instqueue_reg_13__7_ );
   not U46557 ( n37130,n38633 );
   nand U46558 ( n38633,n45205,n45206 );
   nor U46559 ( n45206,n45207,n45208 );
   nand U46560 ( n45208,n45209,n45210 );
   nor U46561 ( n45210,n45211,n45212 );
   nor U46562 ( n45212,n45029,n40560 );
   not U46563 ( n40560,p2_instqueue_reg_15__3_ );
   nor U46564 ( n45211,n45041,n40581 );
   not U46565 ( n40581,p2_instqueue_reg_9__3_ );
   nor U46566 ( n45209,n45213,n45214 );
   nor U46567 ( n45214,n45044,n40585 );
   not U46568 ( n40585,p2_instqueue_reg_6__3_ );
   nor U46569 ( n45213,n45045,n40564 );
   not U46570 ( n40564,p2_instqueue_reg_7__3_ );
   nand U46571 ( n45207,n45215,n45216 );
   nor U46572 ( n45216,n45217,n45218 );
   nor U46573 ( n45218,n45050,n40595 );
   not U46574 ( n40595,p2_instqueue_reg_12__3_ );
   nor U46575 ( n45217,n45051,n40596 );
   not U46576 ( n40596,p2_instqueue_reg_10__3_ );
   nor U46577 ( n45215,n45219,n45220 );
   nor U46578 ( n45220,n45054,n40570 );
   not U46579 ( n40570,p2_instqueue_reg_4__3_ );
   nor U46580 ( n45219,n45055,n40571 );
   not U46581 ( n40571,p2_instqueue_reg_2__3_ );
   nor U46582 ( n45205,n45221,n45222 );
   nand U46583 ( n45222,n45223,n45224 );
   nor U46584 ( n45224,n45225,n45226 );
   nor U46585 ( n45226,n45062,n40574 );
   not U46586 ( n40574,p2_instqueue_reg_1__3_ );
   nor U46587 ( n45225,n45063,n40582 );
   not U46588 ( n40582,p2_instqueue_reg_8__3_ );
   nor U46589 ( n45223,n45227,n45228 );
   nor U46590 ( n45228,n45066,n38638 );
   not U46591 ( n38638,p2_instqueue_reg_0__3_ );
   nor U46592 ( n45227,n45067,n40561 );
   not U46593 ( n40561,p2_instqueue_reg_11__3_ );
   nand U46594 ( n45221,n45229,n45230 );
   nor U46595 ( n45230,n45231,n45232 );
   nor U46596 ( n45232,n45072,n40586 );
   not U46597 ( n40586,p2_instqueue_reg_5__3_ );
   nor U46598 ( n45231,n45073,n40591 );
   not U46599 ( n40591,p2_instqueue_reg_14__3_ );
   nor U46600 ( n45229,n45233,n45234 );
   nor U46601 ( n45234,n45076,n40565 );
   not U46602 ( n40565,p2_instqueue_reg_3__3_ );
   nor U46603 ( n45233,n45077,n40592 );
   not U46604 ( n40592,p2_instqueue_reg_13__3_ );
   nor U46605 ( n45174,n38617,n38649 );
   nand U46606 ( n38649,n45235,n45236 );
   nor U46607 ( n45236,n45237,n45238 );
   nand U46608 ( n45238,n45239,n45240 );
   nor U46609 ( n45240,n45241,n45242 );
   nor U46610 ( n45242,n45029,n40741 );
   not U46611 ( n40741,p2_instqueue_reg_15__2_ );
   nor U46612 ( n45241,n45041,n40720 );
   not U46613 ( n40720,p2_instqueue_reg_9__2_ );
   nor U46614 ( n45239,n45243,n45244 );
   nor U46615 ( n45244,n45044,n40724 );
   not U46616 ( n40724,p2_instqueue_reg_6__2_ );
   nor U46617 ( n45243,n45045,n40745 );
   not U46618 ( n40745,p2_instqueue_reg_7__2_ );
   nand U46619 ( n45237,n45245,n45246 );
   nor U46620 ( n45246,n45247,n45248 );
   nor U46621 ( n45248,n45050,n40714 );
   not U46622 ( n40714,p2_instqueue_reg_12__2_ );
   nor U46623 ( n45247,n45051,n40715 );
   not U46624 ( n40715,p2_instqueue_reg_10__2_ );
   nor U46625 ( n45245,n45249,n45250 );
   nor U46626 ( n45250,n45054,n40732 );
   not U46627 ( n40732,p2_instqueue_reg_4__2_ );
   nor U46628 ( n45249,n45055,n40733 );
   not U46629 ( n40733,p2_instqueue_reg_2__2_ );
   nor U46630 ( n45235,n45251,n45252 );
   nand U46631 ( n45252,n45253,n45254 );
   nor U46632 ( n45254,n45255,n45256 );
   nor U46633 ( n45256,n45062,n40736 );
   not U46634 ( n40736,p2_instqueue_reg_1__2_ );
   nor U46635 ( n45255,n45063,n40721 );
   not U46636 ( n40721,p2_instqueue_reg_8__2_ );
   nor U46637 ( n45253,n45257,n45258 );
   nor U46638 ( n45258,n45066,n38654 );
   not U46639 ( n38654,p2_instqueue_reg_0__2_ );
   nor U46640 ( n45257,n45067,n40742 );
   not U46641 ( n40742,p2_instqueue_reg_11__2_ );
   nand U46642 ( n45251,n45259,n45260 );
   nor U46643 ( n45260,n45261,n45262 );
   nor U46644 ( n45262,n45072,n40725 );
   not U46645 ( n40725,p2_instqueue_reg_5__2_ );
   nor U46646 ( n45261,n45073,n40710 );
   not U46647 ( n40710,p2_instqueue_reg_14__2_ );
   nor U46648 ( n45259,n45263,n45264 );
   nor U46649 ( n45264,n45076,n40746 );
   not U46650 ( n40746,p2_instqueue_reg_3__2_ );
   nor U46651 ( n45263,n45077,n40711 );
   not U46652 ( n40711,p2_instqueue_reg_13__2_ );
   nand U46653 ( n38617,n45265,n45266 );
   nor U46654 ( n45266,n45267,n45268 );
   nand U46655 ( n45268,n45269,n45270 );
   nor U46656 ( n45270,n45271,n45272 );
   nor U46657 ( n45272,n45029,n40848 );
   not U46658 ( n40848,p2_instqueue_reg_15__4_ );
   nand U46659 ( n45029,n42580,p2_instqueuerd_addr_reg_3_ );
   nor U46660 ( n45271,n45041,n40823 );
   not U46661 ( n40823,p2_instqueue_reg_9__4_ );
   nand U46662 ( n45041,n45273,n42582 );
   nor U46663 ( n45273,p2_instqueuerd_addr_reg_2_,n37139 );
   nor U46664 ( n45269,n45274,n45275 );
   nor U46665 ( n45275,n45044,n40828 );
   not U46666 ( n40828,p2_instqueue_reg_6__4_ );
   nand U46667 ( n45044,n42585,n37139 );
   nor U46668 ( n45274,n45045,n40852 );
   not U46669 ( n40852,p2_instqueue_reg_7__4_ );
   nand U46670 ( n45045,n42580,n37139 );
   nor U46671 ( n42580,n37155,n37154 );
   nand U46672 ( n45267,n45276,n45277 );
   nor U46673 ( n45277,n45278,n45279 );
   nor U46674 ( n45279,n45050,n40816 );
   not U46675 ( n40816,p2_instqueue_reg_12__4_ );
   nand U46676 ( n45050,n42592,p2_instqueuerd_addr_reg_3_ );
   nor U46677 ( n45278,n45051,n40817 );
   not U46678 ( n40817,p2_instqueue_reg_10__4_ );
   nand U46679 ( n45051,n42591,p2_instqueuerd_addr_reg_3_ );
   nor U46680 ( n45276,n45280,n45281 );
   nor U46681 ( n45281,n45054,n40838 );
   not U46682 ( n40838,p2_instqueue_reg_4__4_ );
   nand U46683 ( n45054,n42592,n37139 );
   nor U46684 ( n42592,n45282,n37154 );
   nor U46685 ( n45280,n45055,n40839 );
   not U46686 ( n40839,p2_instqueue_reg_2__4_ );
   nand U46687 ( n45055,n42591,n37139 );
   and U46688 ( n42591,n44530,n37154 );
   nor U46689 ( n44530,n37120,p2_instqueuerd_addr_reg_0_ );
   nor U46690 ( n45265,n45283,n45284 );
   nand U46691 ( n45284,n45285,n45286 );
   nor U46692 ( n45286,n45287,n45288 );
   nor U46693 ( n45288,n45062,n40842 );
   not U46694 ( n40842,p2_instqueue_reg_1__4_ );
   nand U46695 ( n45062,n45289,n42582 );
   nor U46696 ( n45289,p2_instqueuerd_addr_reg_3_,p2_instqueuerd_addr_reg_2_ );
   nor U46697 ( n45287,n45063,n40825 );
   not U46698 ( n40825,p2_instqueue_reg_8__4_ );
   nand U46699 ( n45063,n42449,p2_instqueuerd_addr_reg_3_ );
   nor U46700 ( n45285,n45290,n45291 );
   nor U46701 ( n45291,n45066,n38622 );
   not U46702 ( n38622,p2_instqueue_reg_0__4_ );
   nand U46703 ( n45066,n42449,n37139 );
   nor U46704 ( n42449,n45282,p2_instqueuerd_addr_reg_2_ );
   not U46705 ( n45282,n42450 );
   nor U46706 ( n42450,p2_instqueuerd_addr_reg_0_,p2_instqueuerd_addr_reg_1_ );
   nor U46707 ( n45290,n45067,n40849 );
   not U46708 ( n40849,p2_instqueue_reg_11__4_ );
   nand U46709 ( n45067,n42605,p2_instqueuerd_addr_reg_3_ );
   nand U46710 ( n45283,n45292,n45293 );
   nor U46711 ( n45293,n45294,n45295 );
   nor U46712 ( n45295,n45072,n40830 );
   not U46713 ( n40830,p2_instqueue_reg_5__4_ );
   nand U46714 ( n45072,n42610,n37139 );
   nor U46715 ( n45294,n45073,n40808 );
   not U46716 ( n40808,p2_instqueue_reg_14__4_ );
   nand U46717 ( n45073,n42585,p2_instqueuerd_addr_reg_3_ );
   nor U46718 ( n42585,n36779,p2_instqueuerd_addr_reg_0_ );
   nand U46719 ( n36779,p2_instqueuerd_addr_reg_2_,p2_instqueuerd_addr_reg_1_ );
   nor U46720 ( n45292,n45296,n45297 );
   nor U46721 ( n45297,n45076,n40853 );
   not U46722 ( n40853,p2_instqueue_reg_3__4_ );
   nand U46723 ( n45076,n42605,n37139 );
   nor U46724 ( n42605,n37155,p2_instqueuerd_addr_reg_2_ );
   not U46725 ( n37155,n44506 );
   nor U46726 ( n44506,n37120,n37114 );
   nor U46727 ( n45296,n45077,n40811 );
   not U46728 ( n40811,p2_instqueue_reg_13__4_ );
   nand U46729 ( n45077,n42610,p2_instqueuerd_addr_reg_3_ );
   nor U46730 ( n42610,n42602,n37154 );
   not U46731 ( n42602,n42582 );
   nor U46732 ( n42582,n37114,p2_instqueuerd_addr_reg_1_ );
   and U46733 ( n37213,n44693,n45298 );
   nand U46734 ( n45298,n45299,n45300 );
   nor U46735 ( n45300,n44697,n44707 );
   xor U46736 ( n44707,n45301,n45302 );
   xor U46737 ( n45301,n37607,n37154 );
   not U46738 ( n37154,p2_instqueuerd_addr_reg_2_ );
   xor U46739 ( n44697,n45303,n45304 );
   xor U46740 ( n45303,p2_instqueuewr_addr_reg_4_,p2_instqueuerd_addr_reg_4_ );
   nor U46741 ( n45299,n44699,n44704 );
   xor U46742 ( n44704,n45305,n44990 );
   xor U46743 ( n45305,n37096,n37120 );
   xor U46744 ( n44699,n45306,n45307 );
   xor U46745 ( n45306,n37606,n37139 );
   not U46746 ( n37139,p2_instqueuerd_addr_reg_3_ );
   nand U46747 ( n44693,n45308,n45309 );
   nand U46748 ( n45309,p2_instqueuewr_addr_reg_4_,n45310 );
   nand U46749 ( n45310,p2_instqueuerd_addr_reg_4_,n45304 );
   or U46750 ( n45308,n45304,p2_instqueuerd_addr_reg_4_ );
   nand U46751 ( n45304,n45311,n45312 );
   nand U46752 ( n45312,n45313,n37606 );
   not U46753 ( n37606,p2_instqueuewr_addr_reg_3_ );
   or U46754 ( n45313,n45307,p2_instqueuerd_addr_reg_3_ );
   nand U46755 ( n45311,p2_instqueuerd_addr_reg_3_,n45307 );
   nand U46756 ( n45307,n45314,n45315 );
   nand U46757 ( n45315,n45316,n37607 );
   not U46758 ( n37607,p2_instqueuewr_addr_reg_2_ );
   or U46759 ( n45316,n45302,p2_instqueuerd_addr_reg_2_ );
   nand U46760 ( n45314,p2_instqueuerd_addr_reg_2_,n45302 );
   nand U46761 ( n45302,n45317,n45318 );
   nand U46762 ( n45318,n45319,n37096 );
   not U46763 ( n37096,p2_instqueuewr_addr_reg_1_ );
   nand U46764 ( n45319,n37120,n44950 );
   not U46765 ( n44950,n44990 );
   not U46766 ( n37120,p2_instqueuerd_addr_reg_1_ );
   nand U46767 ( n45317,p2_instqueuerd_addr_reg_1_,n44990 );
   nor U46768 ( n44990,n37114,p2_instqueuewr_addr_reg_0_ );
   not U46769 ( n37114,p2_instqueuerd_addr_reg_0_ );
   nor U46770 ( n39574,n38704,p2_state2_reg_1_ );
   not U46771 ( n38704,n36628 );
   nor U46772 ( n36628,p2_state2_reg_2_,p2_state2_reg_3_ );
   nand U46773 ( n45321,n45322,p1_readrequest_reg );
   nand U46774 ( n45320,n45323,n45324 );
   not U46775 ( n45324,n45322 );
   nor U46776 ( n45322,n45325,n45326 );
   nand U46777 ( n45323,n45327,p1_state2_reg_2_ );
   nor U46778 ( n45327,n45328,n45329 );
   nand U46779 ( n45331,p1_m_io_n_reg,n28378 );
   nand U46780 ( n45330,p1_memoryfetch_reg,n45333 );
   or U46781 ( n45335,n45336,n45337 );
   nand U46782 ( n45334,n45338,n45336 );
   nand U46783 ( n45336,n45339,n45340 );
   nor U46784 ( n45340,n45341,n45342 );
   nor U46785 ( n45339,n45325,n45343 );
   nor U46786 ( n45343,n45344,n45345 );
   nand U46787 ( n45345,n45346,n28094 );
   nand U46788 ( n45338,n45348,n45349 );
   nand U46789 ( n45349,n45350,n45351 );
   nor U46790 ( n45348,n45352,n45353 );
   nor U46791 ( n45353,n45354,n45347 );
   nor U46792 ( n45354,n45355,n45356 );
   nand U46793 ( n45356,n45357,n45346 );
   nand U46794 ( n45357,n45358,n45359 );
   nand U46795 ( n45359,p1_statebs16_reg,n45360 );
   nand U46796 ( n45362,n45363,n45364 );
   not U46797 ( n45363,n45365 );
   nand U46798 ( n45361,p1_more_reg,n45365 );
   or U46799 ( n45367,n45332,p1_readrequest_reg );
   nand U46800 ( n45366,p1_w_r_n_reg,n28378 );
   nor U46801 ( n45368,n45370,n45371 );
   nor U46802 ( n45371,n45372,n45373 );
   and U46803 ( n45370,n45372,p1_byteenable_reg_0_ );
   nand U46804 ( n45375,n45376,p1_reip_reg_0_ );
   nor U46805 ( n45374,n45377,n45378 );
   nor U46806 ( n45378,n45372,n45379 );
   nand U46807 ( n45379,n45380,n45381 );
   nand U46808 ( n45381,p1_reip_reg_0_,p1_datawidth_reg_0_ );
   nor U46809 ( n45380,p1_reip_reg_1_,p1_datawidth_reg_1_ );
   and U46810 ( n45377,n45372,p1_byteenable_reg_2_ );
   nand U46811 ( n45383,n45384,p1_instqueuewr_addr_reg_0_ );
   nand U46812 ( n45382,n45385,n45386 );
   nand U46813 ( n45385,n45387,n45388 );
   nand U46814 ( n45388,n45341,n45389 );
   nor U46815 ( n45387,n45390,n45391 );
   nor U46816 ( n45391,n45344,n45392 );
   nor U46817 ( n45390,n45393,n45394 );
   nand U46818 ( n45396,n45384,p1_instqueuewr_addr_reg_1_ );
   nand U46819 ( n45395,n45397,n45386 );
   nand U46820 ( n45397,n45398,n45399 );
   nand U46821 ( n45399,n45400,n45401 );
   nor U46822 ( n45398,n45402,n45403 );
   nor U46823 ( n45403,n45393,n45404 );
   nor U46824 ( n45402,n45405,n45406 );
   nor U46825 ( n45405,n45407,n45408 );
   nand U46826 ( n45410,n45384,p1_instqueuewr_addr_reg_2_ );
   nand U46827 ( n45409,n45411,n45386 );
   nand U46828 ( n45411,n45412,n45413 );
   nand U46829 ( n45413,n45400,n45414 );
   nor U46830 ( n45412,n45415,n45416 );
   nor U46831 ( n45416,n45393,n45417 );
   nor U46832 ( n45415,n45406,n45418 );
   nand U46833 ( n45418,n45419,n45420 );
   or U46834 ( n45419,n45421,n45422 );
   nand U46835 ( n45424,n45384,p1_instqueuewr_addr_reg_3_ );
   nand U46836 ( n45423,n45425,n45386 );
   nand U46837 ( n45425,n45426,n45427 );
   nand U46838 ( n45427,n45428,n45400 );
   nor U46839 ( n45426,n45429,n45430 );
   nor U46840 ( n45430,n45393,n45431 );
   nor U46841 ( n45393,n45432,p1_state2_reg_3_ );
   nor U46842 ( n45429,n45433,n45406 );
   nor U46843 ( n45433,n45434,n45435 );
   nor U46844 ( n45434,n45436,n45437 );
   nand U46845 ( n45439,p1_instqueuerd_addr_reg_0_,n45440 );
   nand U46846 ( n45440,n45441,n45442 );
   nand U46847 ( n45442,n45443,n45444 );
   nand U46848 ( n45438,n45445,n45441 );
   nand U46849 ( n45445,n45446,n45447 );
   nand U46850 ( n45447,p1_state2_reg_1_,n45448 );
   nor U46851 ( n45446,n45449,n45450 );
   and U46852 ( n45450,n45451,n45452 );
   and U46853 ( n45449,n45453,n45443 );
   nand U46854 ( n45455,n45456,p1_instqueuerd_addr_reg_1_ );
   nand U46855 ( n45454,n45457,n45441 );
   nand U46856 ( n45457,n45458,n45459 );
   nand U46857 ( n45459,n45452,n45460 );
   nor U46858 ( n45458,n45461,n45462 );
   nor U46859 ( n45462,n45463,n45464 );
   nor U46860 ( n45461,n45448,n45465 );
   nand U46861 ( n45465,p1_state2_reg_1_,n45466 );
   nand U46862 ( n45468,n45456,p1_instqueuerd_addr_reg_2_ );
   nand U46863 ( n45467,n45469,n45441 );
   nand U46864 ( n45469,n45470,n45471 );
   nand U46865 ( n45471,n45452,n45472 );
   nor U46866 ( n45470,n45473,n45474 );
   nor U46867 ( n45474,n45475,n45464 );
   nor U46868 ( n45473,n45466,n45476 );
   nand U46869 ( n45476,p1_instaddrpointer_reg_0_,p1_state2_reg_1_ );
   nand U46870 ( n45466,n45477,n45478 );
   nand U46871 ( n45478,n45479,n45480 );
   nand U46872 ( n45477,p1_instaddrpointer_reg_31_,n45481 );
   nand U46873 ( n45483,n45456,p1_instqueuerd_addr_reg_3_ );
   nand U46874 ( n45482,n45484,n45441 );
   nand U46875 ( n45484,n45485,n45486 );
   nand U46876 ( n45486,n45443,n45487 );
   nand U46877 ( n45485,n45452,n45488 );
   nand U46878 ( n45490,n45491,n45441 );
   nor U46879 ( n45491,n45464,n45492 );
   nand U46880 ( n45489,n45456,p1_instqueuerd_addr_reg_4_ );
   not U46881 ( n45456,n45441 );
   nand U46882 ( n45441,n45493,n45494 );
   nand U46883 ( n45494,p1_state2_reg_3_,n45347 );
   nor U46884 ( n45493,n45495,n45496 );
   nor U46885 ( n45496,n45497,n45498 );
   or U46886 ( n45500,n45501,n45502 );
   nand U46887 ( n45499,n45502,n45503 );
   nand U46888 ( n45505,n45506,p1_datawidth_reg_1_ );
   nand U46889 ( n45504,n45507,n28156 );
   nand U46890 ( n45507,n28898,n45509 );
   nand U46891 ( n45511,n45512,n45508 );
   nor U46892 ( n45512,bs16,n45513 );
   nand U46893 ( n45510,n45506,p1_datawidth_reg_0_ );
   nand U46894 ( n45515,p1_be_n_reg_0_,n45332 );
   nand U46895 ( n45514,p1_byteenable_reg_0_,n45333 );
   nand U46896 ( n45517,p1_be_n_reg_1_,n45332 );
   nand U46897 ( n45516,p1_byteenable_reg_1_,n45333 );
   nand U46898 ( n45519,p1_be_n_reg_2_,n28378 );
   nand U46899 ( n45518,p1_byteenable_reg_2_,n45333 );
   nand U46900 ( n45521,p1_be_n_reg_3_,n28378 );
   nand U46901 ( n45520,p1_byteenable_reg_3_,n45333 );
   nand U46902 ( n45523,p1_address_reg_29_,n28378 );
   nor U46903 ( n45522,n45524,n45525 );
   nor U46904 ( n45525,n28137,n45527 );
   nor U46905 ( n45524,n45528,n45529 );
   nand U46906 ( n45531,p1_address_reg_28_,n28378 );
   nor U46907 ( n45530,n45532,n45533 );
   nor U46908 ( n45533,n45529,n28138 );
   nor U46909 ( n45532,n28393,n45534 );
   nand U46910 ( n45536,p1_address_reg_27_,n45332 );
   nor U46911 ( n45535,n45537,n45538 );
   nor U46912 ( n45538,n28138,n45534 );
   nor U46913 ( n45537,n45528,n45539 );
   nand U46914 ( n45541,p1_address_reg_26_,n28378 );
   nor U46915 ( n45540,n45542,n45543 );
   nor U46916 ( n45543,n45526,n45539 );
   nor U46917 ( n45542,n28394,n45544 );
   nand U46918 ( n45546,p1_address_reg_25_,n28378 );
   nor U46919 ( n45545,n45547,n45548 );
   nor U46920 ( n45548,n28137,n45544 );
   nor U46921 ( n45547,n28393,n45549 );
   nand U46922 ( n45551,p1_address_reg_24_,n28378 );
   nor U46923 ( n45550,n45552,n45553 );
   nor U46924 ( n45553,n28138,n45549 );
   nor U46925 ( n45552,n28393,n45554 );
   nand U46926 ( n45556,p1_address_reg_23_,n28378 );
   nor U46927 ( n45555,n45557,n45558 );
   nor U46928 ( n45558,n45526,n45554 );
   nor U46929 ( n45557,n45528,n45559 );
   nand U46930 ( n45561,p1_address_reg_22_,n28378 );
   nor U46931 ( n45560,n45562,n45563 );
   nor U46932 ( n45563,n45526,n45559 );
   nor U46933 ( n45562,n28394,n45564 );
   nand U46934 ( n45566,p1_address_reg_21_,n28378 );
   nor U46935 ( n45565,n45567,n45568 );
   nor U46936 ( n45568,n28137,n45564 );
   nor U46937 ( n45567,n28393,n45569 );
   nand U46938 ( n45571,p1_address_reg_20_,n45332 );
   nor U46939 ( n45570,n45572,n45573 );
   nor U46940 ( n45573,n28138,n45569 );
   nor U46941 ( n45572,n45528,n45574 );
   nand U46942 ( n45576,p1_address_reg_19_,n28378 );
   nor U46943 ( n45575,n45577,n45578 );
   nor U46944 ( n45578,n45526,n45574 );
   nor U46945 ( n45577,n28394,n45579 );
   nand U46946 ( n45581,p1_address_reg_18_,n45332 );
   nor U46947 ( n45580,n45582,n45583 );
   nor U46948 ( n45583,n28137,n45579 );
   nor U46949 ( n45582,n28393,n45584 );
   nand U46950 ( n45586,p1_address_reg_17_,n28378 );
   nor U46951 ( n45585,n45587,n45588 );
   nor U46952 ( n45588,n28138,n45584 );
   nor U46953 ( n45587,n45528,n45589 );
   nand U46954 ( n45591,p1_address_reg_16_,n28378 );
   nor U46955 ( n45590,n45592,n45593 );
   nor U46956 ( n45593,n45526,n45589 );
   nor U46957 ( n45592,n28394,n45594 );
   nand U46958 ( n45596,p1_address_reg_15_,n28378 );
   nor U46959 ( n45595,n45597,n45598 );
   nor U46960 ( n45598,n28137,n45594 );
   nor U46961 ( n45597,n28394,n45599 );
   nand U46962 ( n45601,p1_address_reg_14_,n28378 );
   nor U46963 ( n45600,n45602,n45603 );
   nor U46964 ( n45603,n28138,n45599 );
   nor U46965 ( n45602,n28394,n45604 );
   nand U46966 ( n45606,p1_address_reg_13_,n28378 );
   nor U46967 ( n45605,n45607,n45608 );
   nor U46968 ( n45608,n28137,n45604 );
   nor U46969 ( n45607,n45528,n45609 );
   nand U46970 ( n45611,p1_address_reg_12_,n45332 );
   nor U46971 ( n45610,n45612,n45613 );
   nor U46972 ( n45613,n45526,n45609 );
   nor U46973 ( n45612,n28393,n45614 );
   nand U46974 ( n45616,p1_address_reg_11_,n28378 );
   nor U46975 ( n45615,n45617,n45618 );
   nor U46976 ( n45618,n45526,n45614 );
   nor U46977 ( n45617,n28393,n45619 );
   nand U46978 ( n45621,p1_address_reg_10_,n28378 );
   nor U46979 ( n45620,n45622,n45623 );
   nor U46980 ( n45623,n28137,n45619 );
   nor U46981 ( n45622,n45528,n45624 );
   nand U46982 ( n45626,p1_address_reg_9_,n45332 );
   nor U46983 ( n45625,n45627,n45628 );
   nor U46984 ( n45628,n28138,n45624 );
   nor U46985 ( n45627,n28394,n45629 );
   nand U46986 ( n45631,p1_address_reg_8_,n45332 );
   nor U46987 ( n45630,n45632,n45633 );
   nor U46988 ( n45633,n45526,n45629 );
   nor U46989 ( n45632,n28393,n45634 );
   nand U46990 ( n45636,p1_address_reg_7_,n28378 );
   nor U46991 ( n45635,n45637,n45638 );
   nor U46992 ( n45638,n28137,n45634 );
   nor U46993 ( n45637,n45528,n45639 );
   nand U46994 ( n45641,p1_address_reg_6_,n45332 );
   nor U46995 ( n45640,n45642,n45643 );
   nor U46996 ( n45643,n28138,n45639 );
   nor U46997 ( n45642,n28394,n45644 );
   nand U46998 ( n45646,p1_address_reg_5_,n28378 );
   nor U46999 ( n45645,n45647,n45648 );
   nor U47000 ( n45648,n45526,n45644 );
   nor U47001 ( n45647,n28393,n45649 );
   nand U47002 ( n45651,p1_address_reg_4_,n45332 );
   nor U47003 ( n45650,n45652,n45653 );
   nor U47004 ( n45653,n28137,n45649 );
   nor U47005 ( n45652,n45528,n45654 );
   nand U47006 ( n45656,p1_address_reg_3_,n45332 );
   nor U47007 ( n45655,n45657,n45658 );
   nor U47008 ( n45658,n28138,n45654 );
   nor U47009 ( n45657,n28394,n45659 );
   nand U47010 ( n45661,p1_address_reg_2_,n45332 );
   nor U47011 ( n45660,n45662,n45663 );
   nor U47012 ( n45663,n45526,n45659 );
   nor U47013 ( n45662,n28393,n45664 );
   nand U47014 ( n45666,p1_address_reg_1_,n28378 );
   nor U47015 ( n45665,n45667,n45668 );
   nor U47016 ( n45668,n28137,n45664 );
   nor U47017 ( n45667,n45528,n45669 );
   nand U47018 ( n45671,p1_address_reg_0_,n45332 );
   nor U47019 ( n45670,n45672,n45673 );
   nor U47020 ( n45673,n28138,n45669 );
   nor U47021 ( n45672,n45674,n28394 );
   not U47022 ( n45528,n45675 );
   nand U47023 ( n45677,n45678,n45679 );
   nor U47024 ( n45679,n45680,n45681 );
   nor U47025 ( n45681,p1_requestpending_reg,hold );
   nor U47026 ( n45680,n45682,n45683 );
   nor U47027 ( n45682,p1_requestpending_reg,n45509 );
   nor U47028 ( n45678,n45684,n45685 );
   nor U47029 ( n45684,n29075,n45686 );
   nor U47030 ( n45676,n45675,n45687 );
   nor U47031 ( n45687,n45688,n45689 );
   nor U47032 ( n45688,n45683,n45690 );
   nand U47033 ( n45690,n45691,n45692 );
   nand U47034 ( n45692,n29075,n45685 );
   not U47035 ( n29075,na );
   nand U47036 ( n45691,p1_state_reg_0_,hold );
   nor U47037 ( n45683,n45686,n45346 );
   nor U47038 ( n45675,n45689,n45332 );
   nor U47039 ( n45694,n45695,n45696 );
   nand U47040 ( n45696,n45697,n28137 );
   nand U47041 ( n45526,n45333,n45689 );
   nand U47042 ( n45697,n45698,p1_state_reg_1_ );
   nor U47043 ( n45698,n45699,n45700 );
   nor U47044 ( n45700,n45701,n45702 );
   nand U47045 ( n45702,n29093,n45337 );
   nor U47046 ( n45699,n45703,n45689 );
   nor U47047 ( n45703,n45704,n45685 );
   nor U47048 ( n45704,n45701,n29093 );
   not U47049 ( n29093,hold );
   nor U47050 ( n45695,n45509,n45705 );
   nand U47051 ( n45705,p1_state_reg_0_,p1_requestpending_reg );
   nor U47052 ( n45693,n45706,n45707 );
   nor U47053 ( n45707,n45332,n45346 );
   nor U47054 ( n45706,n45708,n45689 );
   nor U47055 ( n45708,n45709,n45710 );
   and U47056 ( n45709,n45686,n45711 );
   nand U47057 ( n45713,n45710,na );
   nor U47058 ( n45712,n45714,n45715 );
   nor U47059 ( n45715,p1_state_reg_2_,n45716 );
   nor U47060 ( n45716,n45685,n45717 );
   nand U47061 ( n45717,p1_requestpending_reg,n45718 );
   nand U47062 ( n45718,n45701,p1_state_reg_1_ );
   nor U47063 ( n45714,n45711,n45719 );
   nand U47064 ( n45719,n45720,n45721 );
   nand U47065 ( n45721,n45686,n45689 );
   not U47066 ( n45689,p1_state_reg_2_ );
   nand U47067 ( n45720,p1_state_reg_1_,n45685 );
   nor U47068 ( n45711,n45337,hold );
   not U47069 ( n45337,p1_requestpending_reg );
   nor U47070 ( n53143,n28155,n45722 );
   nor U47071 ( n53144,n45508,n45723 );
   nor U47072 ( n53145,n28156,n45724 );
   nor U47073 ( n53146,n28155,n45725 );
   nor U47074 ( n53147,n45508,n45726 );
   nor U47075 ( n53148,n28156,n45727 );
   nor U47076 ( n53149,n28156,n45728 );
   nor U47077 ( n53150,n28155,n45729 );
   nor U47078 ( n53151,n45508,n45730 );
   nor U47079 ( n53152,n28156,n45731 );
   nor U47080 ( n53153,n28155,n45732 );
   nor U47081 ( n53154,n45508,n45733 );
   nor U47082 ( n53155,n28155,n45734 );
   nor U47083 ( n53156,n45508,n45735 );
   nor U47084 ( n53157,n45508,n45736 );
   nor U47085 ( n53158,n28155,n45737 );
   nor U47086 ( n53159,n28156,n45738 );
   nor U47087 ( n53160,n45508,n45739 );
   nor U47088 ( n53161,n28155,n45740 );
   nor U47089 ( n53162,n28156,n45741 );
   nor U47090 ( n53163,n28155,n45742 );
   nor U47091 ( n53164,n45508,n45743 );
   nor U47092 ( n53165,n28156,n45744 );
   nor U47093 ( n53166,n28155,n45745 );
   nor U47094 ( n53167,n45508,n45746 );
   nor U47095 ( n53168,n28156,n45747 );
   nor U47096 ( n53169,n28155,n45748 );
   nor U47097 ( n53170,n28156,n45750 );
   nor U47098 ( n45753,n45754,n45755 );
   nor U47099 ( n45755,n28094,n45756 );
   or U47100 ( n45756,n45757,n45701 );
   nor U47101 ( n45754,p1_state2_reg_0_,n45758 );
   nand U47102 ( n45758,p1_statebs16_reg,p1_state2_reg_1_ );
   nor U47103 ( n45752,n45759,n45760 );
   nor U47104 ( n45760,n45502,n28374 );
   nor U47105 ( n45502,n45347,n45761 );
   nand U47106 ( n45763,p1_state2_reg_1_,n45764 );
   nand U47107 ( n45764,n45765,n45766 );
   nor U47108 ( n45762,n45767,n45768 );
   nor U47109 ( n45768,n45761,n45769 );
   nor U47110 ( n45769,n45770,n45771 );
   nor U47111 ( n45770,n45701,n45772 );
   nor U47112 ( n45774,n45775,n45776 );
   nand U47113 ( n45776,n45766,n45777 );
   nand U47114 ( n45766,n45778,n45701 );
   nor U47115 ( n45778,p1_state2_reg_2_,n28094 );
   nor U47116 ( n45775,n45779,n45392 );
   not U47117 ( n45779,n45780 );
   nor U47118 ( n45773,n45781,n45782 );
   nand U47119 ( n45782,n45783,n45784 );
   nand U47120 ( n45784,n45785,n45347 );
   nor U47121 ( n45785,n45761,n45786 );
   and U47122 ( n45786,n45452,n45352 );
   nand U47123 ( n45783,n45761,p1_state2_reg_0_ );
   not U47124 ( n45761,n45765 );
   nand U47125 ( n45765,n45787,n45788 );
   nor U47126 ( n45788,n45789,n45790 );
   nor U47127 ( n45790,p1_state2_reg_0_,n45791 );
   nor U47128 ( n45791,n45432,n45346 );
   nor U47129 ( n45789,n45792,n28094 );
   nor U47130 ( n45792,p1_state2_reg_1_,n45793 );
   nor U47131 ( n45787,n45794,n45355 );
   nor U47132 ( n45794,n45795,n45796 );
   not U47133 ( n45796,n45797 );
   and U47134 ( n45781,n45793,n45771 );
   nand U47135 ( n45793,n45798,n45799 );
   nor U47136 ( n45799,n45800,n45801 );
   nand U47137 ( n45801,n45802,n45803 );
   nand U47138 ( n45802,n45804,n45805 );
   nand U47139 ( n45805,n45806,p1_instqueuewr_addr_reg_3_ );
   nor U47140 ( n45804,p1_instqueuewr_addr_reg_4_,n45807 );
   nor U47141 ( n45807,n45808,n45809 );
   nand U47142 ( n45809,n45810,n45811 );
   nand U47143 ( n45811,n45812,n45813 );
   nor U47144 ( n45812,p1_instqueuewr_addr_reg_2_,n45814 );
   nand U47145 ( n45810,n45815,n45816 );
   nand U47146 ( n45816,n45817,n45818 );
   nand U47147 ( n45818,n45819,n45820 );
   nand U47148 ( n45819,n45821,p1_instqueuewr_addr_reg_0_ );
   nor U47149 ( n45821,n45822,n45823 );
   nor U47150 ( n45823,n45497,n45463 );
   not U47151 ( n45463,n45824 );
   nor U47152 ( n45822,n45825,n45826 );
   nor U47153 ( n45817,n45827,n45828 );
   nor U47154 ( n45828,n45497,n45829 );
   nor U47155 ( n45829,n45830,n45453 );
   nand U47156 ( n45453,n45831,n45832 );
   nand U47157 ( n45832,n45833,n45451 );
   nand U47158 ( n45831,n45834,n45835 );
   nor U47159 ( n45830,n45451,n45836 );
   nor U47160 ( n45827,n45451,n45826 );
   nor U47161 ( n45815,n45837,n45838 );
   nor U47162 ( n45838,n45839,n45840 );
   nor U47163 ( n45839,n45841,n45814 );
   nor U47164 ( n45837,n45842,n45843 );
   nand U47165 ( n45843,n45844,n45845 );
   nand U47166 ( n45845,n45497,p1_instqueuerd_addr_reg_1_ );
   nand U47167 ( n45844,n45824,n45826 );
   nand U47168 ( n45824,n45846,n45847 );
   nand U47169 ( n45847,n45444,n45825 );
   nor U47170 ( n45846,n45848,n45849 );
   nor U47171 ( n45849,n45850,n45404 );
   and U47172 ( n45848,n45833,n45460 );
   nand U47173 ( n45833,n45851,n45852 );
   nand U47174 ( n45852,n45853,n45328 );
   nor U47175 ( n45808,p1_instqueuewr_addr_reg_3_,n45806 );
   not U47176 ( n45806,n45854 );
   nor U47177 ( n45800,n45855,n45856 );
   nor U47178 ( n45855,p1_flush_reg,p1_more_reg );
   nor U47179 ( n45798,n45364,n45857 );
   nand U47180 ( n45857,n45858,n45859 );
   nand U47181 ( n45859,n45860,n45861 );
   nand U47182 ( n45364,n45862,n45863 );
   nand U47183 ( n45863,n45864,n45865 );
   nor U47184 ( n45862,n45866,n45867 );
   nor U47185 ( n45867,n45868,n45869 );
   nor U47186 ( n45868,n45870,n45871 );
   nand U47187 ( n45871,n45872,n45836 );
   nand U47188 ( n45870,n45873,n45803 );
   nand U47189 ( n45803,n45874,n45875 );
   nor U47190 ( n45875,n45876,n45877 );
   nor U47191 ( n45874,n45878,n45879 );
   nor U47192 ( n45866,n45880,n45851 );
   nor U47193 ( n45882,n45883,n45884 );
   nand U47194 ( n45884,n45885,n45886 );
   nand U47195 ( n45886,n45887,n45888 );
   nand U47196 ( n45885,p1_instqueue_reg_15__7_,n45889 );
   nor U47197 ( n45883,n28192,n45891 );
   nor U47198 ( n45881,n45892,n45893 );
   nor U47199 ( n45893,n45894,n45895 );
   nor U47200 ( n45892,n45896,n28189 );
   nor U47201 ( n45899,n45900,n45901 );
   nand U47202 ( n45901,n45902,n45903 );
   nand U47203 ( n45903,n45904,n45888 );
   nand U47204 ( n45902,p1_instqueue_reg_15__6_,n45889 );
   nor U47205 ( n45900,n28198,n45891 );
   nor U47206 ( n45898,n45906,n45907 );
   nor U47207 ( n45907,n45908,n45895 );
   nor U47208 ( n45906,n45896,n28194 );
   nor U47209 ( n45911,n45912,n45913 );
   nand U47210 ( n45913,n45914,n45915 );
   nand U47211 ( n45915,n45916,n45888 );
   nand U47212 ( n45914,p1_instqueue_reg_15__5_,n45889 );
   nor U47213 ( n45912,n28204,n45891 );
   nor U47214 ( n45910,n45918,n45919 );
   nor U47215 ( n45919,n45920,n45895 );
   nor U47216 ( n45918,n45896,n28200 );
   nor U47217 ( n45923,n45924,n45925 );
   nand U47218 ( n45925,n45926,n45927 );
   nand U47219 ( n45927,n45928,n45888 );
   nand U47220 ( n45926,p1_instqueue_reg_15__4_,n45889 );
   nor U47221 ( n45924,n28211,n45891 );
   nor U47222 ( n45922,n45930,n45931 );
   nor U47223 ( n45931,n45932,n45895 );
   nor U47224 ( n45930,n45896,n28207 );
   nor U47225 ( n45935,n45936,n45937 );
   nand U47226 ( n45937,n45938,n45939 );
   nand U47227 ( n45939,n45940,n45888 );
   nand U47228 ( n45938,p1_instqueue_reg_15__3_,n45889 );
   nor U47229 ( n45936,n28219,n45891 );
   nor U47230 ( n45934,n45942,n45943 );
   nor U47231 ( n45943,n45944,n45895 );
   nor U47232 ( n45942,n45896,n28215 );
   nor U47233 ( n45947,n45948,n45949 );
   nand U47234 ( n45949,n45950,n45951 );
   nand U47235 ( n45951,n45952,n45888 );
   nand U47236 ( n45950,p1_instqueue_reg_15__2_,n45889 );
   nor U47237 ( n45948,n28231,n45891 );
   nor U47238 ( n45946,n45954,n45955 );
   nor U47239 ( n45955,n45956,n45895 );
   nor U47240 ( n45954,n45896,n28227 );
   nor U47241 ( n45959,n45960,n45961 );
   nand U47242 ( n45961,n45962,n45963 );
   nand U47243 ( n45963,n45964,n45888 );
   nand U47244 ( n45962,p1_instqueue_reg_15__1_,n45889 );
   nor U47245 ( n45960,n28249,n45891 );
   nor U47246 ( n45958,n45966,n45967 );
   nor U47247 ( n45967,n45968,n45895 );
   nor U47248 ( n45966,n45896,n28245 );
   nor U47249 ( n45971,n45972,n45973 );
   nand U47250 ( n45973,n45974,n45975 );
   nand U47251 ( n45975,n45976,n45888 );
   nand U47252 ( n45888,n45977,n45978 );
   nand U47253 ( n45978,p1_state2_reg_2_,n45979 );
   nand U47254 ( n45977,n45980,n45981 );
   nand U47255 ( n45974,p1_instqueue_reg_15__0_,n45889 );
   nand U47256 ( n45889,n45982,n45983 );
   nand U47257 ( n45983,p1_state2_reg_3_,n45896 );
   nor U47258 ( n45982,n45984,n45985 );
   nor U47259 ( n45985,n45986,n45987 );
   nand U47260 ( n45987,n45988,n45989 );
   nand U47261 ( n45988,n45990,n45991 );
   nand U47262 ( n45991,n45895,n45891 );
   and U47263 ( n45986,n45981,n45992 );
   nand U47264 ( n45981,n45896,n45993 );
   nand U47265 ( n45993,n45994,n45995 );
   nor U47266 ( n45984,n45355,n45979 );
   nand U47267 ( n45979,n45896,n45996 );
   nand U47268 ( n45996,n45997,n45998 );
   nor U47269 ( n45972,n28273,n45891 );
   nand U47270 ( n45891,n46000,n46001 );
   nor U47271 ( n45970,n46002,n46003 );
   nor U47272 ( n46003,n46004,n45895 );
   nand U47273 ( n45895,n45436,n46005 );
   not U47274 ( n45436,n45420 );
   nor U47275 ( n46002,n45896,n28325 );
   nand U47276 ( n45896,n46007,n46008 );
   nor U47277 ( n46010,n46011,n46012 );
   nand U47278 ( n46012,n46013,n46014 );
   nand U47279 ( n46014,n45887,n46015 );
   nand U47280 ( n46013,p1_instqueue_reg_14__7_,n46016 );
   nor U47281 ( n46011,n45890,n46017 );
   nor U47282 ( n46009,n46018,n46019 );
   nor U47283 ( n46019,n45894,n46020 );
   nor U47284 ( n46018,n28189,n46021 );
   nor U47285 ( n46023,n46024,n46025 );
   nand U47286 ( n46025,n46026,n46027 );
   nand U47287 ( n46027,n45904,n46015 );
   nand U47288 ( n46026,p1_instqueue_reg_14__6_,n46016 );
   nor U47289 ( n46024,n45905,n46017 );
   nor U47290 ( n46022,n46028,n46029 );
   nor U47291 ( n46029,n45908,n46020 );
   nor U47292 ( n46028,n28194,n46021 );
   nor U47293 ( n46031,n46032,n46033 );
   nand U47294 ( n46033,n46034,n46035 );
   nand U47295 ( n46035,n45916,n46015 );
   nand U47296 ( n46034,p1_instqueue_reg_14__5_,n46016 );
   nor U47297 ( n46032,n45917,n46017 );
   nor U47298 ( n46030,n46036,n46037 );
   nor U47299 ( n46037,n45920,n46020 );
   nor U47300 ( n46036,n28200,n46021 );
   nor U47301 ( n46039,n46040,n46041 );
   nand U47302 ( n46041,n46042,n46043 );
   nand U47303 ( n46043,n45928,n46015 );
   nand U47304 ( n46042,p1_instqueue_reg_14__4_,n46016 );
   nor U47305 ( n46040,n45929,n46017 );
   nor U47306 ( n46038,n46044,n46045 );
   nor U47307 ( n46045,n45932,n46020 );
   nor U47308 ( n46044,n28207,n46021 );
   nor U47309 ( n46047,n46048,n46049 );
   nand U47310 ( n46049,n46050,n46051 );
   nand U47311 ( n46051,n45940,n46015 );
   nand U47312 ( n46050,p1_instqueue_reg_14__3_,n46016 );
   nor U47313 ( n46048,n45941,n46017 );
   nor U47314 ( n46046,n46052,n46053 );
   nor U47315 ( n46053,n45944,n46020 );
   nor U47316 ( n46052,n28215,n46021 );
   nor U47317 ( n46055,n46056,n46057 );
   nand U47318 ( n46057,n46058,n46059 );
   nand U47319 ( n46059,n45952,n46015 );
   nand U47320 ( n46058,p1_instqueue_reg_14__2_,n46016 );
   nor U47321 ( n46056,n45953,n46017 );
   nor U47322 ( n46054,n46060,n46061 );
   nor U47323 ( n46061,n45956,n46020 );
   nor U47324 ( n46060,n28227,n46021 );
   nor U47325 ( n46063,n46064,n46065 );
   nand U47326 ( n46065,n46066,n46067 );
   nand U47327 ( n46067,n45964,n46015 );
   nand U47328 ( n46066,p1_instqueue_reg_14__1_,n46016 );
   nor U47329 ( n46064,n45965,n46017 );
   nor U47330 ( n46062,n46068,n46069 );
   nor U47331 ( n46069,n45968,n46020 );
   nor U47332 ( n46068,n28245,n46021 );
   nor U47333 ( n46071,n46072,n46073 );
   nand U47334 ( n46073,n46074,n46075 );
   nand U47335 ( n46075,n45976,n46015 );
   nand U47336 ( n46015,n46076,n46077 );
   nand U47337 ( n46077,n46078,n45998 );
   nand U47338 ( n46076,n46079,n45980 );
   not U47339 ( n46079,n46080 );
   nand U47340 ( n46074,p1_instqueue_reg_14__0_,n46016 );
   nand U47341 ( n46016,n46081,n46082 );
   nand U47342 ( n46082,p1_state2_reg_3_,n46021 );
   nor U47343 ( n46081,n46083,n46084 );
   nor U47344 ( n46084,n46085,n46086 );
   nand U47345 ( n46086,n46087,n45989 );
   nand U47346 ( n46087,n45990,n46088 );
   nand U47347 ( n46088,n46020,n46017 );
   nor U47348 ( n46085,n46080,n46089 );
   nand U47349 ( n46080,n45994,n46090 );
   nor U47350 ( n46083,n46091,n28374 );
   nor U47351 ( n46091,n46092,n46093 );
   nor U47352 ( n46072,n45999,n46017 );
   nand U47353 ( n46017,n46094,n46000 );
   nor U47354 ( n46070,n46095,n46096 );
   nor U47355 ( n46096,n46004,n46020 );
   nand U47356 ( n46020,n45407,n46097 );
   nor U47357 ( n46095,n28325,n46021 );
   nand U47358 ( n46021,n46098,n46007 );
   nor U47359 ( n46100,n46101,n46102 );
   nand U47360 ( n46102,n46103,n46104 );
   nand U47361 ( n46104,n45887,n46105 );
   nand U47362 ( n46103,p1_instqueue_reg_13__7_,n46106 );
   nor U47363 ( n46101,n28192,n46107 );
   nor U47364 ( n46099,n46108,n46109 );
   nor U47365 ( n46109,n28316,n46110 );
   nor U47366 ( n46108,n28189,n46111 );
   nor U47367 ( n46113,n46114,n46115 );
   nand U47368 ( n46115,n46116,n46117 );
   nand U47369 ( n46117,n45904,n46105 );
   nand U47370 ( n46116,p1_instqueue_reg_13__6_,n46106 );
   nor U47371 ( n46114,n28198,n46107 );
   nor U47372 ( n46112,n46118,n46119 );
   nor U47373 ( n46119,n28317,n46110 );
   nor U47374 ( n46118,n28194,n46111 );
   nor U47375 ( n46121,n46122,n46123 );
   nand U47376 ( n46123,n46124,n46125 );
   nand U47377 ( n46125,n45916,n46105 );
   nand U47378 ( n46124,p1_instqueue_reg_13__5_,n46106 );
   nor U47379 ( n46122,n28204,n46107 );
   nor U47380 ( n46120,n46126,n46127 );
   nor U47381 ( n46127,n28318,n46110 );
   nor U47382 ( n46126,n28200,n46111 );
   nor U47383 ( n46129,n46130,n46131 );
   nand U47384 ( n46131,n46132,n46133 );
   nand U47385 ( n46133,n45928,n46105 );
   nand U47386 ( n46132,p1_instqueue_reg_13__4_,n46106 );
   nor U47387 ( n46130,n28211,n46107 );
   nor U47388 ( n46128,n46134,n46135 );
   nor U47389 ( n46135,n28319,n46110 );
   nor U47390 ( n46134,n28207,n46111 );
   nor U47391 ( n46137,n46138,n46139 );
   nand U47392 ( n46139,n46140,n46141 );
   nand U47393 ( n46141,n45940,n46105 );
   nand U47394 ( n46140,p1_instqueue_reg_13__3_,n46106 );
   nor U47395 ( n46138,n28219,n46107 );
   nor U47396 ( n46136,n46142,n46143 );
   nor U47397 ( n46143,n28320,n46110 );
   nor U47398 ( n46142,n28215,n46111 );
   nor U47399 ( n46145,n46146,n46147 );
   nand U47400 ( n46147,n46148,n46149 );
   nand U47401 ( n46149,n45952,n46105 );
   nand U47402 ( n46148,p1_instqueue_reg_13__2_,n46106 );
   nor U47403 ( n46146,n28231,n46107 );
   nor U47404 ( n46144,n46150,n46151 );
   nor U47405 ( n46151,n28321,n46110 );
   nor U47406 ( n46150,n28227,n46111 );
   nor U47407 ( n46153,n46154,n46155 );
   nand U47408 ( n46155,n46156,n46157 );
   nand U47409 ( n46157,n45964,n46105 );
   nand U47410 ( n46156,p1_instqueue_reg_13__1_,n46106 );
   nor U47411 ( n46154,n28249,n46107 );
   nor U47412 ( n46152,n46158,n46159 );
   nor U47413 ( n46159,n28322,n46110 );
   nor U47414 ( n46158,n28245,n46111 );
   nor U47415 ( n46161,n46162,n46163 );
   nand U47416 ( n46163,n46164,n46165 );
   nand U47417 ( n46165,n45976,n46105 );
   nand U47418 ( n46105,n46166,n46167 );
   nand U47419 ( n46167,p1_state2_reg_2_,n46168 );
   nand U47420 ( n46166,n46169,n45980 );
   nand U47421 ( n46164,p1_instqueue_reg_13__0_,n46106 );
   nand U47422 ( n46106,n46170,n46171 );
   nand U47423 ( n46171,p1_state2_reg_3_,n46111 );
   nor U47424 ( n46170,n46172,n46173 );
   nor U47425 ( n46173,n46174,n46175 );
   nand U47426 ( n46175,n46176,n45989 );
   nand U47427 ( n46176,n45990,n46177 );
   nand U47428 ( n46177,n46110,n46107 );
   and U47429 ( n46174,n46169,n45992 );
   nand U47430 ( n46169,n46111,n46178 );
   nand U47431 ( n46178,n46179,n45994 );
   nor U47432 ( n46172,n28375,n46168 );
   nand U47433 ( n46168,n46111,n46180 );
   nand U47434 ( n46180,n46181,n45997 );
   nor U47435 ( n46162,n28273,n46107 );
   nand U47436 ( n46107,n46182,n46000 );
   nor U47437 ( n46160,n46183,n46184 );
   nor U47438 ( n46184,n28323,n46110 );
   nand U47439 ( n46110,n45408,n46097 );
   nor U47440 ( n46183,n28325,n46111 );
   nand U47441 ( n46111,n46185,n46007 );
   nor U47442 ( n46187,n46188,n46189 );
   nand U47443 ( n46189,n46190,n46191 );
   nand U47444 ( n46191,n45887,n46192 );
   nand U47445 ( n46190,p1_instqueue_reg_12__7_,n46193 );
   nor U47446 ( n46188,n28192,n46194 );
   nor U47447 ( n46186,n46195,n46196 );
   nor U47448 ( n46196,n28316,n46197 );
   nor U47449 ( n46195,n45897,n46198 );
   nor U47450 ( n46200,n46201,n46202 );
   nand U47451 ( n46202,n46203,n46204 );
   nand U47452 ( n46204,n45904,n46192 );
   nand U47453 ( n46203,p1_instqueue_reg_12__6_,n46193 );
   nor U47454 ( n46201,n28198,n46194 );
   nor U47455 ( n46199,n46205,n46206 );
   nor U47456 ( n46206,n28317,n46197 );
   nor U47457 ( n46205,n45909,n46198 );
   nor U47458 ( n46208,n46209,n46210 );
   nand U47459 ( n46210,n46211,n46212 );
   nand U47460 ( n46212,n45916,n46192 );
   nand U47461 ( n46211,p1_instqueue_reg_12__5_,n46193 );
   nor U47462 ( n46209,n28204,n46194 );
   nor U47463 ( n46207,n46213,n46214 );
   nor U47464 ( n46214,n28318,n46197 );
   nor U47465 ( n46213,n45921,n46198 );
   nor U47466 ( n46216,n46217,n46218 );
   nand U47467 ( n46218,n46219,n46220 );
   nand U47468 ( n46220,n45928,n46192 );
   nand U47469 ( n46219,p1_instqueue_reg_12__4_,n46193 );
   nor U47470 ( n46217,n28211,n46194 );
   nor U47471 ( n46215,n46221,n46222 );
   nor U47472 ( n46222,n28319,n46197 );
   nor U47473 ( n46221,n45933,n46198 );
   nor U47474 ( n46224,n46225,n46226 );
   nand U47475 ( n46226,n46227,n46228 );
   nand U47476 ( n46228,n45940,n46192 );
   nand U47477 ( n46227,p1_instqueue_reg_12__3_,n46193 );
   nor U47478 ( n46225,n28219,n46194 );
   nor U47479 ( n46223,n46229,n46230 );
   nor U47480 ( n46230,n28320,n46197 );
   nor U47481 ( n46229,n45945,n46198 );
   nor U47482 ( n46232,n46233,n46234 );
   nand U47483 ( n46234,n46235,n46236 );
   nand U47484 ( n46236,n45952,n46192 );
   nand U47485 ( n46235,p1_instqueue_reg_12__2_,n46193 );
   nor U47486 ( n46233,n28231,n46194 );
   nor U47487 ( n46231,n46237,n46238 );
   nor U47488 ( n46238,n28321,n46197 );
   nor U47489 ( n46237,n45957,n46198 );
   nor U47490 ( n46240,n46241,n46242 );
   nand U47491 ( n46242,n46243,n46244 );
   nand U47492 ( n46244,n45964,n46192 );
   nand U47493 ( n46243,p1_instqueue_reg_12__1_,n46193 );
   nor U47494 ( n46241,n28249,n46194 );
   nor U47495 ( n46239,n46245,n46246 );
   nor U47496 ( n46246,n28322,n46197 );
   nor U47497 ( n46245,n45969,n46198 );
   nor U47498 ( n46248,n46249,n46250 );
   nand U47499 ( n46250,n46251,n46252 );
   nand U47500 ( n46252,n45976,n46192 );
   nand U47501 ( n46192,n46253,n46254 );
   nand U47502 ( n46254,n46181,n46078 );
   nand U47503 ( n46253,n46255,n45980 );
   not U47504 ( n46255,n46256 );
   nand U47505 ( n46251,p1_instqueue_reg_12__0_,n46193 );
   nand U47506 ( n46193,n46257,n46258 );
   nand U47507 ( n46258,p1_state2_reg_3_,n46198 );
   nor U47508 ( n46257,n46259,n46260 );
   nor U47509 ( n46260,n46261,n46262 );
   nand U47510 ( n46262,n46263,n45989 );
   nand U47511 ( n46263,n45990,n46264 );
   nand U47512 ( n46264,n46197,n46194 );
   nor U47513 ( n46261,n46256,n46089 );
   nand U47514 ( n46256,n45994,n45404 );
   nor U47515 ( n45994,n45431,n45417 );
   nor U47516 ( n46259,n46265,n28374 );
   nor U47517 ( n46265,n46092,n46266 );
   nor U47518 ( n46249,n28273,n46194 );
   nand U47519 ( n46194,n46267,n46000 );
   nor U47520 ( n46000,n46268,n46269 );
   nor U47521 ( n46247,n46270,n46271 );
   nor U47522 ( n46271,n28323,n46197 );
   nand U47523 ( n46197,n46272,n46097 );
   nor U47524 ( n46097,n46273,n45437 );
   nor U47525 ( n46270,n46006,n46198 );
   nand U47526 ( n46198,n46274,n46007 );
   nor U47527 ( n46007,n45840,n46275 );
   nor U47528 ( n46277,n46278,n46279 );
   nand U47529 ( n46279,n46280,n46281 );
   nand U47530 ( n46281,n45887,n46282 );
   nand U47531 ( n46280,p1_instqueue_reg_11__7_,n46283 );
   nor U47532 ( n46278,n28192,n46284 );
   nor U47533 ( n46276,n46285,n46286 );
   nor U47534 ( n46286,n28316,n46287 );
   nor U47535 ( n46285,n45897,n46288 );
   nor U47536 ( n46290,n46291,n46292 );
   nand U47537 ( n46292,n46293,n46294 );
   nand U47538 ( n46294,n45904,n46282 );
   nand U47539 ( n46293,p1_instqueue_reg_11__6_,n46283 );
   nor U47540 ( n46291,n28198,n46284 );
   nor U47541 ( n46289,n46295,n46296 );
   nor U47542 ( n46296,n28317,n46287 );
   nor U47543 ( n46295,n45909,n46288 );
   nor U47544 ( n46298,n46299,n46300 );
   nand U47545 ( n46300,n46301,n46302 );
   nand U47546 ( n46302,n45916,n46282 );
   nand U47547 ( n46301,p1_instqueue_reg_11__5_,n46283 );
   nor U47548 ( n46299,n28204,n46284 );
   nor U47549 ( n46297,n46303,n46304 );
   nor U47550 ( n46304,n28318,n46287 );
   nor U47551 ( n46303,n45921,n46288 );
   nor U47552 ( n46306,n46307,n46308 );
   nand U47553 ( n46308,n46309,n46310 );
   nand U47554 ( n46310,n45928,n46282 );
   nand U47555 ( n46309,p1_instqueue_reg_11__4_,n46283 );
   nor U47556 ( n46307,n28211,n46284 );
   nor U47557 ( n46305,n46311,n46312 );
   nor U47558 ( n46312,n28319,n46287 );
   nor U47559 ( n46311,n45933,n46288 );
   nor U47560 ( n46314,n46315,n46316 );
   nand U47561 ( n46316,n46317,n46318 );
   nand U47562 ( n46318,n45940,n46282 );
   nand U47563 ( n46317,p1_instqueue_reg_11__3_,n46283 );
   nor U47564 ( n46315,n28219,n46284 );
   nor U47565 ( n46313,n46319,n46320 );
   nor U47566 ( n46320,n28320,n46287 );
   nor U47567 ( n46319,n45945,n46288 );
   nor U47568 ( n46322,n46323,n46324 );
   nand U47569 ( n46324,n46325,n46326 );
   nand U47570 ( n46326,n45952,n46282 );
   nand U47571 ( n46325,p1_instqueue_reg_11__2_,n46283 );
   nor U47572 ( n46323,n28231,n46284 );
   nor U47573 ( n46321,n46327,n46328 );
   nor U47574 ( n46328,n28321,n46287 );
   nor U47575 ( n46327,n45957,n46288 );
   nor U47576 ( n46330,n46331,n46332 );
   nand U47577 ( n46332,n46333,n46334 );
   nand U47578 ( n46334,n45964,n46282 );
   nand U47579 ( n46333,p1_instqueue_reg_11__1_,n46283 );
   nor U47580 ( n46331,n28249,n46284 );
   nor U47581 ( n46329,n46335,n46336 );
   nor U47582 ( n46336,n28322,n46287 );
   nor U47583 ( n46335,n45969,n46288 );
   nor U47584 ( n46338,n46339,n46340 );
   nand U47585 ( n46340,n46341,n46342 );
   nand U47586 ( n46342,n45976,n46282 );
   nand U47587 ( n46282,n46343,n46344 );
   nand U47588 ( n46344,p1_state2_reg_2_,n46345 );
   nand U47589 ( n46343,n46346,n45980 );
   nand U47590 ( n46341,p1_instqueue_reg_11__0_,n46283 );
   nand U47591 ( n46283,n46347,n46348 );
   nand U47592 ( n46348,p1_state2_reg_3_,n46288 );
   nor U47593 ( n46347,n46349,n46350 );
   nor U47594 ( n46350,n46351,n46352 );
   nand U47595 ( n46352,n46353,n45989 );
   nand U47596 ( n46353,n45990,n46354 );
   nand U47597 ( n46354,n46287,n46284 );
   and U47598 ( n46351,n46346,n45992 );
   nand U47599 ( n46346,n46288,n46355 );
   nand U47600 ( n46355,n46356,n45995 );
   nor U47601 ( n46349,n28375,n46345 );
   nand U47602 ( n46345,n46288,n46357 );
   nand U47603 ( n46357,n46358,n45998 );
   nor U47604 ( n46339,n28273,n46284 );
   nand U47605 ( n46284,n46359,n46001 );
   nor U47606 ( n46337,n46360,n46361 );
   nor U47607 ( n46361,n28323,n46287 );
   nand U47608 ( n46287,n46362,n45422 );
   nor U47609 ( n46360,n46006,n46288 );
   nand U47610 ( n46288,n46363,n46008 );
   nor U47611 ( n46365,n46366,n46367 );
   nand U47612 ( n46367,n46368,n46369 );
   nand U47613 ( n46369,n45887,n46370 );
   nand U47614 ( n46368,p1_instqueue_reg_10__7_,n46371 );
   nor U47615 ( n46366,n28192,n46372 );
   nor U47616 ( n46364,n46373,n46374 );
   nor U47617 ( n46374,n28316,n46375 );
   nor U47618 ( n46373,n45897,n46376 );
   nor U47619 ( n46378,n46379,n46380 );
   nand U47620 ( n46380,n46381,n46382 );
   nand U47621 ( n46382,n45904,n46370 );
   nand U47622 ( n46381,p1_instqueue_reg_10__6_,n46371 );
   nor U47623 ( n46379,n28198,n46372 );
   nor U47624 ( n46377,n46383,n46384 );
   nor U47625 ( n46384,n28317,n46375 );
   nor U47626 ( n46383,n45909,n46376 );
   nor U47627 ( n46386,n46387,n46388 );
   nand U47628 ( n46388,n46389,n46390 );
   nand U47629 ( n46390,n45916,n46370 );
   nand U47630 ( n46389,p1_instqueue_reg_10__5_,n46371 );
   nor U47631 ( n46387,n28204,n46372 );
   nor U47632 ( n46385,n46391,n46392 );
   nor U47633 ( n46392,n28318,n46375 );
   nor U47634 ( n46391,n45921,n46376 );
   nor U47635 ( n46394,n46395,n46396 );
   nand U47636 ( n46396,n46397,n46398 );
   nand U47637 ( n46398,n45928,n46370 );
   nand U47638 ( n46397,p1_instqueue_reg_10__4_,n46371 );
   nor U47639 ( n46395,n28211,n46372 );
   nor U47640 ( n46393,n46399,n46400 );
   nor U47641 ( n46400,n28319,n46375 );
   nor U47642 ( n46399,n45933,n46376 );
   nor U47643 ( n46402,n46403,n46404 );
   nand U47644 ( n46404,n46405,n46406 );
   nand U47645 ( n46406,n45940,n46370 );
   nand U47646 ( n46405,p1_instqueue_reg_10__3_,n46371 );
   nor U47647 ( n46403,n28219,n46372 );
   nor U47648 ( n46401,n46407,n46408 );
   nor U47649 ( n46408,n28320,n46375 );
   nor U47650 ( n46407,n45945,n46376 );
   nor U47651 ( n46410,n46411,n46412 );
   nand U47652 ( n46412,n46413,n46414 );
   nand U47653 ( n46414,n45952,n46370 );
   nand U47654 ( n46413,p1_instqueue_reg_10__2_,n46371 );
   nor U47655 ( n46411,n28231,n46372 );
   nor U47656 ( n46409,n46415,n46416 );
   nor U47657 ( n46416,n28321,n46375 );
   nor U47658 ( n46415,n45957,n46376 );
   nor U47659 ( n46418,n46419,n46420 );
   nand U47660 ( n46420,n46421,n46422 );
   nand U47661 ( n46422,n45964,n46370 );
   nand U47662 ( n46421,p1_instqueue_reg_10__1_,n46371 );
   nor U47663 ( n46419,n28249,n46372 );
   nor U47664 ( n46417,n46423,n46424 );
   nor U47665 ( n46424,n28322,n46375 );
   nor U47666 ( n46423,n45969,n46376 );
   nor U47667 ( n46426,n46427,n46428 );
   nand U47668 ( n46428,n46429,n46430 );
   nand U47669 ( n46430,n45976,n46370 );
   nand U47670 ( n46370,n46431,n46432 );
   nand U47671 ( n46432,n46433,n45998 );
   nand U47672 ( n46431,n46434,n45980 );
   not U47673 ( n46434,n46435 );
   nand U47674 ( n46429,p1_instqueue_reg_10__0_,n46371 );
   nand U47675 ( n46371,n46436,n46437 );
   nand U47676 ( n46437,p1_state2_reg_3_,n46376 );
   nor U47677 ( n46436,n46438,n46439 );
   nor U47678 ( n46439,n46440,n46441 );
   nand U47679 ( n46441,n46442,n45989 );
   nand U47680 ( n46442,n45990,n46443 );
   nand U47681 ( n46443,n46375,n46372 );
   nor U47682 ( n46440,n46435,n28281 );
   nand U47683 ( n46435,n46356,n46090 );
   nor U47684 ( n46438,n46444,n28374 );
   nor U47685 ( n46444,n46093,n46445 );
   not U47686 ( n46093,n45998 );
   nor U47687 ( n45998,n46446,n46447 );
   nor U47688 ( n46427,n28273,n46372 );
   nand U47689 ( n46372,n46359,n46094 );
   nor U47690 ( n46425,n46448,n46449 );
   nor U47691 ( n46449,n28323,n46375 );
   nand U47692 ( n46375,n46362,n45407 );
   nor U47693 ( n46448,n46006,n46376 );
   nand U47694 ( n46376,n46363,n46098 );
   nor U47695 ( n46451,n46452,n46453 );
   nand U47696 ( n46453,n46454,n46455 );
   nand U47697 ( n46455,n45887,n46456 );
   nand U47698 ( n46454,p1_instqueue_reg_9__7_,n46457 );
   nor U47699 ( n46452,n28192,n46458 );
   nor U47700 ( n46450,n46459,n46460 );
   nor U47701 ( n46460,n28316,n46461 );
   nor U47702 ( n46459,n28189,n46462 );
   nor U47703 ( n46464,n46465,n46466 );
   nand U47704 ( n46466,n46467,n46468 );
   nand U47705 ( n46468,n45904,n46456 );
   nand U47706 ( n46467,p1_instqueue_reg_9__6_,n46457 );
   nor U47707 ( n46465,n28198,n46458 );
   nor U47708 ( n46463,n46469,n46470 );
   nor U47709 ( n46470,n28317,n46461 );
   nor U47710 ( n46469,n28194,n46462 );
   nor U47711 ( n46472,n46473,n46474 );
   nand U47712 ( n46474,n46475,n46476 );
   nand U47713 ( n46476,n45916,n46456 );
   nand U47714 ( n46475,p1_instqueue_reg_9__5_,n46457 );
   nor U47715 ( n46473,n28204,n46458 );
   nor U47716 ( n46471,n46477,n46478 );
   nor U47717 ( n46478,n28318,n46461 );
   nor U47718 ( n46477,n28200,n46462 );
   nor U47719 ( n46480,n46481,n46482 );
   nand U47720 ( n46482,n46483,n46484 );
   nand U47721 ( n46484,n45928,n46456 );
   nand U47722 ( n46483,p1_instqueue_reg_9__4_,n46457 );
   nor U47723 ( n46481,n28211,n46458 );
   nor U47724 ( n46479,n46485,n46486 );
   nor U47725 ( n46486,n28319,n46461 );
   nor U47726 ( n46485,n28207,n46462 );
   nor U47727 ( n46488,n46489,n46490 );
   nand U47728 ( n46490,n46491,n46492 );
   nand U47729 ( n46492,n45940,n46456 );
   nand U47730 ( n46491,p1_instqueue_reg_9__3_,n46457 );
   nor U47731 ( n46489,n28219,n46458 );
   nor U47732 ( n46487,n46493,n46494 );
   nor U47733 ( n46494,n28320,n46461 );
   nor U47734 ( n46493,n28215,n46462 );
   nor U47735 ( n46496,n46497,n46498 );
   nand U47736 ( n46498,n46499,n46500 );
   nand U47737 ( n46500,n45952,n46456 );
   nand U47738 ( n46499,p1_instqueue_reg_9__2_,n46457 );
   nor U47739 ( n46497,n28231,n46458 );
   nor U47740 ( n46495,n46501,n46502 );
   nor U47741 ( n46502,n28321,n46461 );
   nor U47742 ( n46501,n28227,n46462 );
   nor U47743 ( n46504,n46505,n46506 );
   nand U47744 ( n46506,n46507,n46508 );
   nand U47745 ( n46508,n45964,n46456 );
   nand U47746 ( n46507,p1_instqueue_reg_9__1_,n46457 );
   nor U47747 ( n46505,n28249,n46458 );
   nor U47748 ( n46503,n46509,n46510 );
   nor U47749 ( n46510,n28322,n46461 );
   nor U47750 ( n46509,n28245,n46462 );
   nor U47751 ( n46512,n46513,n46514 );
   nand U47752 ( n46514,n46515,n46516 );
   nand U47753 ( n46516,n45976,n46456 );
   nand U47754 ( n46456,n46517,n46518 );
   nand U47755 ( n46518,p1_state2_reg_2_,n46519 );
   nand U47756 ( n46517,n46520,n45980 );
   nand U47757 ( n46515,p1_instqueue_reg_9__0_,n46457 );
   nand U47758 ( n46457,n46521,n46522 );
   nand U47759 ( n46522,p1_state2_reg_3_,n46462 );
   nor U47760 ( n46521,n46523,n46524 );
   nor U47761 ( n46524,n46525,n46526 );
   nand U47762 ( n46526,n46527,n45989 );
   nand U47763 ( n46527,n45990,n46528 );
   nand U47764 ( n46528,n46461,n46458 );
   and U47765 ( n46525,n46520,n45992 );
   nand U47766 ( n46520,n46462,n46529 );
   nand U47767 ( n46529,n46356,n46179 );
   nor U47768 ( n46523,n28375,n46519 );
   nand U47769 ( n46519,n46462,n46530 );
   nand U47770 ( n46530,n46358,n46181 );
   nor U47771 ( n46513,n28273,n46458 );
   nand U47772 ( n46458,n46359,n46182 );
   nor U47773 ( n46511,n46531,n46532 );
   nor U47774 ( n46532,n28323,n46461 );
   nand U47775 ( n46461,n46362,n45408 );
   nor U47776 ( n46531,n28325,n46462 );
   nand U47777 ( n46462,n46363,n46185 );
   nor U47778 ( n46534,n46535,n46536 );
   nand U47779 ( n46536,n46537,n46538 );
   nand U47780 ( n46538,n45887,n46539 );
   nand U47781 ( n46537,p1_instqueue_reg_8__7_,n46540 );
   nor U47782 ( n46535,n45890,n46541 );
   nor U47783 ( n46533,n46542,n46543 );
   nor U47784 ( n46543,n45894,n46544 );
   nor U47785 ( n46542,n28189,n46545 );
   nor U47786 ( n46547,n46548,n46549 );
   nand U47787 ( n46549,n46550,n46551 );
   nand U47788 ( n46551,n45904,n46539 );
   nand U47789 ( n46550,p1_instqueue_reg_8__6_,n46540 );
   nor U47790 ( n46548,n45905,n46541 );
   nor U47791 ( n46546,n46552,n46553 );
   nor U47792 ( n46553,n45908,n46544 );
   nor U47793 ( n46552,n28194,n46545 );
   nor U47794 ( n46555,n46556,n46557 );
   nand U47795 ( n46557,n46558,n46559 );
   nand U47796 ( n46559,n45916,n46539 );
   nand U47797 ( n46558,p1_instqueue_reg_8__5_,n46540 );
   nor U47798 ( n46556,n45917,n46541 );
   nor U47799 ( n46554,n46560,n46561 );
   nor U47800 ( n46561,n45920,n46544 );
   nor U47801 ( n46560,n28200,n46545 );
   nor U47802 ( n46563,n46564,n46565 );
   nand U47803 ( n46565,n46566,n46567 );
   nand U47804 ( n46567,n45928,n46539 );
   nand U47805 ( n46566,p1_instqueue_reg_8__4_,n46540 );
   nor U47806 ( n46564,n45929,n46541 );
   nor U47807 ( n46562,n46568,n46569 );
   nor U47808 ( n46569,n45932,n46544 );
   nor U47809 ( n46568,n28207,n46545 );
   nor U47810 ( n46571,n46572,n46573 );
   nand U47811 ( n46573,n46574,n46575 );
   nand U47812 ( n46575,n45940,n46539 );
   nand U47813 ( n46574,p1_instqueue_reg_8__3_,n46540 );
   nor U47814 ( n46572,n45941,n46541 );
   nor U47815 ( n46570,n46576,n46577 );
   nor U47816 ( n46577,n45944,n46544 );
   nor U47817 ( n46576,n28215,n46545 );
   nor U47818 ( n46579,n46580,n46581 );
   nand U47819 ( n46581,n46582,n46583 );
   nand U47820 ( n46583,n45952,n46539 );
   nand U47821 ( n46582,p1_instqueue_reg_8__2_,n46540 );
   nor U47822 ( n46580,n45953,n46541 );
   nor U47823 ( n46578,n46584,n46585 );
   nor U47824 ( n46585,n45956,n46544 );
   nor U47825 ( n46584,n28227,n46545 );
   nor U47826 ( n46587,n46588,n46589 );
   nand U47827 ( n46589,n46590,n46591 );
   nand U47828 ( n46591,n45964,n46539 );
   nand U47829 ( n46590,p1_instqueue_reg_8__1_,n46540 );
   nor U47830 ( n46588,n45965,n46541 );
   nor U47831 ( n46586,n46592,n46593 );
   nor U47832 ( n46593,n45968,n46544 );
   nor U47833 ( n46592,n28245,n46545 );
   nor U47834 ( n46595,n46596,n46597 );
   nand U47835 ( n46597,n46598,n46599 );
   nand U47836 ( n46599,n45976,n46539 );
   nand U47837 ( n46539,n46600,n46601 );
   nand U47838 ( n46601,n46433,n46181 );
   nand U47839 ( n46600,n46602,n45980 );
   not U47840 ( n46602,n46603 );
   nand U47841 ( n46598,p1_instqueue_reg_8__0_,n46540 );
   nand U47842 ( n46540,n46604,n46605 );
   nand U47843 ( n46605,p1_state2_reg_3_,n46545 );
   nor U47844 ( n46604,n46606,n46607 );
   nor U47845 ( n46607,n46608,n46609 );
   nand U47846 ( n46609,n46610,n45989 );
   nand U47847 ( n46610,n45990,n46611 );
   nand U47848 ( n46611,n46544,n46541 );
   nor U47849 ( n46608,n46603,n46089 );
   nand U47850 ( n46603,n46356,n45404 );
   nor U47851 ( n46356,n46612,n45431 );
   nor U47852 ( n46606,n46613,n45355 );
   nor U47853 ( n46613,n46266,n46445 );
   not U47854 ( n46266,n46181 );
   nor U47855 ( n46181,n46614,n46446 );
   nor U47856 ( n46596,n45999,n46541 );
   nand U47857 ( n46541,n46359,n46267 );
   nor U47858 ( n46594,n46615,n46616 );
   nor U47859 ( n46616,n46004,n46544 );
   nand U47860 ( n46544,n46362,n46272 );
   nor U47861 ( n46362,n45421,n45437 );
   not U47862 ( n45437,n46005 );
   nor U47863 ( n46615,n28325,n46545 );
   nand U47864 ( n46545,n46363,n46274 );
   nor U47865 ( n46618,n46619,n46620 );
   nand U47866 ( n46620,n46621,n46622 );
   nand U47867 ( n46622,n45887,n46623 );
   nand U47868 ( n46621,p1_instqueue_reg_7__7_,n46624 );
   nor U47869 ( n46619,n45894,n46625 );
   nor U47870 ( n46617,n46626,n46627 );
   nor U47871 ( n46627,n45890,n46628 );
   nor U47872 ( n46626,n45897,n46629 );
   nor U47873 ( n46631,n46632,n46633 );
   nand U47874 ( n46633,n46634,n46635 );
   nand U47875 ( n46635,n45904,n46623 );
   nand U47876 ( n46634,p1_instqueue_reg_7__6_,n46624 );
   nor U47877 ( n46632,n45908,n46625 );
   nor U47878 ( n46630,n46636,n46637 );
   nor U47879 ( n46637,n45905,n46628 );
   nor U47880 ( n46636,n45909,n46629 );
   nor U47881 ( n46639,n46640,n46641 );
   nand U47882 ( n46641,n46642,n46643 );
   nand U47883 ( n46643,n45916,n46623 );
   nand U47884 ( n46642,p1_instqueue_reg_7__5_,n46624 );
   nor U47885 ( n46640,n45920,n46625 );
   nor U47886 ( n46638,n46644,n46645 );
   nor U47887 ( n46645,n45917,n46628 );
   nor U47888 ( n46644,n45921,n46629 );
   nor U47889 ( n46647,n46648,n46649 );
   nand U47890 ( n46649,n46650,n46651 );
   nand U47891 ( n46651,n45928,n46623 );
   nand U47892 ( n46650,p1_instqueue_reg_7__4_,n46624 );
   nor U47893 ( n46648,n45932,n46625 );
   nor U47894 ( n46646,n46652,n46653 );
   nor U47895 ( n46653,n45929,n46628 );
   nor U47896 ( n46652,n45933,n46629 );
   nor U47897 ( n46655,n46656,n46657 );
   nand U47898 ( n46657,n46658,n46659 );
   nand U47899 ( n46659,n45940,n46623 );
   nand U47900 ( n46658,p1_instqueue_reg_7__3_,n46624 );
   nor U47901 ( n46656,n45944,n46625 );
   nor U47902 ( n46654,n46660,n46661 );
   nor U47903 ( n46661,n45941,n46628 );
   nor U47904 ( n46660,n45945,n46629 );
   nor U47905 ( n46663,n46664,n46665 );
   nand U47906 ( n46665,n46666,n46667 );
   nand U47907 ( n46667,n45952,n46623 );
   nand U47908 ( n46666,p1_instqueue_reg_7__2_,n46624 );
   nor U47909 ( n46664,n45956,n46625 );
   nor U47910 ( n46662,n46668,n46669 );
   nor U47911 ( n46669,n45953,n46628 );
   nor U47912 ( n46668,n45957,n46629 );
   nor U47913 ( n46671,n46672,n46673 );
   nand U47914 ( n46673,n46674,n46675 );
   nand U47915 ( n46675,n45964,n46623 );
   nand U47916 ( n46674,p1_instqueue_reg_7__1_,n46624 );
   nor U47917 ( n46672,n45968,n46625 );
   nor U47918 ( n46670,n46676,n46677 );
   nor U47919 ( n46677,n45965,n46628 );
   nor U47920 ( n46676,n45969,n46629 );
   nor U47921 ( n46679,n46680,n46681 );
   nand U47922 ( n46681,n46682,n46683 );
   nand U47923 ( n46683,n45976,n46623 );
   nand U47924 ( n46623,n46684,n46685 );
   nand U47925 ( n46685,p1_state2_reg_2_,n46686 );
   nand U47926 ( n46684,n46687,n45980 );
   nand U47927 ( n46682,p1_instqueue_reg_7__0_,n46624 );
   nand U47928 ( n46624,n46688,n46689 );
   nor U47929 ( n46689,n46690,n46691 );
   nor U47930 ( n46691,n45355,n46686 );
   nand U47931 ( n46686,n46629,n46692 );
   nand U47932 ( n46692,n46693,n45997 );
   nor U47933 ( n46690,n46687,n46694 );
   nand U47934 ( n46694,n46695,n46696 );
   nand U47935 ( n46695,n46697,n46698 );
   nand U47936 ( n46698,n46628,n46625 );
   nand U47937 ( n46687,n46629,n46699 );
   nand U47938 ( n46699,n46700,n45995 );
   nor U47939 ( n46688,n46701,n46089 );
   nor U47940 ( n46701,n46702,n45501 );
   nor U47941 ( n46680,n46004,n46625 );
   not U47942 ( n46625,n45435 );
   nor U47943 ( n45435,n45420,n46005 );
   nand U47944 ( n45420,n45422,n45421 );
   nor U47945 ( n46678,n46703,n46704 );
   nor U47946 ( n46704,n45999,n46628 );
   nor U47947 ( n46703,n46006,n46629 );
   nor U47948 ( n46706,n46707,n46708 );
   nand U47949 ( n46708,n46709,n46710 );
   nand U47950 ( n46710,n45887,n46711 );
   nand U47951 ( n46709,p1_instqueue_reg_6__7_,n46712 );
   nor U47952 ( n46707,n45890,n46713 );
   nor U47953 ( n46705,n46714,n46715 );
   nor U47954 ( n46715,n45894,n46716 );
   nor U47955 ( n46714,n28189,n46717 );
   nor U47956 ( n46719,n46720,n46721 );
   nand U47957 ( n46721,n46722,n46723 );
   nand U47958 ( n46723,n45904,n46711 );
   nand U47959 ( n46722,p1_instqueue_reg_6__6_,n46712 );
   nor U47960 ( n46720,n45905,n46713 );
   nor U47961 ( n46718,n46724,n46725 );
   nor U47962 ( n46725,n45908,n46716 );
   nor U47963 ( n46724,n28194,n46717 );
   nor U47964 ( n46727,n46728,n46729 );
   nand U47965 ( n46729,n46730,n46731 );
   nand U47966 ( n46731,n45916,n46711 );
   nand U47967 ( n46730,p1_instqueue_reg_6__5_,n46712 );
   nor U47968 ( n46728,n45917,n46713 );
   nor U47969 ( n46726,n46732,n46733 );
   nor U47970 ( n46733,n45920,n46716 );
   nor U47971 ( n46732,n28200,n46717 );
   nor U47972 ( n46735,n46736,n46737 );
   nand U47973 ( n46737,n46738,n46739 );
   nand U47974 ( n46739,n45928,n46711 );
   nand U47975 ( n46738,p1_instqueue_reg_6__4_,n46712 );
   nor U47976 ( n46736,n45929,n46713 );
   nor U47977 ( n46734,n46740,n46741 );
   nor U47978 ( n46741,n45932,n46716 );
   nor U47979 ( n46740,n28207,n46717 );
   nor U47980 ( n46743,n46744,n46745 );
   nand U47981 ( n46745,n46746,n46747 );
   nand U47982 ( n46747,n45940,n46711 );
   nand U47983 ( n46746,p1_instqueue_reg_6__3_,n46712 );
   nor U47984 ( n46744,n45941,n46713 );
   nor U47985 ( n46742,n46748,n46749 );
   nor U47986 ( n46749,n45944,n46716 );
   nor U47987 ( n46748,n28215,n46717 );
   nor U47988 ( n46751,n46752,n46753 );
   nand U47989 ( n46753,n46754,n46755 );
   nand U47990 ( n46755,n45952,n46711 );
   nand U47991 ( n46754,p1_instqueue_reg_6__2_,n46712 );
   nor U47992 ( n46752,n45953,n46713 );
   nor U47993 ( n46750,n46756,n46757 );
   nor U47994 ( n46757,n45956,n46716 );
   nor U47995 ( n46756,n28227,n46717 );
   nor U47996 ( n46759,n46760,n46761 );
   nand U47997 ( n46761,n46762,n46763 );
   nand U47998 ( n46763,n45964,n46711 );
   nand U47999 ( n46762,p1_instqueue_reg_6__1_,n46712 );
   nor U48000 ( n46760,n45965,n46713 );
   nor U48001 ( n46758,n46764,n46765 );
   nor U48002 ( n46765,n45968,n46716 );
   nor U48003 ( n46764,n28245,n46717 );
   nor U48004 ( n46767,n46768,n46769 );
   nand U48005 ( n46769,n46770,n46771 );
   nand U48006 ( n46771,n45976,n46711 );
   nand U48007 ( n46711,n46772,n46773 );
   nand U48008 ( n46773,n46693,n46078 );
   nand U48009 ( n46772,n46774,n45980 );
   not U48010 ( n46774,n46775 );
   nand U48011 ( n46770,p1_instqueue_reg_6__0_,n46712 );
   nand U48012 ( n46712,n46776,n46777 );
   nand U48013 ( n46777,p1_state2_reg_3_,n46717 );
   nor U48014 ( n46776,n46778,n46779 );
   nor U48015 ( n46779,n46780,n46781 );
   nand U48016 ( n46781,n46782,n45989 );
   nand U48017 ( n46782,n45990,n46783 );
   nand U48018 ( n46783,n46716,n46713 );
   nor U48019 ( n46780,n46775,n46089 );
   nand U48020 ( n46775,n46700,n46090 );
   nor U48021 ( n46778,n46784,n28375 );
   nor U48022 ( n46784,n46092,n46785 );
   nor U48023 ( n46768,n45999,n46713 );
   nand U48024 ( n46713,n46094,n46786 );
   nor U48025 ( n46766,n46787,n46788 );
   nor U48026 ( n46788,n46004,n46716 );
   nand U48027 ( n46716,n46789,n45407 );
   nor U48028 ( n46787,n28325,n46717 );
   nand U48029 ( n46717,n46098,n46790 );
   nor U48030 ( n46792,n46793,n46794 );
   nand U48031 ( n46794,n46795,n46796 );
   nand U48032 ( n46796,n45887,n46797 );
   nand U48033 ( n46795,p1_instqueue_reg_5__7_,n46798 );
   nor U48034 ( n46793,n45890,n46799 );
   nor U48035 ( n46791,n46800,n46801 );
   nor U48036 ( n46801,n45894,n46802 );
   nor U48037 ( n46800,n45897,n46803 );
   nor U48038 ( n46805,n46806,n46807 );
   nand U48039 ( n46807,n46808,n46809 );
   nand U48040 ( n46809,n45904,n46797 );
   nand U48041 ( n46808,p1_instqueue_reg_5__6_,n46798 );
   nor U48042 ( n46806,n45905,n46799 );
   nor U48043 ( n46804,n46810,n46811 );
   nor U48044 ( n46811,n45908,n46802 );
   nor U48045 ( n46810,n45909,n46803 );
   nor U48046 ( n46813,n46814,n46815 );
   nand U48047 ( n46815,n46816,n46817 );
   nand U48048 ( n46817,n45916,n46797 );
   nand U48049 ( n46816,p1_instqueue_reg_5__5_,n46798 );
   nor U48050 ( n46814,n45917,n46799 );
   nor U48051 ( n46812,n46818,n46819 );
   nor U48052 ( n46819,n45920,n46802 );
   nor U48053 ( n46818,n45921,n46803 );
   nor U48054 ( n46821,n46822,n46823 );
   nand U48055 ( n46823,n46824,n46825 );
   nand U48056 ( n46825,n45928,n46797 );
   nand U48057 ( n46824,p1_instqueue_reg_5__4_,n46798 );
   nor U48058 ( n46822,n45929,n46799 );
   nor U48059 ( n46820,n46826,n46827 );
   nor U48060 ( n46827,n45932,n46802 );
   nor U48061 ( n46826,n45933,n46803 );
   nor U48062 ( n46829,n46830,n46831 );
   nand U48063 ( n46831,n46832,n46833 );
   nand U48064 ( n46833,n45940,n46797 );
   nand U48065 ( n46832,p1_instqueue_reg_5__3_,n46798 );
   nor U48066 ( n46830,n45941,n46799 );
   nor U48067 ( n46828,n46834,n46835 );
   nor U48068 ( n46835,n45944,n46802 );
   nor U48069 ( n46834,n45945,n46803 );
   nor U48070 ( n46837,n46838,n46839 );
   nand U48071 ( n46839,n46840,n46841 );
   nand U48072 ( n46841,n45952,n46797 );
   nand U48073 ( n46840,p1_instqueue_reg_5__2_,n46798 );
   nor U48074 ( n46838,n45953,n46799 );
   nor U48075 ( n46836,n46842,n46843 );
   nor U48076 ( n46843,n45956,n46802 );
   nor U48077 ( n46842,n45957,n46803 );
   nor U48078 ( n46845,n46846,n46847 );
   nand U48079 ( n46847,n46848,n46849 );
   nand U48080 ( n46849,n45964,n46797 );
   nand U48081 ( n46848,p1_instqueue_reg_5__1_,n46798 );
   nor U48082 ( n46846,n45965,n46799 );
   nor U48083 ( n46844,n46850,n46851 );
   nor U48084 ( n46851,n45968,n46802 );
   nor U48085 ( n46850,n45969,n46803 );
   nor U48086 ( n46853,n46854,n46855 );
   nand U48087 ( n46855,n46856,n46857 );
   nand U48088 ( n46857,n45976,n46797 );
   nand U48089 ( n46797,n46858,n46859 );
   nand U48090 ( n46859,p1_state2_reg_2_,n46860 );
   nand U48091 ( n46858,n46861,n45980 );
   nand U48092 ( n46856,p1_instqueue_reg_5__0_,n46798 );
   nand U48093 ( n46798,n46862,n46863 );
   nand U48094 ( n46863,p1_state2_reg_3_,n46803 );
   nor U48095 ( n46862,n46864,n46865 );
   nor U48096 ( n46865,n46866,n46867 );
   nand U48097 ( n46867,n46868,n45989 );
   nand U48098 ( n46868,n45990,n46869 );
   nand U48099 ( n46869,n46802,n46799 );
   and U48100 ( n46866,n46861,n45992 );
   nand U48101 ( n46861,n46803,n46870 );
   nand U48102 ( n46870,n46700,n46179 );
   nor U48103 ( n46864,n28375,n46860 );
   nand U48104 ( n46860,n46803,n46871 );
   nand U48105 ( n46871,n46872,n45997 );
   nor U48106 ( n45997,n46092,p1_instqueuewr_addr_reg_0_ );
   nor U48107 ( n46854,n45999,n46799 );
   nand U48108 ( n46799,n46182,n46786 );
   nor U48109 ( n46852,n46873,n46874 );
   nor U48110 ( n46874,n46004,n46802 );
   nand U48111 ( n46802,n46789,n45408 );
   nor U48112 ( n46873,n46006,n46803 );
   nand U48113 ( n46803,n46185,n46790 );
   nor U48114 ( n46876,n46877,n46878 );
   nand U48115 ( n46878,n46879,n46880 );
   nand U48116 ( n46880,n45887,n46881 );
   nand U48117 ( n46879,p1_instqueue_reg_4__7_,n46882 );
   nor U48118 ( n46877,n45890,n46883 );
   nor U48119 ( n46875,n46884,n46885 );
   nor U48120 ( n46885,n45894,n46886 );
   nor U48121 ( n46884,n45897,n46887 );
   nor U48122 ( n46889,n46890,n46891 );
   nand U48123 ( n46891,n46892,n46893 );
   nand U48124 ( n46893,n45904,n46881 );
   nand U48125 ( n46892,p1_instqueue_reg_4__6_,n46882 );
   nor U48126 ( n46890,n45905,n46883 );
   nor U48127 ( n46888,n46894,n46895 );
   nor U48128 ( n46895,n45908,n46886 );
   nor U48129 ( n46894,n45909,n46887 );
   nor U48130 ( n46897,n46898,n46899 );
   nand U48131 ( n46899,n46900,n46901 );
   nand U48132 ( n46901,n45916,n46881 );
   nand U48133 ( n46900,p1_instqueue_reg_4__5_,n46882 );
   nor U48134 ( n46898,n45917,n46883 );
   nor U48135 ( n46896,n46902,n46903 );
   nor U48136 ( n46903,n45920,n46886 );
   nor U48137 ( n46902,n45921,n46887 );
   nor U48138 ( n46905,n46906,n46907 );
   nand U48139 ( n46907,n46908,n46909 );
   nand U48140 ( n46909,n45928,n46881 );
   nand U48141 ( n46908,p1_instqueue_reg_4__4_,n46882 );
   nor U48142 ( n46906,n45929,n46883 );
   nor U48143 ( n46904,n46910,n46911 );
   nor U48144 ( n46911,n45932,n46886 );
   nor U48145 ( n46910,n45933,n46887 );
   nor U48146 ( n46913,n46914,n46915 );
   nand U48147 ( n46915,n46916,n46917 );
   nand U48148 ( n46917,n45940,n46881 );
   nand U48149 ( n46916,p1_instqueue_reg_4__3_,n46882 );
   nor U48150 ( n46914,n45941,n46883 );
   nor U48151 ( n46912,n46918,n46919 );
   nor U48152 ( n46919,n45944,n46886 );
   nor U48153 ( n46918,n45945,n46887 );
   nor U48154 ( n46921,n46922,n46923 );
   nand U48155 ( n46923,n46924,n46925 );
   nand U48156 ( n46925,n45952,n46881 );
   nand U48157 ( n46924,p1_instqueue_reg_4__2_,n46882 );
   nor U48158 ( n46922,n45953,n46883 );
   nor U48159 ( n46920,n46926,n46927 );
   nor U48160 ( n46927,n45956,n46886 );
   nor U48161 ( n46926,n45957,n46887 );
   nor U48162 ( n46929,n46930,n46931 );
   nand U48163 ( n46931,n46932,n46933 );
   nand U48164 ( n46933,n45964,n46881 );
   nand U48165 ( n46932,p1_instqueue_reg_4__1_,n46882 );
   nor U48166 ( n46930,n45965,n46883 );
   nor U48167 ( n46928,n46934,n46935 );
   nor U48168 ( n46935,n45968,n46886 );
   nor U48169 ( n46934,n45969,n46887 );
   nor U48170 ( n46937,n46938,n46939 );
   nand U48171 ( n46939,n46940,n46941 );
   nand U48172 ( n46941,n45976,n46881 );
   nand U48173 ( n46881,n46942,n46943 );
   nand U48174 ( n46943,n46872,n46078 );
   nor U48175 ( n46078,n45355,n46092 );
   nand U48176 ( n46942,n46944,n45980 );
   not U48177 ( n46944,n46945 );
   nand U48178 ( n46940,p1_instqueue_reg_4__0_,n46882 );
   nand U48179 ( n46882,n46946,n46947 );
   nand U48180 ( n46947,p1_state2_reg_3_,n46887 );
   nor U48181 ( n46946,n46948,n46949 );
   nor U48182 ( n46949,n46950,n46951 );
   nand U48183 ( n46951,n46952,n45989 );
   nand U48184 ( n46952,n45990,n46953 );
   nand U48185 ( n46953,n46886,n46883 );
   nor U48186 ( n46950,n46945,n28281 );
   nand U48187 ( n46945,n46700,n45404 );
   nor U48188 ( n46700,n45417,n46954 );
   nor U48189 ( n46948,n46955,n28375 );
   nor U48190 ( n46955,n46092,n46956 );
   not U48191 ( n46092,n46445 );
   nor U48192 ( n46938,n45999,n46883 );
   nand U48193 ( n46883,n46267,n46786 );
   nor U48194 ( n46936,n46957,n46958 );
   nor U48195 ( n46958,n46004,n46886 );
   nand U48196 ( n46886,n46789,n46272 );
   nor U48197 ( n46789,n46005,n46273 );
   nor U48198 ( n46957,n46006,n46887 );
   nand U48199 ( n46887,n46274,n46790 );
   nor U48200 ( n46960,n46961,n46962 );
   nand U48201 ( n46962,n46963,n46964 );
   nand U48202 ( n46964,n45887,n46965 );
   nand U48203 ( n46963,p1_instqueue_reg_3__7_,n46966 );
   nor U48204 ( n46961,n45890,n46967 );
   nor U48205 ( n46959,n46968,n46969 );
   nor U48206 ( n46969,n45894,n46970 );
   nor U48207 ( n46968,n45897,n46971 );
   nor U48208 ( n46973,n46974,n46975 );
   nand U48209 ( n46975,n46976,n46977 );
   nand U48210 ( n46977,n45904,n46965 );
   nand U48211 ( n46976,p1_instqueue_reg_3__6_,n46966 );
   nor U48212 ( n46974,n45905,n46967 );
   nor U48213 ( n46972,n46978,n46979 );
   nor U48214 ( n46979,n45908,n46970 );
   nor U48215 ( n46978,n45909,n46971 );
   nor U48216 ( n46981,n46982,n46983 );
   nand U48217 ( n46983,n46984,n46985 );
   nand U48218 ( n46985,n45916,n46965 );
   nand U48219 ( n46984,p1_instqueue_reg_3__5_,n46966 );
   nor U48220 ( n46982,n45917,n46967 );
   nor U48221 ( n46980,n46986,n46987 );
   nor U48222 ( n46987,n45920,n46970 );
   nor U48223 ( n46986,n45921,n46971 );
   nor U48224 ( n46989,n46990,n46991 );
   nand U48225 ( n46991,n46992,n46993 );
   nand U48226 ( n46993,n45928,n46965 );
   nand U48227 ( n46992,p1_instqueue_reg_3__4_,n46966 );
   nor U48228 ( n46990,n45929,n46967 );
   nor U48229 ( n46988,n46994,n46995 );
   nor U48230 ( n46995,n45932,n46970 );
   nor U48231 ( n46994,n45933,n46971 );
   nor U48232 ( n46997,n46998,n46999 );
   nand U48233 ( n46999,n47000,n47001 );
   nand U48234 ( n47001,n45940,n46965 );
   nand U48235 ( n47000,p1_instqueue_reg_3__3_,n46966 );
   nor U48236 ( n46998,n45941,n46967 );
   nor U48237 ( n46996,n47002,n47003 );
   nor U48238 ( n47003,n45944,n46970 );
   nor U48239 ( n47002,n45945,n46971 );
   nor U48240 ( n47005,n47006,n47007 );
   nand U48241 ( n47007,n47008,n47009 );
   nand U48242 ( n47009,n45952,n46965 );
   nand U48243 ( n47008,p1_instqueue_reg_3__2_,n46966 );
   nor U48244 ( n47006,n45953,n46967 );
   nor U48245 ( n47004,n47010,n47011 );
   nor U48246 ( n47011,n45956,n46970 );
   nor U48247 ( n47010,n45957,n46971 );
   nor U48248 ( n47013,n47014,n47015 );
   nand U48249 ( n47015,n47016,n47017 );
   nand U48250 ( n47017,n45964,n46965 );
   nand U48251 ( n47016,p1_instqueue_reg_3__1_,n46966 );
   nor U48252 ( n47014,n45965,n46967 );
   nor U48253 ( n47012,n47018,n47019 );
   nor U48254 ( n47019,n45968,n46970 );
   nor U48255 ( n47018,n45969,n46971 );
   nor U48256 ( n47021,n47022,n47023 );
   nand U48257 ( n47023,n47024,n47025 );
   nand U48258 ( n47025,n45976,n46965 );
   nand U48259 ( n46965,n47026,n47027 );
   nand U48260 ( n47027,p1_state2_reg_2_,n47028 );
   nand U48261 ( n47026,n47029,n45980 );
   nand U48262 ( n47024,p1_instqueue_reg_3__0_,n46966 );
   nand U48263 ( n46966,n47030,n47031 );
   nand U48264 ( n47031,p1_state2_reg_3_,n46971 );
   nor U48265 ( n47030,n47032,n47033 );
   nor U48266 ( n47033,n47034,n47035 );
   nand U48267 ( n47035,n47036,n45989 );
   nand U48268 ( n47036,n45990,n47037 );
   nand U48269 ( n47037,n46970,n46967 );
   and U48270 ( n47034,n47029,n45992 );
   nand U48271 ( n47029,n46971,n47038 );
   nand U48272 ( n47038,n47039,n45995 );
   nor U48273 ( n45995,n45394,n45404 );
   nor U48274 ( n47032,n28374,n47028 );
   nand U48275 ( n47028,n46971,n47040 );
   nand U48276 ( n47040,n46693,n46358 );
   nor U48277 ( n47022,n45999,n46967 );
   nand U48278 ( n46967,n47041,n46001 );
   nor U48279 ( n47020,n47042,n47043 );
   nor U48280 ( n47043,n46004,n46970 );
   nand U48281 ( n46970,n47044,n45422 );
   nor U48282 ( n45422,n45389,n47045 );
   nor U48283 ( n47042,n46006,n46971 );
   nand U48284 ( n46971,n47046,n46008 );
   nor U48285 ( n47048,n47049,n47050 );
   nand U48286 ( n47050,n47051,n47052 );
   nand U48287 ( n47052,n45887,n47053 );
   nand U48288 ( n47051,p1_instqueue_reg_2__7_,n47054 );
   nor U48289 ( n47049,n45890,n47055 );
   nor U48290 ( n47047,n47056,n47057 );
   nor U48291 ( n47057,n45894,n47058 );
   nor U48292 ( n47056,n45897,n47059 );
   nor U48293 ( n47061,n47062,n47063 );
   nand U48294 ( n47063,n47064,n47065 );
   nand U48295 ( n47065,n45904,n47053 );
   nand U48296 ( n47064,p1_instqueue_reg_2__6_,n47054 );
   nor U48297 ( n47062,n45905,n47055 );
   nor U48298 ( n47060,n47066,n47067 );
   nor U48299 ( n47067,n45908,n47058 );
   nor U48300 ( n47066,n45909,n47059 );
   nor U48301 ( n47069,n47070,n47071 );
   nand U48302 ( n47071,n47072,n47073 );
   nand U48303 ( n47073,n45916,n47053 );
   nand U48304 ( n47072,p1_instqueue_reg_2__5_,n47054 );
   nor U48305 ( n47070,n45917,n47055 );
   nor U48306 ( n47068,n47074,n47075 );
   nor U48307 ( n47075,n45920,n47058 );
   nor U48308 ( n47074,n45921,n47059 );
   nor U48309 ( n47077,n47078,n47079 );
   nand U48310 ( n47079,n47080,n47081 );
   nand U48311 ( n47081,n45928,n47053 );
   nand U48312 ( n47080,p1_instqueue_reg_2__4_,n47054 );
   nor U48313 ( n47078,n45929,n47055 );
   nor U48314 ( n47076,n47082,n47083 );
   nor U48315 ( n47083,n45932,n47058 );
   nor U48316 ( n47082,n45933,n47059 );
   nor U48317 ( n47085,n47086,n47087 );
   nand U48318 ( n47087,n47088,n47089 );
   nand U48319 ( n47089,n45940,n47053 );
   nand U48320 ( n47088,p1_instqueue_reg_2__3_,n47054 );
   nor U48321 ( n47086,n45941,n47055 );
   nor U48322 ( n47084,n47090,n47091 );
   nor U48323 ( n47091,n45944,n47058 );
   nor U48324 ( n47090,n45945,n47059 );
   nor U48325 ( n47093,n47094,n47095 );
   nand U48326 ( n47095,n47096,n47097 );
   nand U48327 ( n47097,n45952,n47053 );
   nand U48328 ( n47096,p1_instqueue_reg_2__2_,n47054 );
   nor U48329 ( n47094,n45953,n47055 );
   nor U48330 ( n47092,n47098,n47099 );
   nor U48331 ( n47099,n45956,n47058 );
   nor U48332 ( n47098,n45957,n47059 );
   nor U48333 ( n47101,n47102,n47103 );
   nand U48334 ( n47103,n47104,n47105 );
   nand U48335 ( n47105,n45964,n47053 );
   nand U48336 ( n47104,p1_instqueue_reg_2__1_,n47054 );
   nor U48337 ( n47102,n45965,n47055 );
   nor U48338 ( n47100,n47106,n47107 );
   nor U48339 ( n47107,n45968,n47058 );
   nor U48340 ( n47106,n45969,n47059 );
   nor U48341 ( n47109,n47110,n47111 );
   nand U48342 ( n47111,n47112,n47113 );
   nand U48343 ( n47113,n45976,n47053 );
   nand U48344 ( n47053,n47114,n47115 );
   nand U48345 ( n47115,n46693,n46433 );
   nand U48346 ( n47114,n47116,n45980 );
   not U48347 ( n47116,n47117 );
   nand U48348 ( n47112,p1_instqueue_reg_2__0_,n47054 );
   nand U48349 ( n47054,n47118,n47119 );
   nand U48350 ( n47119,p1_state2_reg_3_,n47059 );
   nor U48351 ( n47118,n47120,n47121 );
   nor U48352 ( n47121,n47122,n47123 );
   nand U48353 ( n47123,n47124,n45989 );
   nand U48354 ( n47124,n45990,n47125 );
   nand U48355 ( n47125,n47058,n47055 );
   nor U48356 ( n47122,n47117,n28281 );
   nand U48357 ( n47117,n47039,n46090 );
   nor U48358 ( n47120,n47126,n28375 );
   nor U48359 ( n47126,n46445,n46785 );
   not U48360 ( n46785,n46693 );
   nor U48361 ( n46693,n47127,n46447 );
   nor U48362 ( n47110,n45999,n47055 );
   nand U48363 ( n47055,n47041,n46094 );
   nor U48364 ( n47108,n47128,n47129 );
   nor U48365 ( n47129,n46004,n47058 );
   nand U48366 ( n47058,n47044,n45407 );
   nor U48367 ( n45407,n47130,n47045 );
   nor U48368 ( n47128,n46006,n47059 );
   nand U48369 ( n47059,n47046,n46098 );
   nor U48370 ( n47132,n47133,n47134 );
   nand U48371 ( n47134,n47135,n47136 );
   nand U48372 ( n47136,n45887,n47137 );
   nand U48373 ( n47135,p1_instqueue_reg_1__7_,n47138 );
   nor U48374 ( n47133,n45890,n47139 );
   nor U48375 ( n47131,n47140,n47141 );
   nor U48376 ( n47141,n45894,n47142 );
   not U48377 ( n45894,n47143 );
   nor U48378 ( n47140,n45897,n47144 );
   nor U48379 ( n47146,n47147,n47148 );
   nand U48380 ( n47148,n47149,n47150 );
   nand U48381 ( n47150,n45904,n47137 );
   nand U48382 ( n47149,p1_instqueue_reg_1__6_,n47138 );
   nor U48383 ( n47147,n45905,n47139 );
   nor U48384 ( n47145,n47151,n47152 );
   nor U48385 ( n47152,n45908,n47142 );
   not U48386 ( n45908,n47153 );
   nor U48387 ( n47151,n45909,n47144 );
   nor U48388 ( n47155,n47156,n47157 );
   nand U48389 ( n47157,n47158,n47159 );
   nand U48390 ( n47159,n45916,n47137 );
   nand U48391 ( n47158,p1_instqueue_reg_1__5_,n47138 );
   nor U48392 ( n47156,n45917,n47139 );
   nor U48393 ( n47154,n47160,n47161 );
   nor U48394 ( n47161,n45920,n47142 );
   not U48395 ( n45920,n47162 );
   nor U48396 ( n47160,n45921,n47144 );
   nor U48397 ( n47164,n47165,n47166 );
   nand U48398 ( n47166,n47167,n47168 );
   nand U48399 ( n47168,n45928,n47137 );
   nand U48400 ( n47167,p1_instqueue_reg_1__4_,n47138 );
   nor U48401 ( n47165,n45929,n47139 );
   nor U48402 ( n47163,n47169,n47170 );
   nor U48403 ( n47170,n45932,n47142 );
   not U48404 ( n45932,n47171 );
   nor U48405 ( n47169,n45933,n47144 );
   nor U48406 ( n47173,n47174,n47175 );
   nand U48407 ( n47175,n47176,n47177 );
   nand U48408 ( n47177,n45940,n47137 );
   nand U48409 ( n47176,p1_instqueue_reg_1__3_,n47138 );
   nor U48410 ( n47174,n45941,n47139 );
   nor U48411 ( n47172,n47178,n47179 );
   nor U48412 ( n47179,n45944,n47142 );
   not U48413 ( n45944,n47180 );
   nor U48414 ( n47178,n45945,n47144 );
   nor U48415 ( n47182,n47183,n47184 );
   nand U48416 ( n47184,n47185,n47186 );
   nand U48417 ( n47186,n45952,n47137 );
   nand U48418 ( n47185,p1_instqueue_reg_1__2_,n47138 );
   nor U48419 ( n47183,n45953,n47139 );
   nor U48420 ( n47181,n47187,n47188 );
   nor U48421 ( n47188,n45956,n47142 );
   not U48422 ( n45956,n47189 );
   nor U48423 ( n47187,n45957,n47144 );
   nor U48424 ( n47191,n47192,n47193 );
   nand U48425 ( n47193,n47194,n47195 );
   nand U48426 ( n47195,n45964,n47137 );
   nand U48427 ( n47194,p1_instqueue_reg_1__1_,n47138 );
   nor U48428 ( n47192,n45965,n47139 );
   nor U48429 ( n47190,n47196,n47197 );
   nor U48430 ( n47197,n45968,n47142 );
   not U48431 ( n45968,n47198 );
   nor U48432 ( n47196,n45969,n47144 );
   nor U48433 ( n47200,n47201,n47202 );
   nand U48434 ( n47202,n47203,n47204 );
   nand U48435 ( n47204,n45976,n47137 );
   nand U48436 ( n47137,n47205,n47206 );
   nand U48437 ( n47206,p1_state2_reg_2_,n47207 );
   nand U48438 ( n47205,n47208,n45980 );
   nand U48439 ( n47203,p1_instqueue_reg_1__0_,n47138 );
   nand U48440 ( n47138,n47209,n47210 );
   nand U48441 ( n47210,p1_state2_reg_3_,n47144 );
   nor U48442 ( n47209,n47211,n47212 );
   nor U48443 ( n47212,n47213,n47214 );
   nand U48444 ( n47214,n47215,n45989 );
   nand U48445 ( n47215,n45990,n47216 );
   nand U48446 ( n47216,n47142,n47139 );
   and U48447 ( n47213,n47208,n45992 );
   nand U48448 ( n47208,n47144,n47217 );
   nand U48449 ( n47217,n47039,n46179 );
   nor U48450 ( n46179,n45394,n46090 );
   nor U48451 ( n47211,n28374,n47207 );
   nand U48452 ( n47207,n47144,n47218 );
   nand U48453 ( n47218,n46872,n46358 );
   nor U48454 ( n46358,n46445,p1_instqueuewr_addr_reg_0_ );
   nor U48455 ( n47201,n45999,n47139 );
   nand U48456 ( n47139,n47041,n46182 );
   nor U48457 ( n47199,n47219,n47220 );
   nor U48458 ( n47220,n46004,n47142 );
   nand U48459 ( n47142,n47044,n45408 );
   nor U48460 ( n45408,n47221,n45389 );
   not U48461 ( n46004,n47222 );
   nor U48462 ( n47219,n46006,n47144 );
   nand U48463 ( n47144,n47046,n46185 );
   nor U48464 ( n47224,n47225,n47226 );
   nand U48465 ( n47226,n47227,n47228 );
   nand U48466 ( n47228,n47229,n47143 );
   nand U48467 ( n47143,n47230,n47231 );
   nand U48468 ( n47231,datai_31_,n47232 );
   nand U48469 ( n47230,n47233,buf1_reg_31_ );
   or U48470 ( n47227,n47234,n28189 );
   nand U48471 ( n45897,n47235,n47236 );
   nor U48472 ( n47225,n28192,n47237 );
   and U48473 ( n45890,n47238,n47239 );
   nand U48474 ( n47239,datai_23_,n47232 );
   nand U48475 ( n47238,n47233,buf1_reg_23_ );
   nor U48476 ( n47223,n47240,n47241 );
   nor U48477 ( n47241,n47242,n47243 );
   nor U48478 ( n47240,n47244,n47245 );
   not U48479 ( n47245,n45887 );
   nor U48480 ( n45887,n46089,n47246 );
   nor U48481 ( n47248,n47249,n47250 );
   nand U48482 ( n47250,n47251,n47252 );
   nand U48483 ( n47252,n47229,n47153 );
   nand U48484 ( n47153,n47253,n47254 );
   nand U48485 ( n47254,datai_30_,n47232 );
   nand U48486 ( n47253,n47233,buf1_reg_30_ );
   or U48487 ( n47251,n47234,n28194 );
   nand U48488 ( n45909,n47235,n47255 );
   nor U48489 ( n47249,n28198,n47237 );
   and U48490 ( n45905,n47256,n47257 );
   nand U48491 ( n47257,datai_22_,n47232 );
   nand U48492 ( n47256,n47233,buf1_reg_22_ );
   nor U48493 ( n47247,n47258,n47259 );
   nor U48494 ( n47259,n47242,n47260 );
   nor U48495 ( n47258,n47244,n47261 );
   not U48496 ( n47261,n45904 );
   nor U48497 ( n45904,n47262,n28281 );
   nor U48498 ( n47264,n47265,n47266 );
   nand U48499 ( n47266,n47267,n47268 );
   nand U48500 ( n47268,n47229,n47162 );
   nand U48501 ( n47162,n47269,n47270 );
   nand U48502 ( n47270,datai_29_,n47232 );
   nand U48503 ( n47269,n47233,buf1_reg_29_ );
   or U48504 ( n47267,n47234,n28200 );
   nand U48505 ( n45921,n47235,n47271 );
   nor U48506 ( n47265,n28204,n47237 );
   and U48507 ( n45917,n47272,n47273 );
   nand U48508 ( n47273,datai_21_,n47232 );
   nand U48509 ( n47272,n47233,buf1_reg_21_ );
   nor U48510 ( n47263,n47274,n47275 );
   nor U48511 ( n47275,n47242,n47276 );
   nor U48512 ( n47274,n47244,n47277 );
   not U48513 ( n47277,n45916 );
   nor U48514 ( n45916,n47278,n46089 );
   nor U48515 ( n47280,n47281,n47282 );
   nand U48516 ( n47282,n47283,n47284 );
   nand U48517 ( n47284,n47229,n47171 );
   nand U48518 ( n47171,n47285,n47286 );
   nand U48519 ( n47286,datai_28_,n47232 );
   nand U48520 ( n47285,n47233,buf1_reg_28_ );
   or U48521 ( n47283,n47234,n28207 );
   nand U48522 ( n45933,n47235,n47287 );
   nor U48523 ( n47281,n28211,n47237 );
   and U48524 ( n45929,n47288,n47289 );
   nand U48525 ( n47289,datai_20_,n47232 );
   nand U48526 ( n47288,n47233,buf1_reg_20_ );
   nor U48527 ( n47279,n47290,n47291 );
   nor U48528 ( n47291,n47242,n47292 );
   nor U48529 ( n47290,n47244,n47293 );
   not U48530 ( n47293,n45928 );
   nor U48531 ( n45928,n47294,n28281 );
   nor U48532 ( n47296,n47297,n47298 );
   nand U48533 ( n47298,n47299,n47300 );
   nand U48534 ( n47300,n47229,n47180 );
   nand U48535 ( n47180,n47301,n47302 );
   nand U48536 ( n47302,datai_27_,n47232 );
   nand U48537 ( n47301,n47233,buf1_reg_27_ );
   or U48538 ( n47299,n47234,n28215 );
   nand U48539 ( n45945,n47235,n47303 );
   nor U48540 ( n47297,n28219,n47237 );
   and U48541 ( n45941,n47304,n47305 );
   nand U48542 ( n47305,datai_19_,n47232 );
   nand U48543 ( n47304,n47233,buf1_reg_19_ );
   nor U48544 ( n47295,n47306,n47307 );
   nor U48545 ( n47307,n47242,n47308 );
   nor U48546 ( n47306,n47244,n47309 );
   not U48547 ( n47309,n45940 );
   nor U48548 ( n45940,n47310,n28281 );
   nor U48549 ( n47312,n47313,n47314 );
   nand U48550 ( n47314,n47315,n47316 );
   nand U48551 ( n47316,n47229,n47189 );
   nand U48552 ( n47189,n47317,n47318 );
   nand U48553 ( n47318,datai_26_,n47232 );
   nand U48554 ( n47317,n47233,buf1_reg_26_ );
   or U48555 ( n47315,n47234,n28227 );
   nand U48556 ( n45957,n47235,n45878 );
   nor U48557 ( n47313,n28231,n47237 );
   and U48558 ( n45953,n47319,n47320 );
   nand U48559 ( n47320,datai_18_,n47232 );
   nand U48560 ( n47319,n47233,buf1_reg_18_ );
   nor U48561 ( n47311,n47321,n47322 );
   nor U48562 ( n47322,n47242,n47323 );
   nor U48563 ( n47321,n47244,n47324 );
   not U48564 ( n47324,n45952 );
   nor U48565 ( n45952,n47325,n28281 );
   nor U48566 ( n47327,n47328,n47329 );
   nand U48567 ( n47329,n47330,n47331 );
   nand U48568 ( n47331,n47229,n47198 );
   nand U48569 ( n47198,n47332,n47333 );
   nand U48570 ( n47333,datai_25_,n47232 );
   nand U48571 ( n47332,n47233,buf1_reg_25_ );
   or U48572 ( n47330,n47234,n28245 );
   nand U48573 ( n45969,n47235,n47334 );
   nor U48574 ( n47328,n28249,n47237 );
   and U48575 ( n45965,n47335,n47336 );
   nand U48576 ( n47336,datai_17_,n47232 );
   nand U48577 ( n47335,n47233,buf1_reg_17_ );
   nor U48578 ( n47326,n47337,n47338 );
   nor U48579 ( n47338,n47242,n47339 );
   nor U48580 ( n47337,n47244,n47340 );
   not U48581 ( n47340,n45964 );
   nor U48582 ( n45964,n47341,n28281 );
   nor U48583 ( n47343,n47344,n47345 );
   nand U48584 ( n47345,n47346,n47347 );
   nand U48585 ( n47347,n47229,n47222 );
   nand U48586 ( n47222,n47348,n47349 );
   nand U48587 ( n47349,datai_24_,n47232 );
   nand U48588 ( n47348,n47233,buf1_reg_24_ );
   not U48589 ( n47229,n47350 );
   or U48590 ( n47346,n47234,n28325 );
   nand U48591 ( n46006,n47235,n27892 );
   nor U48592 ( n47235,n46089,n45501 );
   nor U48593 ( n47344,n28273,n47237 );
   and U48594 ( n45999,n47352,n47353 );
   nand U48595 ( n47353,datai_16_,n47232 );
   nor U48596 ( n47232,n47354,n47355 );
   nand U48597 ( n47352,n47233,buf1_reg_16_ );
   nor U48598 ( n47233,n47354,n28765 );
   nor U48599 ( n47342,n47356,n47357 );
   nor U48600 ( n47357,n47244,n47358 );
   not U48601 ( n47358,n45976 );
   nor U48602 ( n45976,n47359,n28281 );
   and U48603 ( n47244,n47360,n47361 );
   nand U48604 ( n47361,n46872,n46433 );
   nor U48605 ( n46433,n46445,n45355 );
   nand U48606 ( n47360,n45980,n47362 );
   not U48607 ( n47362,n47363 );
   nand U48608 ( n45980,n46697,n45406 );
   nor U48609 ( n47356,n47242,n47364 );
   and U48610 ( n47242,n47365,n47366 );
   nand U48611 ( n47366,p1_state2_reg_3_,n47234 );
   nand U48612 ( n47234,n47046,n46274 );
   nor U48613 ( n46274,p1_instqueuewr_addr_reg_1_,p1_instqueuewr_addr_reg_0_ );
   nor U48614 ( n47046,p1_instqueuewr_addr_reg_3_,p1_instqueuewr_addr_reg_2_ );
   nor U48615 ( n47365,n47367,n47368 );
   nor U48616 ( n47368,n47369,n47370 );
   nand U48617 ( n47370,n47371,n45989 );
   or U48618 ( n45989,n46696,n28281 );
   nand U48619 ( n46696,n46697,n47354 );
   or U48620 ( n47354,n46089,n45406 );
   nand U48621 ( n45406,p1_statebs16_reg,n45341 );
   nand U48622 ( n47371,n45990,n47372 );
   nand U48623 ( n47372,n47350,n47237 );
   nand U48624 ( n47237,n47041,n46267 );
   nor U48625 ( n46267,n45389,n45401 );
   nor U48626 ( n47041,n45414,n45428 );
   nand U48627 ( n47350,n47044,n46272 );
   nor U48628 ( n46272,n47221,n47130 );
   not U48629 ( n47221,n47045 );
   nor U48630 ( n47045,n46094,n46182 );
   nor U48631 ( n46182,n45401,n47130 );
   nor U48632 ( n46094,n45389,n47373 );
   nor U48633 ( n47044,n46005,n45421 );
   not U48634 ( n45421,n46273 );
   xor U48635 ( n46273,n46001,n46269 );
   nand U48636 ( n46005,n47374,n47375 );
   or U48637 ( n47375,n46268,n46001 );
   nor U48638 ( n47374,n46359,n47376 );
   not U48639 ( n47376,n46628 );
   nand U48640 ( n46628,n46786,n46001 );
   nor U48641 ( n46001,n47373,n47130 );
   nor U48642 ( n46786,n45428,n46269 );
   nor U48643 ( n46359,n46268,n45414 );
   nor U48644 ( n45990,n46089,n45400 );
   not U48645 ( n45400,n46697 );
   nand U48646 ( n46697,n45341,n47377 );
   nor U48647 ( n47369,n47363,n28281 );
   nand U48648 ( n47363,n47039,n45404 );
   nor U48649 ( n47039,n46612,n46954 );
   nor U48650 ( n47367,n47378,n45355 );
   nor U48651 ( n47378,n46445,n46956 );
   not U48652 ( n46956,n46872 );
   nor U48653 ( n46872,n47127,n46614 );
   not U48654 ( n46614,n46447 );
   not U48655 ( n45384,n45386 );
   nand U48656 ( n45386,n47379,n47380 );
   nand U48657 ( n47380,n45780,n45392 );
   nand U48658 ( n45392,n45858,n47381 );
   nand U48659 ( n47381,n47382,n45860 );
   nand U48660 ( n45860,n47383,n47384 );
   nand U48661 ( n47384,n47385,p1_instqueuerd_addr_reg_3_ );
   nand U48662 ( n47383,n45854,n45432 );
   nand U48663 ( n45854,n47386,n47387 );
   nand U48664 ( n47387,n45497,p1_instqueuerd_addr_reg_3_ );
   nand U48665 ( n47386,n45487,n45826 );
   nand U48666 ( n45487,n47388,n47389 );
   nor U48667 ( n47389,n47390,n47391 );
   nor U48668 ( n47391,n47392,n47393 );
   nor U48669 ( n47390,n47394,n47395 );
   nor U48670 ( n47394,n47396,n47397 );
   nor U48671 ( n47397,p1_instqueuerd_addr_reg_3_,n47398 );
   nor U48672 ( n47398,n47399,n47400 );
   nor U48673 ( n47396,n47399,n47401 );
   nand U48674 ( n47401,n47400,n47402 );
   not U48675 ( n47400,n47403 );
   nor U48676 ( n47388,n47404,n47405 );
   nor U48677 ( n47405,n45836,n47406 );
   nor U48678 ( n47404,n45850,n45431 );
   not U48679 ( n45431,n46954 );
   and U48680 ( n47382,n47407,n45861 );
   nand U48681 ( n45861,n47408,n47409 );
   nand U48682 ( n47409,n47410,n45813 );
   not U48683 ( n45813,n45841 );
   nor U48684 ( n45841,n45826,p1_instqueuerd_addr_reg_2_ );
   nor U48685 ( n47410,p1_state2_reg_1_,n45814 );
   and U48686 ( n45814,n45475,n45826 );
   and U48687 ( n45475,n47411,n47412 );
   nor U48688 ( n47412,n47413,n47414 );
   nor U48689 ( n47414,n47395,n45472 );
   nor U48690 ( n47395,n47415,n47416 );
   nor U48691 ( n47413,n47417,n47393 );
   nand U48692 ( n47393,n47418,n47419 );
   nor U48693 ( n47418,n47334,n47420 );
   nor U48694 ( n47411,n47421,n47422 );
   nor U48695 ( n47422,n47423,n45836 );
   nor U48696 ( n47421,n45850,n45417 );
   not U48697 ( n45850,n45835 );
   nand U48698 ( n45835,n47424,n47425 );
   nor U48699 ( n47425,n47426,n47427 );
   nand U48700 ( n47427,n47428,n47429 );
   nor U48701 ( n47424,n47430,n47431 );
   nand U48702 ( n47431,n47432,n47433 );
   nand U48703 ( n47408,n47385,p1_instqueuerd_addr_reg_2_ );
   and U48704 ( n45858,n47434,n47435 );
   nand U48705 ( n47435,n47436,n45432 );
   nand U48706 ( n47436,n45492,n47437 );
   nand U48707 ( n47437,n45497,p1_instqueuerd_addr_reg_4_ );
   not U48708 ( n45497,n45826 );
   nand U48709 ( n45826,n47438,n47439 );
   nor U48710 ( n47439,n47440,n47441 );
   nand U48711 ( n47441,n47442,n47443 );
   nand U48712 ( n47442,n47444,n45864 );
   nor U48713 ( n47440,n47351,n47445 );
   nand U48714 ( n47445,n47446,n47334 );
   nor U48715 ( n47438,n47447,n47448 );
   nand U48716 ( n47448,n47449,n47450 );
   nand U48717 ( n47449,n47451,n45869 );
   nand U48718 ( n47451,n45872,n47452 );
   nand U48719 ( n47452,n47453,n45346 );
   nand U48720 ( n47453,n47454,n47455 );
   nand U48721 ( n47455,n45360,n47456 );
   nand U48722 ( n47456,n47433,n45836 );
   not U48723 ( n47454,n47457 );
   nand U48724 ( n45492,n45864,n47458 );
   nand U48725 ( n47434,n47385,p1_instqueuerd_addr_reg_4_ );
   nor U48726 ( n47385,n45432,p1_flush_reg );
   nor U48727 ( n47379,n45495,n45992 );
   not U48728 ( n45992,n46089 );
   nand U48729 ( n46089,n45347,n47459 );
   nand U48730 ( n47459,n47460,n45757 );
   nand U48731 ( n45757,p1_state2_reg_1_,n45355 );
   nor U48732 ( n47460,n45759,n45452 );
   nor U48733 ( n45452,n45501,n45880 );
   and U48734 ( n45495,p1_flush_reg,n45780 );
   nor U48735 ( n45780,n45344,n28094 );
   not U48736 ( n45344,n45503 );
   nor U48737 ( n47462,n47463,n47464 );
   nor U48738 ( n47464,n45373,n47465 );
   nor U48739 ( n47463,n28305,n47467 );
   nor U48740 ( n47461,n47468,n47469 );
   nand U48741 ( n47469,n47470,n47471 );
   nand U48742 ( n47470,p1_instaddrpointer_reg_0_,n47472 );
   nand U48743 ( n47472,n47473,n28253 );
   nor U48744 ( n47468,n28293,n47475 );
   nor U48745 ( n47477,n47478,n47479 );
   nand U48746 ( n47479,n47480,n47481 );
   not U48747 ( n47481,n47482 );
   or U48748 ( n47480,n47483,n28305 );
   nor U48749 ( n47478,n45674,n47465 );
   nor U48750 ( n47476,n47484,n47485 );
   nand U48751 ( n47485,n47486,n47487 );
   nand U48752 ( n47487,p1_instaddrpointer_reg_1_,n47488 );
   nand U48753 ( n47488,n47473,n47471 );
   nand U48754 ( n47471,n47489,n45448 );
   not U48755 ( n47489,n47490 );
   nand U48756 ( n47486,n47491,n45479 );
   nor U48757 ( n47491,n47490,n45448 );
   nor U48758 ( n47484,n28294,n47492 );
   nor U48759 ( n47494,n47495,n47496 );
   nand U48760 ( n47496,n47497,n47498 );
   nand U48761 ( n47498,n47499,n47500 );
   nand U48762 ( n47500,n47501,n47502 );
   nand U48763 ( n47497,n47503,n28213 );
   nor U48764 ( n47495,n45669,n28113 );
   nor U48765 ( n47493,n47505,n47506 );
   nand U48766 ( n47506,n47507,n47508 );
   nand U48767 ( n47508,p1_instaddrpointer_reg_2_,n47509 );
   nand U48768 ( n47509,n47510,n47511 );
   nand U48769 ( n47511,n47512,n47513 );
   nor U48770 ( n47510,n47514,n47482 );
   nand U48771 ( n47507,n47515,n47516 );
   nor U48772 ( n47515,n47517,n45479 );
   nor U48773 ( n47517,n47518,n47519 );
   nor U48774 ( n47518,n45448,n47520 );
   nor U48775 ( n47505,n28296,n47521 );
   nor U48776 ( n47523,n47524,n47525 );
   nor U48777 ( n47525,n45664,n28114 );
   nor U48778 ( n47524,n47466,n47526 );
   nor U48779 ( n47522,n47527,n47528 );
   nand U48780 ( n47528,n47529,n47530 );
   nand U48781 ( n47530,p1_instaddrpointer_reg_3_,n47531 );
   nand U48782 ( n47531,n47532,n47533 );
   nor U48783 ( n47532,n47482,n47534 );
   nor U48784 ( n47534,p1_instaddrpointer_reg_2_,n47474 );
   nor U48785 ( n47482,n28253,p1_instaddrpointer_reg_1_ );
   nand U48786 ( n47529,n47535,n47536 );
   nand U48787 ( n47535,n47537,n47538 );
   nand U48788 ( n47538,n47539,p1_instaddrpointer_reg_2_ );
   nor U48789 ( n47539,n45479,n47474 );
   not U48790 ( n47537,n47540 );
   nor U48791 ( n47527,n28296,n47541 );
   nor U48792 ( n47543,n47544,n47545 );
   nor U48793 ( n47545,n45659,n47465 );
   nor U48794 ( n47544,n28305,n47546 );
   nor U48795 ( n47542,n47547,n47548 );
   nand U48796 ( n47548,n47549,n47550 );
   nand U48797 ( n47550,p1_instaddrpointer_reg_4_,n47551 );
   nand U48798 ( n47551,n47552,n47533 );
   and U48799 ( n47533,n47553,n47554 );
   nand U48800 ( n47554,n47555,n47499 );
   nor U48801 ( n47553,n47514,n47556 );
   nor U48802 ( n47556,n47557,n47520 );
   nor U48803 ( n47552,n47558,n47559 );
   nor U48804 ( n47559,p1_instaddrpointer_reg_3_,n47490 );
   nor U48805 ( n47558,n47560,n28253 );
   nand U48806 ( n47549,n47561,n47562 );
   nand U48807 ( n47561,n47563,n47564 );
   nand U48808 ( n47564,p1_instaddrpointer_reg_3_,n47540 );
   nand U48809 ( n47540,n47565,n47566 );
   nand U48810 ( n47566,n47557,n47512 );
   nand U48811 ( n47565,n47499,n47501 );
   not U48812 ( n47501,n47555 );
   nand U48813 ( n47563,n47560,n28338 );
   nor U48814 ( n47547,n28293,n47567 );
   nor U48815 ( n47569,n47570,n47571 );
   nor U48816 ( n47571,n45654,n28113 );
   nor U48817 ( n47570,n28305,n47572 );
   nor U48818 ( n47568,n47573,n47574 );
   nand U48819 ( n47574,n47575,n47576 );
   nand U48820 ( n47576,p1_instaddrpointer_reg_5_,n47577 );
   nand U48821 ( n47577,n47578,n47579 );
   nand U48822 ( n47579,n47519,n47580 );
   nand U48823 ( n47575,n47581,n47582 );
   nand U48824 ( n47581,n47583,n47584 );
   or U48825 ( n47584,n47580,n47474 );
   not U48826 ( n47583,n47585 );
   nor U48827 ( n47573,n28293,n47586 );
   nor U48828 ( n47588,n47589,n47590 );
   nor U48829 ( n47590,n45649,n28114 );
   nor U48830 ( n47589,n47466,n47591 );
   nor U48831 ( n47587,n47592,n47593 );
   nand U48832 ( n47593,n47594,n47595 );
   nand U48833 ( n47595,p1_instaddrpointer_reg_6_,n47596 );
   nand U48834 ( n47596,n47597,n47578 );
   and U48835 ( n47578,n47598,n47599 );
   nand U48836 ( n47599,n47499,n47600 );
   nor U48837 ( n47598,n47514,n47601 );
   nor U48838 ( n47601,n47602,n47520 );
   nor U48839 ( n47597,n47603,n47604 );
   nor U48840 ( n47604,p1_instaddrpointer_reg_5_,n47490 );
   nor U48841 ( n47603,n47605,n47474 );
   nand U48842 ( n47594,n47606,n47607 );
   nand U48843 ( n47606,n47608,n47609 );
   nand U48844 ( n47609,p1_instaddrpointer_reg_5_,n47585 );
   nand U48845 ( n47585,n47610,n47611 );
   nand U48846 ( n47611,n47602,n47512 );
   not U48847 ( n47602,n47612 );
   or U48848 ( n47610,n47600,n47613 );
   nand U48849 ( n47608,n47605,n28338 );
   nor U48850 ( n47592,n28295,n47614 );
   nor U48851 ( n47616,n47617,n47618 );
   nor U48852 ( n47618,n45644,n47465 );
   nor U48853 ( n47617,n47466,n47619 );
   nor U48854 ( n47615,n47620,n47621 );
   nand U48855 ( n47621,n47622,n47623 );
   nand U48856 ( n47623,p1_instaddrpointer_reg_7_,n47624 );
   nand U48857 ( n47624,n47625,n47626 );
   nand U48858 ( n47626,n47519,n47627 );
   nand U48859 ( n47622,n47628,n47629 );
   nand U48860 ( n47628,n47630,n47631 );
   or U48861 ( n47631,n47627,n47474 );
   not U48862 ( n47630,n47632 );
   nor U48863 ( n47620,n28295,n47633 );
   nor U48864 ( n47635,n47636,n47637 );
   nor U48865 ( n47637,n45639,n28113 );
   and U48866 ( n47636,n47504,n47638 );
   nor U48867 ( n47634,n47639,n47640 );
   nand U48868 ( n47640,n47641,n47642 );
   nand U48869 ( n47642,p1_instaddrpointer_reg_8_,n47643 );
   nand U48870 ( n47643,n47644,n47625 );
   and U48871 ( n47625,n47645,n47646 );
   nand U48872 ( n47646,n47499,n47647 );
   nor U48873 ( n47645,n28232,n47648 );
   nor U48874 ( n47648,n47649,n47520 );
   nor U48875 ( n47644,n47650,n47651 );
   nor U48876 ( n47651,p1_instaddrpointer_reg_7_,n47490 );
   nor U48877 ( n47650,n47652,n28253 );
   nand U48878 ( n47641,n47653,n47654 );
   nand U48879 ( n47653,n47655,n47656 );
   nand U48880 ( n47656,p1_instaddrpointer_reg_7_,n47632 );
   nand U48881 ( n47632,n47657,n47658 );
   nand U48882 ( n47658,n47649,n47512 );
   not U48883 ( n47649,n47659 );
   or U48884 ( n47657,n47647,n47613 );
   nand U48885 ( n47655,n47652,n28338 );
   nor U48886 ( n47639,n28294,n47660 );
   nor U48887 ( n47662,n47663,n47664 );
   nor U48888 ( n47664,n45634,n28114 );
   and U48889 ( n47663,n47504,n47665 );
   nor U48890 ( n47661,n47666,n47667 );
   nand U48891 ( n47667,n47668,n47669 );
   nand U48892 ( n47669,p1_instaddrpointer_reg_9_,n47670 );
   nand U48893 ( n47670,n47671,n47672 );
   nand U48894 ( n47672,n47519,n47673 );
   nand U48895 ( n47668,n47674,n47675 );
   nand U48896 ( n47674,n47676,n47677 );
   or U48897 ( n47677,n47673,n28253 );
   not U48898 ( n47676,n47678 );
   nor U48899 ( n47666,n28294,n47679 );
   nor U48900 ( n47681,n47682,n47683 );
   nor U48901 ( n47683,n45629,n47465 );
   and U48902 ( n47682,n28213,n47684 );
   nor U48903 ( n47680,n47685,n47686 );
   nand U48904 ( n47686,n47687,n47688 );
   nand U48905 ( n47688,p1_instaddrpointer_reg_10_,n47689 );
   nand U48906 ( n47689,n47690,n47671 );
   and U48907 ( n47671,n47691,n47692 );
   nand U48908 ( n47692,n47499,n47693 );
   nor U48909 ( n47691,n47514,n47694 );
   nor U48910 ( n47694,n47695,n28205 );
   nor U48911 ( n47690,n47696,n47697 );
   nor U48912 ( n47697,p1_instaddrpointer_reg_9_,n28238 );
   nor U48913 ( n47696,n47698,n28253 );
   nand U48914 ( n47687,n47699,n47700 );
   not U48915 ( n47700,p1_instaddrpointer_reg_10_ );
   nand U48916 ( n47699,n47701,n47702 );
   nand U48917 ( n47702,p1_instaddrpointer_reg_9_,n47678 );
   nand U48918 ( n47678,n47703,n47704 );
   nand U48919 ( n47704,n47695,n47512 );
   not U48920 ( n47695,n47705 );
   or U48921 ( n47703,n47693,n47613 );
   nand U48922 ( n47701,n47698,n28338 );
   nor U48923 ( n47685,n28296,n47706 );
   nor U48924 ( n47708,n47709,n47710 );
   nor U48925 ( n47710,n45624,n28113 );
   nor U48926 ( n47709,n47711,n47712 );
   nand U48927 ( n47712,n47713,n28213 );
   nor U48928 ( n47707,n47714,n47715 );
   nand U48929 ( n47715,n47716,n47717 );
   nand U48930 ( n47717,p1_instaddrpointer_reg_11_,n47718 );
   nand U48931 ( n47718,n47719,n47720 );
   nand U48932 ( n47720,n47519,n47721 );
   nand U48933 ( n47716,n47722,n47723 );
   nand U48934 ( n47722,n47724,n47725 );
   or U48935 ( n47725,n47721,n47474 );
   not U48936 ( n47724,n47726 );
   nor U48937 ( n47714,n28296,n47727 );
   nor U48938 ( n47729,n47730,n47731 );
   nor U48939 ( n47731,n45619,n28114 );
   and U48940 ( n47730,n47504,n47732 );
   nor U48941 ( n47728,n47733,n47734 );
   nand U48942 ( n47734,n47735,n47736 );
   nand U48943 ( n47736,p1_instaddrpointer_reg_12_,n47737 );
   nand U48944 ( n47737,n47738,n47719 );
   and U48945 ( n47719,n47739,n47740 );
   nand U48946 ( n47740,n47499,n47741 );
   nor U48947 ( n47739,n47514,n47742 );
   nor U48948 ( n47742,n47743,n28205 );
   nor U48949 ( n47738,n47744,n47745 );
   nor U48950 ( n47745,p1_instaddrpointer_reg_11_,n47490 );
   nor U48951 ( n47744,n47746,n47474 );
   nand U48952 ( n47735,n47747,n47748 );
   nand U48953 ( n47747,n47749,n47750 );
   nand U48954 ( n47750,p1_instaddrpointer_reg_11_,n47726 );
   nand U48955 ( n47726,n47751,n47752 );
   nand U48956 ( n47752,n47743,n47512 );
   not U48957 ( n47743,n47753 );
   or U48958 ( n47751,n47741,n47613 );
   nand U48959 ( n47749,n47746,n28338 );
   nor U48960 ( n47733,n28294,n47754 );
   nor U48961 ( n47756,n47757,n47758 );
   nor U48962 ( n47758,n45614,n28113 );
   and U48963 ( n47757,n47504,n47759 );
   nor U48964 ( n47755,n47760,n47761 );
   nand U48965 ( n47761,n47762,n47763 );
   nand U48966 ( n47763,p1_instaddrpointer_reg_13_,n47764 );
   nand U48967 ( n47764,n47765,n47766 );
   nand U48968 ( n47766,n28338,n47767 );
   nand U48969 ( n47762,n47768,n47769 );
   nand U48970 ( n47768,n47770,n47771 );
   or U48971 ( n47771,n47767,n47474 );
   not U48972 ( n47770,n47772 );
   nor U48973 ( n47760,n28295,n47773 );
   nor U48974 ( n47775,n47776,n47777 );
   nor U48975 ( n47777,n45609,n47465 );
   nor U48976 ( n47776,n47466,n47778 );
   nor U48977 ( n47774,n47779,n47780 );
   nand U48978 ( n47780,n47781,n47782 );
   nand U48979 ( n47782,p1_instaddrpointer_reg_14_,n47783 );
   nand U48980 ( n47783,n47784,n47765 );
   and U48981 ( n47765,n47785,n47786 );
   nand U48982 ( n47786,n47499,n47787 );
   nor U48983 ( n47785,n47514,n47788 );
   nor U48984 ( n47788,n47789,n47520 );
   nor U48985 ( n47784,n47790,n47791 );
   nor U48986 ( n47791,p1_instaddrpointer_reg_13_,n47490 );
   nor U48987 ( n47790,n47792,n47474 );
   nand U48988 ( n47781,n47793,n47794 );
   nand U48989 ( n47793,n47795,n47796 );
   nand U48990 ( n47796,p1_instaddrpointer_reg_13_,n47772 );
   nand U48991 ( n47772,n47797,n47798 );
   nand U48992 ( n47798,n47789,n47512 );
   not U48993 ( n47789,n47799 );
   or U48994 ( n47797,n47787,n47613 );
   nand U48995 ( n47795,n47792,n28338 );
   nor U48996 ( n47779,n28295,n47800 );
   nor U48997 ( n47802,n47803,n47804 );
   nor U48998 ( n47804,n45604,n28114 );
   nor U48999 ( n47803,n47805,n47806 );
   nand U49000 ( n47806,n47807,n28213 );
   nor U49001 ( n47801,n47808,n47809 );
   nand U49002 ( n47809,n47810,n47811 );
   nand U49003 ( n47811,p1_instaddrpointer_reg_15_,n47812 );
   nand U49004 ( n47812,n47813,n47814 );
   nand U49005 ( n47814,n47519,n47815 );
   nand U49006 ( n47810,n47816,n47817 );
   nand U49007 ( n47816,n47818,n47819 );
   or U49008 ( n47819,n47815,n28253 );
   not U49009 ( n47818,n47820 );
   nor U49010 ( n47808,n28293,n47821 );
   nor U49011 ( n47823,n47824,n47825 );
   nor U49012 ( n47825,n45599,n28113 );
   and U49013 ( n47824,n47504,n47826 );
   nor U49014 ( n47822,n47827,n47828 );
   nand U49015 ( n47828,n47829,n47830 );
   nand U49016 ( n47830,p1_instaddrpointer_reg_16_,n47831 );
   nand U49017 ( n47831,n47832,n47813 );
   and U49018 ( n47813,n47833,n47834 );
   nand U49019 ( n47834,n47499,n47835 );
   nor U49020 ( n47833,n47514,n47836 );
   nor U49021 ( n47836,n47837,n47520 );
   nor U49022 ( n47832,n47838,n47839 );
   nor U49023 ( n47839,p1_instaddrpointer_reg_15_,n47490 );
   nor U49024 ( n47838,n47840,n28253 );
   nand U49025 ( n47829,n47841,n47842 );
   nand U49026 ( n47841,n47843,n47844 );
   nand U49027 ( n47844,p1_instaddrpointer_reg_15_,n47820 );
   nand U49028 ( n47820,n47845,n47846 );
   nand U49029 ( n47846,n47837,n47512 );
   not U49030 ( n47837,n47847 );
   or U49031 ( n47845,n47835,n47613 );
   nand U49032 ( n47843,n47840,n28338 );
   nor U49033 ( n47827,n28293,n47848 );
   nor U49034 ( n47850,n47851,n47852 );
   nor U49035 ( n47852,n45594,n47465 );
   nor U49036 ( n47851,n47466,n47853 );
   nor U49037 ( n47849,n47854,n47855 );
   nand U49038 ( n47855,n47856,n47857 );
   nand U49039 ( n47857,p1_instaddrpointer_reg_17_,n47858 );
   nand U49040 ( n47858,n47859,n47860 );
   nand U49041 ( n47860,n47519,n47861 );
   nand U49042 ( n47856,n47862,n47863 );
   nand U49043 ( n47862,n47864,n47865 );
   or U49044 ( n47865,n47861,n28253 );
   not U49045 ( n47864,n47866 );
   nor U49046 ( n47854,n28296,n47867 );
   nor U49047 ( n47869,n47870,n47871 );
   nor U49048 ( n47871,n45589,n28114 );
   nor U49049 ( n47870,n47466,n47872 );
   nor U49050 ( n47868,n47873,n47874 );
   nand U49051 ( n47874,n47875,n47876 );
   nand U49052 ( n47876,p1_instaddrpointer_reg_18_,n47877 );
   nand U49053 ( n47877,n47878,n47859 );
   and U49054 ( n47859,n47879,n47880 );
   nand U49055 ( n47880,n47499,n47881 );
   nor U49056 ( n47879,n47514,n47882 );
   nor U49057 ( n47882,n47883,n47520 );
   nor U49058 ( n47878,n47884,n47885 );
   nor U49059 ( n47885,p1_instaddrpointer_reg_17_,n47490 );
   nor U49060 ( n47884,n47886,n28253 );
   nand U49061 ( n47875,n47887,n47888 );
   not U49062 ( n47888,p1_instaddrpointer_reg_18_ );
   nand U49063 ( n47887,n47889,n47890 );
   nand U49064 ( n47890,p1_instaddrpointer_reg_17_,n47866 );
   nand U49065 ( n47866,n47891,n47892 );
   nand U49066 ( n47892,n47883,n47512 );
   not U49067 ( n47883,n47893 );
   or U49068 ( n47891,n47881,n47613 );
   nand U49069 ( n47889,n47886,n28338 );
   nor U49070 ( n47873,n28296,n47894 );
   nor U49071 ( n47896,n47897,n47898 );
   nor U49072 ( n47898,n45584,n28113 );
   and U49073 ( n47897,n47504,n47899 );
   nor U49074 ( n47895,n47900,n47901 );
   nand U49075 ( n47901,n47902,n47903 );
   nand U49076 ( n47903,p1_instaddrpointer_reg_19_,n47904 );
   nand U49077 ( n47904,n47905,n47906 );
   nand U49078 ( n47906,n47519,n47907 );
   nand U49079 ( n47902,n47908,n47909 );
   nand U49080 ( n47908,n47910,n47911 );
   or U49081 ( n47911,n47907,n28253 );
   not U49082 ( n47910,n47912 );
   nor U49083 ( n47900,n28294,n47913 );
   nor U49084 ( n47915,n47916,n47917 );
   nor U49085 ( n47917,n45579,n47465 );
   and U49086 ( n47916,n47504,n47918 );
   nor U49087 ( n47914,n47919,n47920 );
   nand U49088 ( n47920,n47921,n47922 );
   nand U49089 ( n47922,p1_instaddrpointer_reg_20_,n47923 );
   nand U49090 ( n47923,n47924,n47905 );
   and U49091 ( n47905,n47925,n47926 );
   nand U49092 ( n47926,n47499,n47927 );
   nor U49093 ( n47925,n47514,n47928 );
   nor U49094 ( n47928,n47929,n47520 );
   nor U49095 ( n47924,n47930,n47931 );
   nor U49096 ( n47931,p1_instaddrpointer_reg_19_,n47490 );
   nor U49097 ( n47930,n47932,n28253 );
   nand U49098 ( n47921,n47933,n47934 );
   nand U49099 ( n47933,n47935,n47936 );
   nand U49100 ( n47936,p1_instaddrpointer_reg_19_,n47912 );
   nand U49101 ( n47912,n47937,n47938 );
   nand U49102 ( n47938,n47929,n47512 );
   not U49103 ( n47929,n47939 );
   or U49104 ( n47937,n47927,n47613 );
   nand U49105 ( n47935,n47932,n28338 );
   nor U49106 ( n47919,n28294,n47940 );
   nor U49107 ( n47942,n47943,n47944 );
   nor U49108 ( n47944,n45574,n28113 );
   and U49109 ( n47943,n47504,n47945 );
   nor U49110 ( n47941,n47946,n47947 );
   nand U49111 ( n47947,n47948,n47949 );
   nand U49112 ( n47949,p1_instaddrpointer_reg_21_,n47950 );
   nand U49113 ( n47950,n47951,n47952 );
   nand U49114 ( n47952,n28338,n47953 );
   nand U49115 ( n47948,n47954,n47955 );
   nand U49116 ( n47954,n47956,n47957 );
   or U49117 ( n47957,n47953,n28253 );
   not U49118 ( n47956,n47958 );
   nor U49119 ( n47946,n28293,n47959 );
   nor U49120 ( n47961,n47962,n47963 );
   nor U49121 ( n47963,n45569,n28114 );
   and U49122 ( n47962,n47504,n47964 );
   nor U49123 ( n47960,n47965,n47966 );
   nand U49124 ( n47966,n47967,n47968 );
   nand U49125 ( n47968,p1_instaddrpointer_reg_22_,n47969 );
   nand U49126 ( n47969,n47970,n47951 );
   and U49127 ( n47951,n47971,n47972 );
   nand U49128 ( n47972,n47499,n47973 );
   nor U49129 ( n47971,n28232,n47974 );
   nor U49130 ( n47974,n47975,n47520 );
   nor U49131 ( n47970,n47976,n47977 );
   nor U49132 ( n47977,p1_instaddrpointer_reg_21_,n47490 );
   nor U49133 ( n47976,n47978,n28253 );
   nand U49134 ( n47967,n47979,n47980 );
   nand U49135 ( n47979,n47981,n47982 );
   nand U49136 ( n47982,p1_instaddrpointer_reg_21_,n47958 );
   nand U49137 ( n47958,n47983,n47984 );
   nand U49138 ( n47984,n47975,n47512 );
   not U49139 ( n47975,n47985 );
   or U49140 ( n47983,n47973,n47613 );
   nand U49141 ( n47981,n47978,n28338 );
   nor U49142 ( n47965,n28295,n47986 );
   nor U49143 ( n47988,n47989,n47990 );
   nor U49144 ( n47990,n45564,n47465 );
   nor U49145 ( n47989,n47466,n47991 );
   nor U49146 ( n47987,n47992,n47993 );
   nand U49147 ( n47993,n47994,n47995 );
   nand U49148 ( n47995,p1_instaddrpointer_reg_23_,n47996 );
   nand U49149 ( n47996,n47997,n47998 );
   nand U49150 ( n47998,n47519,n47999 );
   nand U49151 ( n47994,n48000,n48001 );
   nand U49152 ( n48000,n48002,n48003 );
   or U49153 ( n48003,n47999,n47474 );
   not U49154 ( n48002,n48004 );
   nor U49155 ( n47992,n28295,n48005 );
   nor U49156 ( n48007,n48008,n48009 );
   nor U49157 ( n48009,n45559,n28113 );
   and U49158 ( n48008,n28213,n48010 );
   nor U49159 ( n48006,n48011,n48012 );
   nand U49160 ( n48012,n48013,n48014 );
   nand U49161 ( n48014,p1_instaddrpointer_reg_24_,n48015 );
   nand U49162 ( n48015,n48016,n47997 );
   and U49163 ( n47997,n48017,n48018 );
   nand U49164 ( n48018,n47499,n48019 );
   nor U49165 ( n48017,n28232,n48020 );
   nor U49166 ( n48020,n48021,n28205 );
   nor U49167 ( n48016,n48022,n48023 );
   nor U49168 ( n48023,p1_instaddrpointer_reg_23_,n47490 );
   nor U49169 ( n48022,n48024,n47474 );
   nand U49170 ( n48013,n48025,n48026 );
   nand U49171 ( n48025,n48027,n48028 );
   nand U49172 ( n48028,p1_instaddrpointer_reg_23_,n48004 );
   nand U49173 ( n48004,n48029,n48030 );
   nand U49174 ( n48030,n48021,n47512 );
   not U49175 ( n48021,n48031 );
   or U49176 ( n48029,n48019,n47613 );
   nand U49177 ( n48027,n48024,n28338 );
   nor U49178 ( n48011,n28294,n48032 );
   nor U49179 ( n48034,n48035,n48036 );
   nor U49180 ( n48036,n45554,n28114 );
   and U49181 ( n48035,n47504,n48037 );
   nor U49182 ( n48033,n48038,n48039 );
   nand U49183 ( n48039,n48040,n48041 );
   nand U49184 ( n48041,p1_instaddrpointer_reg_25_,n48042 );
   nand U49185 ( n48042,n48043,n48044 );
   nand U49186 ( n48044,n47519,n48045 );
   nand U49187 ( n48040,n48046,n48047 );
   nand U49188 ( n48046,n48048,n48049 );
   or U49189 ( n48049,n48045,n28253 );
   not U49190 ( n48048,n48050 );
   nor U49191 ( n48038,n28294,n48051 );
   nor U49192 ( n48053,n48054,n48055 );
   nor U49193 ( n48055,n45549,n47465 );
   and U49194 ( n48054,n47504,n48056 );
   nor U49195 ( n48052,n48057,n48058 );
   nand U49196 ( n48058,n48059,n48060 );
   nand U49197 ( n48060,p1_instaddrpointer_reg_26_,n48061 );
   nand U49198 ( n48061,n48062,n48043 );
   and U49199 ( n48043,n48063,n48064 );
   nand U49200 ( n48064,n47499,n48065 );
   nor U49201 ( n48063,n28232,n48066 );
   nor U49202 ( n48066,n48067,n47520 );
   nor U49203 ( n48067,n48031,n48068 );
   nor U49204 ( n48062,n48069,n48070 );
   nor U49205 ( n48070,p1_instaddrpointer_reg_25_,n47490 );
   nor U49206 ( n48069,n48071,n28253 );
   nand U49207 ( n48059,n48072,n48073 );
   nand U49208 ( n48072,n48074,n48075 );
   nand U49209 ( n48075,p1_instaddrpointer_reg_25_,n48050 );
   nand U49210 ( n48050,n48076,n48077 );
   nand U49211 ( n48077,n48078,n48079 );
   nor U49212 ( n48078,n47520,n48031 );
   nand U49213 ( n48076,n48080,n47499 );
   nand U49214 ( n48074,n48071,n28338 );
   nor U49215 ( n48057,n28296,n48081 );
   nor U49216 ( n48083,n48084,n48085 );
   nor U49217 ( n48085,n45544,n28113 );
   nor U49218 ( n48084,n47466,n48086 );
   nor U49219 ( n48082,n48087,n48088 );
   nand U49220 ( n48088,n48089,n48090 );
   nand U49221 ( n48090,p1_instaddrpointer_reg_27_,n48091 );
   nand U49222 ( n48091,n48092,n48093 );
   nand U49223 ( n48093,n47519,n48094 );
   nand U49224 ( n48089,n48095,n48096 );
   nand U49225 ( n48095,n48097,n48098 );
   or U49226 ( n48098,n48094,n47474 );
   not U49227 ( n48097,n48099 );
   nor U49228 ( n48087,n28296,n48100 );
   nor U49229 ( n48102,n48103,n48104 );
   nor U49230 ( n48104,n45539,n28114 );
   and U49231 ( n48103,n28213,n48105 );
   nor U49232 ( n48101,n48106,n48107 );
   nand U49233 ( n48107,n48108,n48109 );
   nand U49234 ( n48109,p1_instaddrpointer_reg_28_,n48110 );
   nand U49235 ( n48110,n48111,n48092 );
   and U49236 ( n48092,n48112,n48113 );
   nand U49237 ( n48113,n47499,n48114 );
   nor U49238 ( n48112,n28232,n48115 );
   nor U49239 ( n48115,n48116,n47520 );
   nor U49240 ( n48111,n48117,n48118 );
   nor U49241 ( n48118,p1_instaddrpointer_reg_27_,n28238 );
   nor U49242 ( n48117,n48119,n47474 );
   nand U49243 ( n48108,n48120,n48121 );
   nand U49244 ( n48120,n48122,n48123 );
   nand U49245 ( n48123,p1_instaddrpointer_reg_27_,n48099 );
   nand U49246 ( n48122,n48119,n28338 );
   nor U49247 ( n48106,n28293,n48124 );
   nor U49248 ( n48126,n48127,n48128 );
   nor U49249 ( n48128,n45534,n47465 );
   nor U49250 ( n48127,n47466,n48129 );
   nor U49251 ( n48125,n48130,n48131 );
   nand U49252 ( n48131,n48132,n48133 );
   nand U49253 ( n48133,n48134,n48135 );
   or U49254 ( n48132,n48135,n48136 );
   not U49255 ( n48135,p1_instaddrpointer_reg_29_ );
   nor U49256 ( n48130,n28293,n48137 );
   nor U49257 ( n48139,n48140,n48141 );
   nor U49258 ( n48141,n45529,n28113 );
   and U49259 ( n48140,n47504,n48142 );
   nor U49260 ( n48138,n48143,n48144 );
   nand U49261 ( n48144,n48145,n48146 );
   or U49262 ( n48146,n48147,p1_instaddrpointer_reg_30_ );
   or U49263 ( n48145,n48148,n48149 );
   nor U49264 ( n48143,n28295,n48150 );
   nor U49265 ( n48152,n48153,n48154 );
   nor U49266 ( n48154,n45527,n28114 );
   nand U49267 ( n47465,n28374,n47473 );
   nor U49268 ( n48153,n28305,n48155 );
   not U49269 ( n47466,n47504 );
   nand U49270 ( n47504,n48156,n48157 );
   nand U49271 ( n48157,n48158,n47287 );
   nand U49272 ( n48156,n48159,n48160 );
   nand U49273 ( n48160,n48161,n48162 );
   nor U49274 ( n48162,n45864,n47457 );
   not U49275 ( n45864,n47429 );
   nor U49276 ( n48161,n47415,n48163 );
   nor U49277 ( n48163,n45879,n48164 );
   nand U49278 ( n48164,n48165,n47446 );
   nand U49279 ( n48165,n48166,n48167 );
   nand U49280 ( n48167,n45329,n47351 );
   nand U49281 ( n48166,n45358,n47303 );
   not U49282 ( n47415,n45872 );
   nand U49283 ( n45872,n48168,n45853 );
   nor U49284 ( n48168,n45877,n48169 );
   nor U49285 ( n48151,n48170,n48171 );
   nand U49286 ( n48171,n48172,n48173 );
   nand U49287 ( n48173,p1_instaddrpointer_reg_31_,n48174 );
   nand U49288 ( n48174,n48148,n48175 );
   nand U49289 ( n48175,n48176,n48149 );
   nand U49290 ( n48176,n28238,n47474 );
   nand U49291 ( n48148,n48177,n48178 );
   nand U49292 ( n48178,n48179,n28238 );
   nor U49293 ( n47490,n28300,n47512 );
   nor U49294 ( n48179,n47519,n48180 );
   nand U49295 ( n48177,n48136,p1_instaddrpointer_reg_29_ );
   nor U49296 ( n48136,n48180,n48181 );
   and U49297 ( n48181,n47519,n48182 );
   nand U49298 ( n48182,n48119,p1_instaddrpointer_reg_28_ );
   not U49299 ( n47519,n47474 );
   nand U49300 ( n48180,n48183,n48184 );
   nand U49301 ( n48184,n47499,n48185 );
   nand U49302 ( n48185,n48186,n48187 );
   nor U49303 ( n48183,n28232,n48188 );
   nor U49304 ( n48188,n48189,n28205 );
   and U49305 ( n48189,n48116,n48186 );
   nand U49306 ( n48172,n48190,n45480 );
   nor U49307 ( n48190,n48149,n48147 );
   nand U49308 ( n48147,p1_instaddrpointer_reg_29_,n48134 );
   nand U49309 ( n48134,n48191,n48192 );
   nand U49310 ( n48192,n48193,n48119 );
   nor U49311 ( n48119,n48094,n48096 );
   nand U49312 ( n48094,n48071,p1_instaddrpointer_reg_26_ );
   nor U49313 ( n48071,n48045,n48047 );
   nand U49314 ( n48045,n48024,p1_instaddrpointer_reg_24_ );
   nor U49315 ( n48024,n47999,n48001 );
   nand U49316 ( n47999,n47978,p1_instaddrpointer_reg_22_ );
   nor U49317 ( n47978,n47953,n47955 );
   nand U49318 ( n47953,n47932,p1_instaddrpointer_reg_20_ );
   nor U49319 ( n47932,n47907,n47909 );
   nand U49320 ( n47907,n47886,p1_instaddrpointer_reg_18_ );
   nor U49321 ( n47886,n47861,n47863 );
   nand U49322 ( n47861,n47840,p1_instaddrpointer_reg_16_ );
   nor U49323 ( n47840,n47815,n47817 );
   nand U49324 ( n47815,n47792,p1_instaddrpointer_reg_14_ );
   nor U49325 ( n47792,n47767,n47769 );
   nand U49326 ( n47767,n47746,p1_instaddrpointer_reg_12_ );
   nor U49327 ( n47746,n47721,n47723 );
   nand U49328 ( n47721,n47698,p1_instaddrpointer_reg_10_ );
   nor U49329 ( n47698,n47673,n47675 );
   nand U49330 ( n47673,n47652,p1_instaddrpointer_reg_8_ );
   nor U49331 ( n47652,n47627,n47629 );
   nand U49332 ( n47627,n47605,p1_instaddrpointer_reg_6_ );
   nor U49333 ( n47605,n47580,n47582 );
   nand U49334 ( n47580,n47560,p1_instaddrpointer_reg_4_ );
   and U49335 ( n47560,n48194,p1_instaddrpointer_reg_3_ );
   nor U49336 ( n48194,n45479,n47516 );
   nor U49337 ( n48193,n47474,n48121 );
   nand U49338 ( n47474,n48159,n45444 );
   nand U49339 ( n48191,n48186,n48099 );
   nand U49340 ( n48099,n48195,n48196 );
   nand U49341 ( n48196,n48116,n47512 );
   not U49342 ( n47512,n47520 );
   nand U49343 ( n47520,n48159,n48197 );
   nand U49344 ( n48197,n48198,n48199 );
   nor U49345 ( n48199,n47426,n48200 );
   nor U49346 ( n48198,n48201,n47430 );
   nand U49347 ( n47430,n48202,n48203 );
   nor U49348 ( n48203,n48204,n48205 );
   nand U49349 ( n48205,n48206,n48207 );
   nand U49350 ( n48204,n48208,n47443 );
   nand U49351 ( n47443,n48209,n27892 );
   not U49352 ( n48208,n48210 );
   nor U49353 ( n48202,n48211,n48212 );
   nand U49354 ( n48212,n48213,n48214 );
   nand U49355 ( n48214,n48215,n47334 );
   nand U49356 ( n48215,n48216,n48217 );
   nand U49357 ( n48217,n48218,n45878 );
   nand U49358 ( n48213,n47351,n45878 );
   nor U49359 ( n48211,n48219,n28405 );
   nor U49360 ( n48201,n47351,n47432 );
   not U49361 ( n47432,n48220 );
   and U49362 ( n48116,n48221,n48222 );
   nor U49363 ( n48222,n48031,n48047 );
   nand U49364 ( n48031,n48223,p1_instaddrpointer_reg_22_ );
   nor U49365 ( n48223,n47955,n47985 );
   nand U49366 ( n47985,n48224,p1_instaddrpointer_reg_20_ );
   nor U49367 ( n48224,n47909,n47939 );
   nand U49368 ( n47939,n48225,p1_instaddrpointer_reg_18_ );
   nor U49369 ( n48225,n47863,n47893 );
   nand U49370 ( n47893,n48226,p1_instaddrpointer_reg_16_ );
   nor U49371 ( n48226,n47817,n47847 );
   nand U49372 ( n47847,n48227,p1_instaddrpointer_reg_14_ );
   nor U49373 ( n48227,n47769,n47799 );
   nand U49374 ( n47799,n48228,p1_instaddrpointer_reg_12_ );
   nor U49375 ( n48228,n47723,n47753 );
   nand U49376 ( n47753,n48229,p1_instaddrpointer_reg_10_ );
   nor U49377 ( n48229,n47675,n47705 );
   nand U49378 ( n47705,n48230,p1_instaddrpointer_reg_8_ );
   nor U49379 ( n48230,n47629,n47659 );
   nand U49380 ( n47659,n48231,p1_instaddrpointer_reg_6_ );
   nor U49381 ( n48231,n47582,n47612 );
   nand U49382 ( n47612,n48232,p1_instaddrpointer_reg_4_ );
   nor U49383 ( n48232,n47536,n47502 );
   not U49384 ( n47502,n47557 );
   nor U49385 ( n47557,n47516,n47513 );
   not U49386 ( n47513,n45481 );
   not U49387 ( n47516,p1_instaddrpointer_reg_2_ );
   nor U49388 ( n48221,n48068,n48073 );
   nand U49389 ( n48195,n48187,n47499 );
   not U49390 ( n47499,n47613 );
   nand U49391 ( n47613,n48159,n47416 );
   not U49392 ( n48187,n48114 );
   nand U49393 ( n48114,n48233,p1_instaddrpointer_reg_26_ );
   nor U49394 ( n48233,n48047,n48065 );
   not U49395 ( n48065,n48080 );
   nor U49396 ( n48080,n48068,n48019 );
   nand U49397 ( n48019,n48234,p1_instaddrpointer_reg_22_ );
   nor U49398 ( n48234,n47955,n47973 );
   nand U49399 ( n47973,n48235,p1_instaddrpointer_reg_20_ );
   nor U49400 ( n48235,n47909,n47927 );
   nand U49401 ( n47927,n48236,p1_instaddrpointer_reg_18_ );
   nor U49402 ( n48236,n47863,n47881 );
   nand U49403 ( n47881,n48237,p1_instaddrpointer_reg_16_ );
   nor U49404 ( n48237,n47817,n47835 );
   nand U49405 ( n47835,n48238,p1_instaddrpointer_reg_14_ );
   nor U49406 ( n48238,n47769,n47787 );
   nand U49407 ( n47787,n48239,p1_instaddrpointer_reg_12_ );
   nor U49408 ( n48239,n47723,n47741 );
   nand U49409 ( n47741,n48240,p1_instaddrpointer_reg_10_ );
   nor U49410 ( n48240,n47675,n47693 );
   nand U49411 ( n47693,n48241,p1_instaddrpointer_reg_8_ );
   nor U49412 ( n48241,n47629,n47647 );
   nand U49413 ( n47647,n48242,p1_instaddrpointer_reg_6_ );
   nor U49414 ( n48242,n47582,n47600 );
   nand U49415 ( n47600,n48243,p1_instaddrpointer_reg_4_ );
   nor U49416 ( n48243,n47555,n47536 );
   nor U49417 ( n47555,p1_instaddrpointer_reg_2_,n45481 );
   nor U49418 ( n45481,n45479,n45448 );
   not U49419 ( n47629,p1_instaddrpointer_reg_7_ );
   not U49420 ( n47723,p1_instaddrpointer_reg_11_ );
   not U49421 ( n48068,n48079 );
   nor U49422 ( n48186,n48121,n48096 );
   nor U49423 ( n48170,n28295,n48244 );
   nand U49424 ( n48246,n48159,n45797 );
   nor U49425 ( n48159,n28374,n28232 );
   nand U49426 ( n48245,n48158,n48247 );
   and U49427 ( n48158,n48248,n48249 );
   nor U49428 ( n48248,n47514,n47428 );
   nand U49429 ( n47428,n48250,n47419 );
   not U49430 ( n47419,n48216 );
   nor U49431 ( n48250,n47334,n47271 );
   not U49432 ( n47514,n47473 );
   nand U49433 ( n47473,n48251,n48252 );
   nor U49434 ( n48252,n48253,n48254 );
   nor U49435 ( n48254,n48255,n45498 );
   not U49436 ( n45498,n45771 );
   nor U49437 ( n48255,n48256,n47447 );
   nand U49438 ( n47447,n48257,n48207 );
   nand U49439 ( n48207,n45358,n48258 );
   nand U49440 ( n48258,n48259,n48260 );
   nor U49441 ( n48257,n48261,n48262 );
   nor U49442 ( n48262,n47446,n48263 );
   nor U49443 ( n48263,n47351,n48264 );
   nor U49444 ( n48261,n48265,n45878 );
   nor U49445 ( n48265,n48266,n48267 );
   nand U49446 ( n48267,n48268,n47303 );
   nand U49447 ( n48268,n45876,n47420 );
   and U49448 ( n48256,n45853,n48269 );
   nor U49449 ( n48253,n48270,n48271 );
   nand U49450 ( n48271,n45759,n48260 );
   nor U49451 ( n48251,n48272,n48273 );
   nand U49452 ( n48273,n48274,n48275 );
   nand U49453 ( n48275,n48276,n45878 );
   nor U49454 ( n48276,n48277,n48278 );
   nand U49455 ( n48278,n45771,n48279 );
   nand U49456 ( n48277,n48280,n45346 );
   nand U49457 ( n48280,n45351,n47334 );
   nand U49458 ( n48274,n48281,n47446 );
   nor U49459 ( n48281,n48282,n48283 );
   nor U49460 ( n48282,n48284,n48285 );
   nand U49461 ( n48285,n48286,n47351 );
   nor U49462 ( n48284,n47433,n48287 );
   nand U49463 ( n48287,n48288,n45346 );
   nand U49464 ( n48288,n48289,n45351 );
   nor U49465 ( n48291,n48292,n48293 );
   nor U49466 ( n48293,n48294,n48295 );
   nor U49467 ( n48294,n48296,n48297 );
   nor U49468 ( n48292,n28268,n47467 );
   nand U49469 ( n47467,n48299,n48300 );
   or U49470 ( n48299,n48301,p1_instaddrpointer_reg_0_ );
   nor U49471 ( n48290,n48302,n48303 );
   nor U49472 ( n48303,n45373,n28120 );
   not U49473 ( n45373,p1_reip_reg_0_ );
   nor U49474 ( n48302,n48304,n48305 );
   nor U49475 ( n48307,n48308,n48309 );
   nor U49476 ( n48309,n48305,n48310 );
   nor U49477 ( n48308,n47483,n28268 );
   xor U49478 ( n47483,n48311,n48312 );
   xor U49479 ( n48312,n48300,p1_instaddrpointer_reg_1_ );
   nor U49480 ( n48306,n48313,n48314 );
   nand U49481 ( n48314,n48315,n48316 );
   nand U49482 ( n48316,n48296,n48317 );
   nand U49483 ( n48315,n48297,p1_phyaddrpointer_reg_1_ );
   nor U49484 ( n48313,n45674,n28120 );
   nor U49485 ( n48319,n48320,n48321 );
   nand U49486 ( n48321,n48322,n48323 );
   nand U49487 ( n48323,n48324,n47503 );
   xor U49488 ( n47503,n48325,n48326 );
   xor U49489 ( n48325,p1_instaddrpointer_reg_2_,n48327 );
   nand U49490 ( n48322,n48328,n48329 );
   nor U49491 ( n48320,n28289,n48331 );
   nor U49492 ( n48318,n48332,n48333 );
   nor U49493 ( n48333,n28396,n48335 );
   nor U49494 ( n48332,n45669,n28119 );
   nor U49495 ( n48337,n48338,n48339 );
   nand U49496 ( n48339,n48340,n48341 );
   or U49497 ( n48341,n48298,n47526 );
   xor U49498 ( n47526,n48342,n48343 );
   xor U49499 ( n48342,n48344,n47536 );
   not U49500 ( n47536,p1_instaddrpointer_reg_3_ );
   nand U49501 ( n48340,n48345,n28344 );
   and U49502 ( n48338,n48346,n48296 );
   nor U49503 ( n48336,n48347,n48348 );
   nor U49504 ( n48348,n28395,n48349 );
   nor U49505 ( n48347,n45664,n28118 );
   nor U49506 ( n48351,n48352,n48353 );
   nand U49507 ( n48353,n48354,n48355 );
   or U49508 ( n48355,n48298,n47546 );
   xor U49509 ( n47546,n48356,n48357 );
   xor U49510 ( n48356,n48358,n47562 );
   not U49511 ( n47562,p1_instaddrpointer_reg_4_ );
   nand U49512 ( n48354,n48359,n28344 );
   nor U49513 ( n48352,n48330,n48360 );
   nor U49514 ( n48350,n48361,n48362 );
   nor U49515 ( n48362,n28395,n48363 );
   nor U49516 ( n48361,n45659,n28120 );
   nor U49517 ( n48365,n48366,n48367 );
   nand U49518 ( n48367,n48368,n48369 );
   or U49519 ( n48369,n48298,n47572 );
   xor U49520 ( n47572,n48370,n48371 );
   xor U49521 ( n48370,n48372,n47582 );
   nand U49522 ( n48368,n48373,n28344 );
   and U49523 ( n48366,n48374,n48296 );
   nor U49524 ( n48364,n48375,n48376 );
   nor U49525 ( n48376,n48334,n48377 );
   nor U49526 ( n48375,n45654,n28119 );
   nor U49527 ( n48379,n48380,n48381 );
   nand U49528 ( n48381,n48382,n48383 );
   or U49529 ( n48383,n48298,n47591 );
   xor U49530 ( n47591,n48384,n48385 );
   xor U49531 ( n48384,n48386,n47607 );
   nand U49532 ( n48382,n48328,n48387 );
   nor U49533 ( n48380,n28290,n48388 );
   nor U49534 ( n48378,n48389,n48390 );
   nor U49535 ( n48390,n28395,n48391 );
   nor U49536 ( n48389,n45649,n28118 );
   nor U49537 ( n48393,n48394,n48395 );
   nand U49538 ( n48395,n48396,n48397 );
   or U49539 ( n48397,n48298,n47619 );
   nand U49540 ( n47619,n48398,n48399 );
   nand U49541 ( n48399,n48400,n48401 );
   nand U49542 ( n48400,n48402,n48403 );
   nand U49543 ( n48398,n48404,n48405 );
   xor U49544 ( n48404,n48406,p1_instaddrpointer_reg_7_ );
   nand U49545 ( n48396,n48407,n28344 );
   and U49546 ( n48394,n48408,n48296 );
   nor U49547 ( n48392,n48409,n48410 );
   nor U49548 ( n48410,n28396,n48411 );
   nor U49549 ( n48409,n45644,n28120 );
   nor U49550 ( n48413,n48414,n48415 );
   nand U49551 ( n48415,n48416,n48417 );
   nand U49552 ( n48417,n48324,n47638 );
   xor U49553 ( n47638,n48418,n48419 );
   nand U49554 ( n48419,n48402,n48420 );
   nand U49555 ( n48420,n48401,n48403 );
   not U49556 ( n48402,n48421 );
   xor U49557 ( n48418,n48422,p1_instaddrpointer_reg_8_ );
   nand U49558 ( n48416,n48328,n48423 );
   nor U49559 ( n48414,n28289,n48424 );
   nor U49560 ( n48412,n48425,n48426 );
   nor U49561 ( n48426,n48334,n48427 );
   nor U49562 ( n48425,n45639,n28119 );
   nor U49563 ( n48429,n48430,n48431 );
   nand U49564 ( n48431,n48432,n48433 );
   nand U49565 ( n48433,n48324,n47665 );
   nand U49566 ( n47665,n48434,n48435 );
   nand U49567 ( n48435,n48436,n48437 );
   nand U49568 ( n48436,n48438,n48439 );
   nand U49569 ( n48434,n48440,n48439 );
   nand U49570 ( n48432,n48328,n48441 );
   and U49571 ( n48430,n48442,n48296 );
   nor U49572 ( n48428,n48443,n48444 );
   nor U49573 ( n48444,n28395,n48445 );
   nor U49574 ( n48443,n45634,n28118 );
   nor U49575 ( n48447,n48448,n48449 );
   nand U49576 ( n48449,n48450,n48451 );
   nand U49577 ( n48451,n48324,n47684 );
   xor U49578 ( n47684,n48452,n48453 );
   nor U49579 ( n48452,n48454,n48455 );
   nand U49580 ( n48450,n48328,n48456 );
   nor U49581 ( n48448,n28290,n48457 );
   nor U49582 ( n48446,n48458,n48459 );
   nor U49583 ( n48459,n28396,n48460 );
   nor U49584 ( n48458,n45629,n28118 );
   nor U49585 ( n48462,n48463,n48464 );
   nand U49586 ( n48464,n48465,n48466 );
   nand U49587 ( n48466,n48467,n27890 );
   nor U49588 ( n48467,n48468,n47711 );
   nor U49589 ( n47711,n48469,n48470 );
   not U49590 ( n48468,n47713 );
   nand U49591 ( n47713,n48471,n48472 );
   nor U49592 ( n48471,n48455,n48473 );
   nor U49593 ( n48473,n48474,n48470 );
   not U49594 ( n48470,n48475 );
   not U49595 ( n48455,n48476 );
   nand U49596 ( n48465,n48328,n48477 );
   and U49597 ( n48463,n48478,n48296 );
   nor U49598 ( n48461,n48479,n48480 );
   nor U49599 ( n48480,n48334,n48481 );
   nor U49600 ( n48479,n45624,n28119 );
   nor U49601 ( n48483,n48484,n48485 );
   nand U49602 ( n48485,n48486,n48487 );
   nand U49603 ( n48487,n48324,n47732 );
   xor U49604 ( n47732,n48488,n48489 );
   and U49605 ( n48488,n48490,n48491 );
   nand U49606 ( n48486,n48328,n48492 );
   nor U49607 ( n48484,n48330,n48493 );
   nor U49608 ( n48482,n48494,n48495 );
   nor U49609 ( n48495,n28395,n48496 );
   nor U49610 ( n48494,n45619,n28118 );
   nor U49611 ( n48498,n48499,n48500 );
   nand U49612 ( n48500,n48501,n48502 );
   nand U49613 ( n48502,n48324,n47759 );
   xor U49614 ( n47759,n48503,n48504 );
   and U49615 ( n48503,n48505,n48506 );
   nand U49616 ( n48501,n48328,n48507 );
   and U49617 ( n48499,n48508,n48296 );
   not U49618 ( n48296,n48330 );
   nor U49619 ( n48497,n48509,n48510 );
   nor U49620 ( n48510,n28396,n48511 );
   nor U49621 ( n48509,n45614,n28119 );
   nor U49622 ( n48513,n48514,n48515 );
   nand U49623 ( n48515,n48516,n48517 );
   or U49624 ( n48517,n48298,n47778 );
   xor U49625 ( n47778,n48518,n48519 );
   nor U49626 ( n48518,n48520,n48521 );
   nand U49627 ( n48516,n28344,n48522 );
   nor U49628 ( n48514,n28289,n48523 );
   nor U49629 ( n48512,n48524,n48525 );
   nor U49630 ( n48525,n28395,n48526 );
   nor U49631 ( n48524,n45609,n28120 );
   nor U49632 ( n48528,n48529,n48530 );
   nand U49633 ( n48530,n48531,n48532 );
   nand U49634 ( n48532,n48533,n27890 );
   nor U49635 ( n48533,n48534,n47805 );
   and U49636 ( n47805,n48535,n48536 );
   xor U49637 ( n48536,n48537,p1_instaddrpointer_reg_15_ );
   nor U49638 ( n48535,n48520,n48538 );
   nor U49639 ( n48538,n48519,n48521 );
   not U49640 ( n48519,n48539 );
   not U49641 ( n48534,n47807 );
   nand U49642 ( n47807,n48540,n48541 );
   nor U49643 ( n48540,n48542,n48543 );
   nor U49644 ( n48543,n48520,n48539 );
   nand U49645 ( n48539,n48544,n48505 );
   not U49646 ( n48505,n48545 );
   nand U49647 ( n48544,n48506,n48504 );
   nand U49648 ( n48504,n48490,n48546 );
   nand U49649 ( n48531,n48328,n48547 );
   nor U49650 ( n48529,n28289,n48548 );
   nor U49651 ( n48527,n48549,n48550 );
   nor U49652 ( n48550,n48334,n48551 );
   nor U49653 ( n48549,n45604,n28118 );
   nor U49654 ( n48553,n48554,n48555 );
   nand U49655 ( n48555,n48556,n48557 );
   nand U49656 ( n48557,n48324,n47826 );
   nand U49657 ( n47826,n48558,n48559 );
   nand U49658 ( n48559,n48560,n48561 );
   nor U49659 ( n48558,n48562,n48563 );
   nor U49660 ( n48563,n47842,n48564 );
   xor U49661 ( n48564,n48565,n48561 );
   not U49662 ( n47842,p1_instaddrpointer_reg_16_ );
   nor U49663 ( n48562,p1_instaddrpointer_reg_16_,n48566 );
   nand U49664 ( n48566,n48567,n48565 );
   nand U49665 ( n48556,n48568,n28344 );
   nor U49666 ( n48554,n28289,n48569 );
   nor U49667 ( n48552,n48570,n48571 );
   nor U49668 ( n48571,n28395,n48572 );
   nor U49669 ( n48570,n45599,n28119 );
   nor U49670 ( n48574,n48575,n48576 );
   nand U49671 ( n48576,n48577,n48578 );
   or U49672 ( n48578,n28268,n47853 );
   xor U49673 ( n47853,n48579,n48580 );
   or U49674 ( n48580,n48581,n48582 );
   nand U49675 ( n48577,n48328,n48583 );
   nor U49676 ( n48575,n48584,n28290 );
   nor U49677 ( n48573,n48585,n48586 );
   nor U49678 ( n48586,n28396,n48587 );
   nor U49679 ( n48585,n45594,n28120 );
   nor U49680 ( n48589,n48590,n48591 );
   nand U49681 ( n48591,n48592,n48593 );
   or U49682 ( n48593,n48298,n47872 );
   xor U49683 ( n47872,n48594,n48595 );
   or U49684 ( n48595,n48596,n48597 );
   nor U49685 ( n48594,n48582,n48598 );
   nor U49686 ( n48598,n48579,n48581 );
   nor U49687 ( n48579,n48560,n48599 );
   and U49688 ( n48599,n48567,n48600 );
   nand U49689 ( n48600,p1_instaddrpointer_reg_16_,n48565 );
   nand U49690 ( n48592,n48601,n28344 );
   nor U49691 ( n48590,n28289,n48602 );
   nor U49692 ( n48588,n48603,n48604 );
   nor U49693 ( n48604,n48334,n48605 );
   nor U49694 ( n48603,n45589,n28118 );
   nor U49695 ( n48607,n48608,n48609 );
   nand U49696 ( n48609,n48610,n48611 );
   nand U49697 ( n48611,n48324,n47899 );
   xor U49698 ( n47899,n48612,n48613 );
   and U49699 ( n48612,n48614,n48615 );
   nand U49700 ( n48610,n48328,n48616 );
   nor U49701 ( n48608,n28290,n48617 );
   nor U49702 ( n48606,n48618,n48619 );
   nor U49703 ( n48619,n48334,n48620 );
   nor U49704 ( n48618,n45584,n28119 );
   nor U49705 ( n48622,n48623,n48624 );
   nand U49706 ( n48624,n48625,n48626 );
   nand U49707 ( n48626,n48324,n47918 );
   xor U49708 ( n47918,n48627,n48628 );
   and U49709 ( n48627,n48629,n48630 );
   nand U49710 ( n48625,n48631,n28344 );
   nor U49711 ( n48623,n28290,n48632 );
   nor U49712 ( n48621,n48633,n48634 );
   nor U49713 ( n48634,n28396,n48635 );
   nor U49714 ( n48633,n45579,n28120 );
   nor U49715 ( n48637,n48638,n48639 );
   nand U49716 ( n48639,n48640,n48641 );
   nand U49717 ( n48641,n48324,n47945 );
   xor U49718 ( n47945,n48642,n48643 );
   nand U49719 ( n48643,n48629,n48644 );
   nand U49720 ( n48644,n48630,n48628 );
   nand U49721 ( n48628,n48614,n48645 );
   nand U49722 ( n48645,n48615,n48613 );
   not U49723 ( n48615,n48646 );
   nand U49724 ( n48614,p1_instaddrpointer_reg_19_,n28341 );
   nand U49725 ( n48629,p1_instaddrpointer_reg_20_,n28341 );
   nor U49726 ( n48642,n48648,n48649 );
   nor U49727 ( n48648,n48650,n47955 );
   not U49728 ( n47955,p1_instaddrpointer_reg_21_ );
   nand U49729 ( n48640,n48651,n28344 );
   nor U49730 ( n48638,n48652,n28289 );
   nor U49731 ( n48636,n48653,n48654 );
   nor U49732 ( n48654,n28395,n48655 );
   nor U49733 ( n48653,n45574,n28119 );
   nor U49734 ( n48657,n48658,n48659 );
   nand U49735 ( n48659,n48660,n48661 );
   nand U49736 ( n48661,n48324,n47964 );
   xor U49737 ( n47964,n48662,n48663 );
   nand U49738 ( n48663,n48664,n48665 );
   nand U49739 ( n48665,n48666,n48613 );
   nand U49740 ( n48613,n48667,n48668 );
   nor U49741 ( n48662,n48669,n48670 );
   nand U49742 ( n48660,n28344,n48671 );
   nor U49743 ( n48658,n48330,n48672 );
   nor U49744 ( n48656,n48673,n48674 );
   nor U49745 ( n48674,n48334,n48675 );
   nor U49746 ( n48673,n45569,n28118 );
   nor U49747 ( n48677,n48678,n48679 );
   nand U49748 ( n48679,n48680,n48681 );
   or U49749 ( n48681,n28268,n47991 );
   nand U49750 ( n47991,n48682,n48683 );
   or U49751 ( n48683,n48684,n48685 );
   nor U49752 ( n48682,n48686,n48687 );
   nor U49753 ( n48687,p1_instaddrpointer_reg_23_,n48688 );
   xor U49754 ( n48688,n48647,n48685 );
   nor U49755 ( n48686,n48001,n48689 );
   nand U49756 ( n48689,n48685,n28265 );
   nand U49757 ( n48680,n28344,n48690 );
   nor U49758 ( n48678,n28289,n48691 );
   nor U49759 ( n48676,n48692,n48693 );
   nor U49760 ( n48693,n28396,n48694 );
   nor U49761 ( n48692,n45564,n28120 );
   nor U49762 ( n48696,n48697,n48698 );
   nand U49763 ( n48698,n48699,n48700 );
   nand U49764 ( n48700,n48324,n48010 );
   xor U49765 ( n48010,n48701,n48702 );
   nand U49766 ( n48702,n48703,n48684 );
   xor U49767 ( n48701,n48026,n48650 );
   nand U49768 ( n48699,n48704,n28344 );
   nor U49769 ( n48697,n28290,n48705 );
   nor U49770 ( n48695,n48706,n48707 );
   nor U49771 ( n48707,n48334,n48708 );
   nor U49772 ( n48706,n45559,n28119 );
   nor U49773 ( n48710,n48711,n48712 );
   nand U49774 ( n48712,n48713,n48714 );
   nand U49775 ( n48714,n48324,n48037 );
   xor U49776 ( n48037,n48715,n48716 );
   or U49777 ( n48716,n48717,n48718 );
   nor U49778 ( n48715,n48719,n48720 );
   nor U49779 ( n48719,n48721,n48703 );
   nand U49780 ( n48703,n48722,n48685 );
   nand U49781 ( n48722,n48001,n28265 );
   nor U49782 ( n48721,n48647,p1_instaddrpointer_reg_24_ );
   nand U49783 ( n48713,n48723,n28344 );
   nor U49784 ( n48711,n48724,n28290 );
   nor U49785 ( n48709,n48725,n48726 );
   nor U49786 ( n48726,n28395,n48727 );
   nor U49787 ( n48725,n45554,n28118 );
   nor U49788 ( n48729,n48730,n48731 );
   nand U49789 ( n48731,n48732,n48733 );
   nand U49790 ( n48733,n48324,n48056 );
   xor U49791 ( n48056,n48734,n48735 );
   nor U49792 ( n48734,n48736,n48737 );
   nand U49793 ( n48732,n48328,n48738 );
   nor U49794 ( n48730,n48330,n48739 );
   nor U49795 ( n48728,n48740,n48741 );
   nor U49796 ( n48741,n48334,n48742 );
   nor U49797 ( n48740,n45549,n28120 );
   nor U49798 ( n48744,n48745,n48746 );
   nand U49799 ( n48746,n48747,n48748 );
   or U49800 ( n48748,n48298,n48086 );
   xor U49801 ( n48086,n48749,n48750 );
   nand U49802 ( n48750,n48751,n48752 );
   nand U49803 ( n48752,n28265,n48096 );
   not U49804 ( n48751,n48753 );
   nor U49805 ( n48749,n48754,n48737 );
   nor U49806 ( n48754,n48736,n48735 );
   nand U49807 ( n48735,n48755,n48756 );
   nor U49808 ( n48755,n48718,n48757 );
   nor U49809 ( n48757,n48758,n48759 );
   nand U49810 ( n48759,n48685,n48760 );
   nor U49811 ( n48718,n48047,n48650 );
   nor U49812 ( n48736,n48650,n48073 );
   nand U49813 ( n48747,n28344,n48761 );
   nor U49814 ( n48745,n48762,n48330 );
   nor U49815 ( n48743,n48763,n48764 );
   and U49816 ( n48764,n48297,p1_phyaddrpointer_reg_27_ );
   nor U49817 ( n48763,n45544,n28119 );
   nor U49818 ( n48766,n48767,n48768 );
   nand U49819 ( n48768,n48769,n48770 );
   nand U49820 ( n48770,n48324,n48105 );
   xor U49821 ( n48105,n48771,n48772 );
   nand U49822 ( n48772,n48773,n48774 );
   nand U49823 ( n48774,n48775,n48685 );
   nand U49824 ( n48685,n48776,n48777 );
   nor U49825 ( n48776,n48778,n48779 );
   nor U49826 ( n48779,n48667,n48780 );
   and U49827 ( n48667,n48781,n48782 );
   xor U49828 ( n48771,n48121,n48650 );
   nand U49829 ( n48769,n48328,n48783 );
   nor U49830 ( n48767,n28290,n48784 );
   nor U49831 ( n48765,n48785,n48786 );
   nor U49832 ( n48786,n28396,n48787 );
   nor U49833 ( n48785,n45539,n28118 );
   nor U49834 ( n48789,n48790,n48791 );
   nand U49835 ( n48791,n48792,n48793 );
   or U49836 ( n48793,n28268,n48129 );
   xor U49837 ( n48129,n48794,n48795 );
   nand U49838 ( n48795,n48796,n48797 );
   nand U49839 ( n48792,n48328,n48798 );
   nor U49840 ( n48790,n48330,n48799 );
   nor U49841 ( n48788,n48800,n48801 );
   nor U49842 ( n48801,n28395,n48802 );
   nor U49843 ( n48800,n45534,n28120 );
   nor U49844 ( n48804,n48805,n48806 );
   nand U49845 ( n48806,n48807,n48808 );
   nand U49846 ( n48808,n48324,n48142 );
   nand U49847 ( n48142,n48809,n48810 );
   nand U49848 ( n48810,n48811,n48812 );
   nor U49849 ( n48809,n48813,n48814 );
   nor U49850 ( n48814,n48149,n48815 );
   xor U49851 ( n48815,n48647,n48812 );
   not U49852 ( n48149,p1_instaddrpointer_reg_30_ );
   nor U49853 ( n48813,p1_instaddrpointer_reg_30_,n48816 );
   or U49854 ( n48816,n48812,n28265 );
   nand U49855 ( n48812,n48817,n48818 );
   nor U49856 ( n48818,n48819,n48820 );
   nand U49857 ( n48820,n48797,n48821 );
   not U49858 ( n48821,n48822 );
   nand U49859 ( n48797,p1_instaddrpointer_reg_29_,n28341 );
   and U49860 ( n48819,n48796,n48823 );
   nand U49861 ( n48807,n48328,n48824 );
   nor U49862 ( n48805,n48330,n48825 );
   nor U49863 ( n48803,n48826,n48827 );
   nor U49864 ( n48827,n48334,n48828 );
   nor U49865 ( n48826,n45529,n28119 );
   nor U49866 ( n48830,n48831,n48832 );
   nand U49867 ( n48832,n48833,n48834 );
   nand U49868 ( n48834,n48835,n28344 );
   not U49869 ( n48328,n48305 );
   nand U49870 ( n48305,n48836,p1_statebs16_reg );
   nor U49871 ( n48836,n48297,n45432 );
   or U49872 ( n48833,n28268,n48155 );
   nand U49873 ( n48155,n48837,n48838 );
   nand U49874 ( n48838,n48839,n48811 );
   nor U49875 ( n48837,n48840,n48841 );
   nor U49876 ( n48841,n48842,n48843 );
   nand U49877 ( n48843,n48817,n48844 );
   nor U49878 ( n48844,n48845,n48846 );
   nor U49879 ( n48846,n48847,n48848 );
   nor U49880 ( n48840,n48849,n48839 );
   not U49881 ( n48839,n48842 );
   xor U49882 ( n48842,n48647,p1_instaddrpointer_reg_31_ );
   nor U49883 ( n48849,n48850,n48845 );
   nor U49884 ( n48845,n48851,n48650 );
   nor U49885 ( n48851,p1_instaddrpointer_reg_30_,p1_instaddrpointer_reg_29_ );
   nor U49886 ( n48850,n48811,n48852 );
   nand U49887 ( n48852,n48794,n48796 );
   not U49888 ( n48796,n48848 );
   nor U49889 ( n48848,n28341,p1_instaddrpointer_reg_29_ );
   nand U49890 ( n48794,n48817,n48847 );
   nor U49891 ( n48847,n48822,n48823 );
   nor U49892 ( n48823,n48853,n48781 );
   nand U49893 ( n48781,n48854,n48855 );
   nor U49894 ( n48855,n48582,n48567 );
   not U49895 ( n48567,n48561 );
   nand U49896 ( n48561,n48856,n48857 );
   nand U49897 ( n48857,n48541,n48858 );
   nand U49898 ( n48858,n48859,n48860 );
   nand U49899 ( n48860,n48861,n48506 );
   not U49900 ( n48861,n48490 );
   nand U49901 ( n48490,n48862,p1_instaddrpointer_reg_12_ );
   nor U49902 ( n48862,n48863,n48864 );
   nor U49903 ( n48859,n48545,n48520 );
   nor U49904 ( n48520,n47794,n48865 );
   nor U49905 ( n48545,n47769,n48866 );
   nor U49906 ( n48856,n48867,n48542 );
   nor U49907 ( n48542,n47817,n48537 );
   nor U49908 ( n48867,n48546,n48868 );
   nand U49909 ( n48868,n48541,n48506 );
   nand U49910 ( n48506,n47769,n48866 );
   nand U49911 ( n48866,n48869,n48870 );
   not U49912 ( n47769,p1_instaddrpointer_reg_13_ );
   nor U49913 ( n48541,n48521,n48871 );
   and U49914 ( n48871,n48537,n47817 );
   not U49915 ( n47817,p1_instaddrpointer_reg_15_ );
   nand U49916 ( n48537,n48872,n48870 );
   nor U49917 ( n48872,n48873,n48874 );
   nor U49918 ( n48874,n48875,n48876 );
   and U49919 ( n48521,n47794,n48865 );
   nand U49920 ( n48865,n48877,n48870 );
   not U49921 ( n47794,p1_instaddrpointer_reg_14_ );
   nand U49922 ( n48546,n48491,n48489 );
   nand U49923 ( n48489,n48469,n48475 );
   nand U49924 ( n48475,p1_instaddrpointer_reg_11_,n48878 );
   or U49925 ( n48469,n48474,n48879 );
   and U49926 ( n48879,n48472,n48476 );
   nand U49927 ( n48476,p1_instaddrpointer_reg_10_,n48880 );
   nand U49928 ( n48472,n48453,n48881 );
   not U49929 ( n48881,n48454 );
   nor U49930 ( n48454,p1_instaddrpointer_reg_10_,n48880 );
   nor U49931 ( n48880,n48882,n48863 );
   nor U49932 ( n48453,n48440,n48883 );
   not U49933 ( n48883,n48439 );
   nand U49934 ( n48439,n47675,n48884 );
   nand U49935 ( n48884,n48885,n48870 );
   not U49936 ( n47675,p1_instaddrpointer_reg_9_ );
   nor U49937 ( n48440,n48437,n48886 );
   not U49938 ( n48886,n48438 );
   nand U49939 ( n48438,n48887,p1_instaddrpointer_reg_9_ );
   nor U49940 ( n48887,n48863,n48888 );
   nand U49941 ( n48437,n48889,n48890 );
   nand U49942 ( n48890,n48891,n48405 );
   not U49943 ( n48405,n48401 );
   nand U49944 ( n48401,n48892,n48893 );
   nand U49945 ( n48893,n48894,n47607 );
   not U49946 ( n47607,p1_instaddrpointer_reg_6_ );
   nand U49947 ( n48894,n48385,n48386 );
   or U49948 ( n48892,n48386,n48385 );
   and U49949 ( n48385,n48895,n48896 );
   nand U49950 ( n48896,n48897,n47582 );
   not U49951 ( n47582,p1_instaddrpointer_reg_5_ );
   nand U49952 ( n48897,n48372,n48371 );
   or U49953 ( n48895,n48371,n48372 );
   nand U49954 ( n48372,n48898,n48899 );
   nand U49955 ( n48899,n48900,n45358 );
   nor U49956 ( n48900,n48901,n48902 );
   nor U49957 ( n48902,n48903,n48904 );
   nand U49958 ( n48898,n48870,n48905 );
   nand U49959 ( n48371,n48906,n48907 );
   nand U49960 ( n48907,p1_instaddrpointer_reg_4_,n48908 );
   or U49961 ( n48908,n48357,n48358 );
   nand U49962 ( n48906,n48357,n48358 );
   nand U49963 ( n48358,n48909,n48910 );
   or U49964 ( n48910,n48911,n48912 );
   xor U49965 ( n48911,n48913,n48914 );
   nand U49966 ( n48914,n48915,n48916 );
   nand U49967 ( n48909,n48917,n48870 );
   nand U49968 ( n48357,n48918,n48919 );
   nand U49969 ( n48919,p1_instaddrpointer_reg_3_,n48920 );
   or U49970 ( n48920,n48343,n48344 );
   nand U49971 ( n48918,n48343,n48344 );
   nand U49972 ( n48344,n48921,n48922 );
   nand U49973 ( n48922,n45358,n48923 );
   xor U49974 ( n48923,n48916,n48915 );
   nand U49975 ( n48921,n45428,n48870 );
   nand U49976 ( n48343,n48924,n48925 );
   nand U49977 ( n48925,p1_instaddrpointer_reg_2_,n48926 );
   nand U49978 ( n48926,n48327,n48326 );
   or U49979 ( n48924,n48326,n48327 );
   and U49980 ( n48327,n48927,n48928 );
   nand U49981 ( n48928,n45358,n48929 );
   nand U49982 ( n48929,n48930,n48916 );
   nand U49983 ( n48930,n48931,n48932 );
   nor U49984 ( n48931,n48933,n48934 );
   nor U49985 ( n48927,n48935,n48936 );
   nor U49986 ( n48936,n46269,n48863 );
   nand U49987 ( n48326,n48937,n48938 );
   nand U49988 ( n48938,n48939,n45479 );
   nand U49989 ( n48939,n48940,n48311 );
   or U49990 ( n48937,n48311,n48940 );
   not U49991 ( n48940,n48300 );
   nand U49992 ( n48300,p1_instaddrpointer_reg_0_,n48301 );
   nand U49993 ( n48301,n48941,n48942 );
   nand U49994 ( n48942,n48933,n45358 );
   nor U49995 ( n48941,n48935,n48943 );
   nor U49996 ( n48943,n47130,n48863 );
   nor U49997 ( n48935,n47351,n45877 );
   nand U49998 ( n48311,n48944,n48945 );
   nor U49999 ( n48945,n45878,n48946 );
   nand U50000 ( n48946,n47303,n47271 );
   nor U50001 ( n48944,n48947,n48948 );
   nor U50002 ( n48948,n48863,n47373 );
   not U50003 ( n47373,n45401 );
   nor U50004 ( n48947,n48949,n48912 );
   xor U50005 ( n48949,n48950,n48934 );
   nand U50006 ( n48386,n48951,n48952 );
   nand U50007 ( n48952,n48953,n45358 );
   xor U50008 ( n48953,n48954,n48901 );
   not U50009 ( n48901,n48955 );
   nand U50010 ( n48951,n48956,n48870 );
   nor U50011 ( n48891,n48421,n48957 );
   nor U50012 ( n48957,p1_instaddrpointer_reg_8_,n48958 );
   nor U50013 ( n48421,n48406,p1_instaddrpointer_reg_7_ );
   nor U50014 ( n48889,n48959,n48960 );
   nor U50015 ( n48960,n48422,n48403 );
   nor U50016 ( n48959,n48961,n47654 );
   not U50017 ( n47654,p1_instaddrpointer_reg_8_ );
   and U50018 ( n48961,n48403,n48422 );
   not U50019 ( n48422,n48958 );
   nand U50020 ( n48958,n48962,n48963 );
   nand U50021 ( n48963,n48964,n48965 );
   nor U50022 ( n48965,n48966,n48967 );
   nor U50023 ( n48964,n48912,n48955 );
   nand U50024 ( n48962,n48870,n48968 );
   xor U50025 ( n48968,n48969,n48970 );
   nand U50026 ( n48403,p1_instaddrpointer_reg_7_,n48406 );
   nand U50027 ( n48406,n48971,n48972 );
   nand U50028 ( n48972,n48973,n48974 );
   nor U50029 ( n48973,n48863,n48975 );
   nand U50030 ( n48971,n48976,n45358 );
   xor U50031 ( n48976,n48977,n48978 );
   nor U50032 ( n48977,n48967,n48955 );
   nand U50033 ( n48955,n48903,n48904 );
   and U50034 ( n48903,n48979,n48913 );
   and U50035 ( n48979,n48915,n48916 );
   nand U50036 ( n48916,n48980,n48981 );
   nand U50037 ( n48981,n48982,n48950 );
   not U50038 ( n48967,n48954 );
   nor U50039 ( n48474,n48878,p1_instaddrpointer_reg_11_ );
   nor U50040 ( n48878,n48983,n48863 );
   nand U50041 ( n48491,n47748,n48984 );
   nand U50042 ( n48984,n48985,n48870 );
   not U50043 ( n47748,p1_instaddrpointer_reg_12_ );
   nor U50044 ( n48582,n48647,p1_instaddrpointer_reg_17_ );
   nor U50045 ( n48854,n48560,n48597 );
   nor U50046 ( n48597,p1_instaddrpointer_reg_18_,n28341 );
   nor U50047 ( n48560,n48565,p1_instaddrpointer_reg_16_ );
   or U50048 ( n48853,n48780,n48986 );
   nor U50049 ( n48822,n48987,n48986 );
   nand U50050 ( n48986,n48775,n48988 );
   nand U50051 ( n48988,n28265,n48121 );
   and U50052 ( n48775,n48989,n48990 );
   nor U50053 ( n48989,n48717,n48758 );
   nor U50054 ( n48758,n48647,n48079 );
   nor U50055 ( n48079,n48026,n48001 );
   not U50056 ( n48001,p1_instaddrpointer_reg_23_ );
   not U50057 ( n48026,p1_instaddrpointer_reg_24_ );
   not U50058 ( n48717,n48760 );
   nand U50059 ( n48760,n48650,n48047 );
   or U50060 ( n48987,n48782,n48780 );
   nand U50061 ( n48780,n48666,n48991 );
   not U50062 ( n48991,n48669 );
   nor U50063 ( n48669,p1_instaddrpointer_reg_22_,n28341 );
   and U50064 ( n48666,n48992,n48630 );
   nand U50065 ( n48630,n47934,n28265 );
   not U50066 ( n47934,p1_instaddrpointer_reg_20_ );
   nor U50067 ( n48992,n48649,n48646 );
   nor U50068 ( n48646,p1_instaddrpointer_reg_19_,n28341 );
   nor U50069 ( n48649,n28341,p1_instaddrpointer_reg_21_ );
   nor U50070 ( n48782,n48581,n48993 );
   and U50071 ( n48993,p1_instaddrpointer_reg_16_,n48565 );
   nand U50072 ( n48565,n28265,n48994 );
   nand U50073 ( n48994,n48995,n48873 );
   nor U50074 ( n48995,n48996,n48863 );
   nor U50075 ( n48581,n47863,n48650 );
   not U50076 ( n47863,p1_instaddrpointer_reg_17_ );
   nor U50077 ( n48817,n48997,n48998 );
   nand U50078 ( n48998,n48999,n48773 );
   nor U50079 ( n48773,n48753,n49000 );
   and U50080 ( n49000,n48990,n49001 );
   nand U50081 ( n49001,n48756,n49002 );
   nand U50082 ( n49002,n28341,n49003 );
   nand U50083 ( n49003,n48047,n48073 );
   not U50084 ( n48073,p1_instaddrpointer_reg_26_ );
   not U50085 ( n48047,p1_instaddrpointer_reg_25_ );
   not U50086 ( n48756,n48720 );
   nand U50087 ( n48720,n48684,n49004 );
   nand U50088 ( n49004,p1_instaddrpointer_reg_24_,n28341 );
   nand U50089 ( n48684,p1_instaddrpointer_reg_23_,n28341 );
   nor U50090 ( n48990,n48737,n49005 );
   nor U50091 ( n49005,n28341,p1_instaddrpointer_reg_27_ );
   nor U50092 ( n48737,n48647,p1_instaddrpointer_reg_26_ );
   nor U50093 ( n48753,n48096,n48650 );
   not U50094 ( n48096,p1_instaddrpointer_reg_27_ );
   nor U50095 ( n48999,n48778,n49006 );
   nor U50096 ( n49006,n48650,n48121 );
   not U50097 ( n48121,p1_instaddrpointer_reg_28_ );
   not U50098 ( n48778,n48664 );
   nand U50099 ( n48664,n28341,n49007 );
   nand U50100 ( n49007,n49008,n47909 );
   not U50101 ( n47909,p1_instaddrpointer_reg_19_ );
   nor U50102 ( n49008,p1_instaddrpointer_reg_21_,p1_instaddrpointer_reg_20_ );
   not U50103 ( n48997,n48777 );
   nor U50104 ( n48777,n48670,n48596 );
   not U50105 ( n48596,n48668 );
   nand U50106 ( n48668,p1_instaddrpointer_reg_18_,n28341 );
   nor U50107 ( n48670,n47980,n48650 );
   not U50108 ( n47980,p1_instaddrpointer_reg_22_ );
   nor U50109 ( n48811,p1_instaddrpointer_reg_30_,n28341 );
   not U50110 ( n48647,n48650 );
   nand U50111 ( n48650,n49009,n48870 );
   not U50112 ( n48298,n48324 );
   nor U50113 ( n48324,n28095,n48297 );
   nor U50114 ( n48831,n49010,n28289 );
   nand U50115 ( n48330,n49011,n49012 );
   nor U50116 ( n49012,n49013,n45352 );
   nor U50117 ( n49011,p1_state2_reg_0_,n48297 );
   not U50118 ( n48297,n28396 );
   nor U50119 ( n48829,n49014,n49015 );
   nor U50120 ( n49015,n28396,n49016 );
   nor U50121 ( n49014,n45527,n28118 );
   nand U50122 ( n48334,n49017,n49018 );
   nand U50123 ( n49018,n45341,n28094 );
   and U50124 ( n49017,n49019,n49020 );
   nand U50125 ( n49022,n28284,p1_eax_reg_15_ );
   nor U50126 ( n49021,n49024,n49025 );
   nor U50127 ( n49025,n28399,n49026 );
   nor U50128 ( n49024,n49027,n28258 );
   nand U50129 ( n49030,n49023,p1_eax_reg_14_ );
   nor U50130 ( n49029,n49031,n49032 );
   nor U50131 ( n49031,n28399,n49033 );
   nand U50132 ( n49035,n49023,p1_eax_reg_13_ );
   nor U50133 ( n49034,n49036,n49037 );
   nor U50134 ( n49036,n28401,n49038 );
   nand U50135 ( n49040,n49023,p1_eax_reg_12_ );
   nor U50136 ( n49039,n49041,n49042 );
   nor U50137 ( n49041,n28401,n49043 );
   nand U50138 ( n49045,n49023,p1_eax_reg_11_ );
   nor U50139 ( n49044,n49046,n49047 );
   nor U50140 ( n49046,n28398,n49048 );
   nand U50141 ( n49050,n49023,p1_eax_reg_10_ );
   nor U50142 ( n49049,n49051,n49052 );
   nor U50143 ( n49051,n28398,n49053 );
   nand U50144 ( n49055,n49023,p1_eax_reg_9_ );
   nor U50145 ( n49054,n49056,n49057 );
   nor U50146 ( n49056,n28400,n49058 );
   nand U50147 ( n49060,n49023,p1_eax_reg_8_ );
   nor U50148 ( n49059,n49061,n49062 );
   nor U50149 ( n49061,n28398,n49063 );
   nand U50150 ( n49065,n49023,p1_eax_reg_7_ );
   nor U50151 ( n49064,n49066,n49067 );
   nor U50152 ( n49066,n28400,n49068 );
   nand U50153 ( n49070,n49023,p1_eax_reg_6_ );
   nor U50154 ( n49069,n49071,n49072 );
   nor U50155 ( n49071,n28400,n49073 );
   nand U50156 ( n49075,n49023,p1_eax_reg_5_ );
   nor U50157 ( n49074,n49076,n49077 );
   nor U50158 ( n49076,n28398,n49078 );
   nand U50159 ( n49080,n49023,p1_eax_reg_4_ );
   nor U50160 ( n49079,n49081,n49082 );
   nor U50161 ( n49081,n28399,n49083 );
   nand U50162 ( n49085,n49023,p1_eax_reg_3_ );
   nor U50163 ( n49084,n49086,n49087 );
   nor U50164 ( n49086,n28398,n49088 );
   nand U50165 ( n49090,n49023,p1_eax_reg_2_ );
   nor U50166 ( n49089,n49091,n49092 );
   nor U50167 ( n49091,n28400,n49093 );
   nand U50168 ( n49095,n49023,p1_eax_reg_1_ );
   nor U50169 ( n49094,n49096,n49097 );
   nor U50170 ( n49096,n28400,n49098 );
   nand U50171 ( n49100,n49023,p1_eax_reg_0_ );
   nor U50172 ( n49099,n49101,n49102 );
   nor U50173 ( n49101,n28400,n49103 );
   nand U50174 ( n49105,n49023,p1_eax_reg_30_ );
   nor U50175 ( n49104,n49106,n49032 );
   nor U50176 ( n49032,n49028,n49107 );
   nor U50177 ( n49106,n28399,n49108 );
   nand U50178 ( n49110,n28284,p1_eax_reg_29_ );
   nor U50179 ( n49109,n49111,n49037 );
   nor U50180 ( n49037,n49028,n49112 );
   nor U50181 ( n49111,n28401,n49113 );
   nand U50182 ( n49115,n28284,p1_eax_reg_28_ );
   nor U50183 ( n49114,n49116,n49042 );
   nor U50184 ( n49042,n49028,n49117 );
   nor U50185 ( n49116,n28401,n49118 );
   nand U50186 ( n49120,n28284,p1_eax_reg_27_ );
   nor U50187 ( n49119,n49121,n49047 );
   nor U50188 ( n49047,n49028,n49122 );
   nor U50189 ( n49121,n28399,n49123 );
   nand U50190 ( n49125,n28284,p1_eax_reg_26_ );
   nor U50191 ( n49124,n49126,n49052 );
   nor U50192 ( n49052,n49028,n49127 );
   nor U50193 ( n49126,n28399,n49128 );
   nand U50194 ( n49130,n28284,p1_eax_reg_25_ );
   nor U50195 ( n49129,n49131,n49057 );
   nor U50196 ( n49057,n49028,n49132 );
   nor U50197 ( n49131,n28398,n49133 );
   nand U50198 ( n49135,n28284,p1_eax_reg_24_ );
   nor U50199 ( n49134,n49136,n49062 );
   nor U50200 ( n49062,n49028,n49137 );
   nor U50201 ( n49136,n28400,n49138 );
   nand U50202 ( n49140,n28284,p1_eax_reg_23_ );
   nor U50203 ( n49139,n49141,n49067 );
   nor U50204 ( n49067,n47246,n28258 );
   nor U50205 ( n49141,n28400,n49142 );
   nand U50206 ( n49144,n28284,p1_eax_reg_22_ );
   nor U50207 ( n49143,n49145,n49072 );
   nor U50208 ( n49072,n47262,n28258 );
   nor U50209 ( n49145,n28399,n49146 );
   nand U50210 ( n49148,n28284,p1_eax_reg_21_ );
   nor U50211 ( n49147,n49149,n49077 );
   nor U50212 ( n49077,n47278,n49028 );
   nor U50213 ( n49149,n28399,n49150 );
   nand U50214 ( n49152,n28284,p1_eax_reg_20_ );
   nor U50215 ( n49151,n49153,n49082 );
   nor U50216 ( n49082,n47294,n49028 );
   nor U50217 ( n49153,n28401,n49154 );
   nand U50218 ( n49156,n28284,p1_eax_reg_19_ );
   nor U50219 ( n49155,n49157,n49087 );
   nor U50220 ( n49087,n47310,n49028 );
   nor U50221 ( n49157,n28401,n49158 );
   nand U50222 ( n49160,n28284,p1_eax_reg_18_ );
   nor U50223 ( n49159,n49161,n49092 );
   nor U50224 ( n49092,n47325,n28258 );
   nor U50225 ( n49161,n28398,n49162 );
   nand U50226 ( n49164,n28284,p1_eax_reg_17_ );
   nor U50227 ( n49163,n49165,n49097 );
   nor U50228 ( n49097,n47341,n28258 );
   nor U50229 ( n49165,n28398,n49166 );
   nand U50230 ( n49168,n28284,p1_eax_reg_16_ );
   and U50231 ( n49023,n28401,n48289 );
   nor U50232 ( n49167,n49169,n49102 );
   nor U50233 ( n49102,n47359,n28258 );
   nand U50234 ( n49028,n28399,n47334 );
   nor U50235 ( n49169,n28401,n49170 );
   nor U50236 ( n49172,n45876,n49173 );
   nor U50237 ( n49173,n45358,n45346 );
   nor U50238 ( n49171,n47433,n48283 );
   nand U50239 ( n49175,n28364,p1_datao_reg_0_ );
   nor U50240 ( n49174,n49177,n49178 );
   nor U50241 ( n49178,n49179,n49180 );
   nor U50242 ( n49177,n49103,n28098 );
   not U50243 ( n49103,p1_lword_reg_0_ );
   nand U50244 ( n49182,n28364,p1_datao_reg_1_ );
   nor U50245 ( n49181,n49183,n49184 );
   and U50246 ( n49184,p1_eax_reg_1_,n49185 );
   nor U50247 ( n49183,n49098,n28096 );
   not U50248 ( n49098,p1_lword_reg_1_ );
   nand U50249 ( n49187,n49176,p1_datao_reg_2_ );
   nor U50250 ( n49186,n49188,n49189 );
   nor U50251 ( n49189,n49190,n49180 );
   nor U50252 ( n49188,n49093,n28097 );
   not U50253 ( n49093,p1_lword_reg_2_ );
   nand U50254 ( n49192,n49176,p1_datao_reg_3_ );
   nor U50255 ( n49191,n49193,n49194 );
   nor U50256 ( n49194,n49195,n49180 );
   nor U50257 ( n49193,n49088,n28098 );
   not U50258 ( n49088,p1_lword_reg_3_ );
   nand U50259 ( n49197,n49176,p1_datao_reg_4_ );
   nor U50260 ( n49196,n49198,n49199 );
   nor U50261 ( n49199,n49200,n49180 );
   nor U50262 ( n49198,n49083,n28096 );
   not U50263 ( n49083,p1_lword_reg_4_ );
   nand U50264 ( n49202,n49176,p1_datao_reg_5_ );
   nor U50265 ( n49201,n49203,n49204 );
   and U50266 ( n49204,p1_eax_reg_5_,n49185 );
   nor U50267 ( n49203,n49078,n28097 );
   not U50268 ( n49078,p1_lword_reg_5_ );
   nand U50269 ( n49206,n49176,p1_datao_reg_6_ );
   nor U50270 ( n49205,n49207,n49208 );
   nor U50271 ( n49208,n49209,n49180 );
   nor U50272 ( n49207,n49073,n28098 );
   not U50273 ( n49073,p1_lword_reg_6_ );
   nand U50274 ( n49211,n49176,p1_datao_reg_7_ );
   nor U50275 ( n49210,n49212,n49213 );
   nor U50276 ( n49213,n49214,n49180 );
   nor U50277 ( n49212,n49068,n28096 );
   not U50278 ( n49068,p1_lword_reg_7_ );
   nand U50279 ( n49216,n49176,p1_datao_reg_8_ );
   nor U50280 ( n49215,n49217,n49218 );
   nor U50281 ( n49218,n49219,n49180 );
   nor U50282 ( n49217,n49063,n28097 );
   not U50283 ( n49063,p1_lword_reg_8_ );
   nand U50284 ( n49221,n49176,p1_datao_reg_9_ );
   nor U50285 ( n49220,n49222,n49223 );
   nor U50286 ( n49223,n49224,n49180 );
   nor U50287 ( n49222,n49058,n28098 );
   not U50288 ( n49058,p1_lword_reg_9_ );
   nand U50289 ( n49226,n49176,p1_datao_reg_10_ );
   nor U50290 ( n49225,n49227,n49228 );
   and U50291 ( n49228,p1_eax_reg_10_,n49185 );
   nor U50292 ( n49227,n49053,n28096 );
   not U50293 ( n49053,p1_lword_reg_10_ );
   nand U50294 ( n49230,n49176,p1_datao_reg_11_ );
   nor U50295 ( n49229,n49231,n49232 );
   nor U50296 ( n49232,n49233,n49180 );
   nor U50297 ( n49231,n49048,n28097 );
   not U50298 ( n49048,p1_lword_reg_11_ );
   nand U50299 ( n49235,n49176,p1_datao_reg_12_ );
   nor U50300 ( n49234,n49236,n49237 );
   nor U50301 ( n49237,n49238,n49180 );
   nor U50302 ( n49236,n49043,n28098 );
   not U50303 ( n49043,p1_lword_reg_12_ );
   nand U50304 ( n49240,n49176,p1_datao_reg_13_ );
   nor U50305 ( n49239,n49241,n49242 );
   nor U50306 ( n49242,n49243,n49180 );
   not U50307 ( n49180,n49185 );
   nor U50308 ( n49241,n49038,n28096 );
   not U50309 ( n49038,p1_lword_reg_13_ );
   nand U50310 ( n49245,n49176,p1_datao_reg_14_ );
   nor U50311 ( n49244,n49246,n49247 );
   and U50312 ( n49247,p1_eax_reg_14_,n49185 );
   nor U50313 ( n49246,n49033,n28097 );
   not U50314 ( n49033,p1_lword_reg_14_ );
   nand U50315 ( n49249,n49176,p1_datao_reg_15_ );
   nor U50316 ( n49248,n49250,n49251 );
   and U50317 ( n49251,p1_eax_reg_15_,n49185 );
   nor U50318 ( n49250,n49026,n28098 );
   not U50319 ( n49026,p1_lword_reg_15_ );
   nand U50320 ( n49253,n28364,p1_datao_reg_16_ );
   nor U50321 ( n49252,n49254,n49255 );
   nor U50322 ( n49255,n49256,n49257 );
   nor U50323 ( n49254,n49170,n28096 );
   not U50324 ( n49170,p1_uword_reg_0_ );
   nand U50325 ( n49259,n28364,p1_datao_reg_17_ );
   nor U50326 ( n49258,n49260,n49261 );
   nor U50327 ( n49261,n49262,n27881 );
   nor U50328 ( n49260,n49166,n28097 );
   not U50329 ( n49166,p1_uword_reg_1_ );
   nand U50330 ( n49264,n28364,p1_datao_reg_18_ );
   nor U50331 ( n49263,n49265,n49266 );
   nor U50332 ( n49266,n49267,n27881 );
   nor U50333 ( n49265,n49162,n28098 );
   not U50334 ( n49162,p1_uword_reg_2_ );
   nand U50335 ( n49269,n28364,p1_datao_reg_19_ );
   nor U50336 ( n49268,n49270,n49271 );
   nor U50337 ( n49271,n49272,n27881 );
   nor U50338 ( n49270,n49158,n28096 );
   not U50339 ( n49158,p1_uword_reg_3_ );
   nand U50340 ( n49274,n28364,p1_datao_reg_20_ );
   nor U50341 ( n49273,n49275,n49276 );
   nor U50342 ( n49276,n49277,n49257 );
   nor U50343 ( n49275,n49154,n28097 );
   not U50344 ( n49154,p1_uword_reg_4_ );
   nand U50345 ( n49279,n28364,p1_datao_reg_21_ );
   nor U50346 ( n49278,n49280,n49281 );
   nor U50347 ( n49281,n49282,n49257 );
   nor U50348 ( n49280,n49150,n28098 );
   not U50349 ( n49150,p1_uword_reg_5_ );
   nand U50350 ( n49284,n28364,p1_datao_reg_22_ );
   nor U50351 ( n49283,n49285,n49286 );
   nor U50352 ( n49286,n49287,n49257 );
   nor U50353 ( n49285,n49146,n28096 );
   not U50354 ( n49146,p1_uword_reg_6_ );
   nand U50355 ( n49289,n28364,p1_datao_reg_23_ );
   nor U50356 ( n49288,n49290,n49291 );
   nor U50357 ( n49291,n49292,n49257 );
   nor U50358 ( n49290,n49142,n28097 );
   not U50359 ( n49142,p1_uword_reg_7_ );
   nand U50360 ( n49294,n28364,p1_datao_reg_24_ );
   nor U50361 ( n49293,n49295,n49296 );
   nor U50362 ( n49296,n49297,n49257 );
   nor U50363 ( n49295,n49138,n28098 );
   not U50364 ( n49138,p1_uword_reg_8_ );
   nand U50365 ( n49299,n28364,p1_datao_reg_25_ );
   nor U50366 ( n49298,n49300,n49301 );
   nor U50367 ( n49301,n49302,n49257 );
   nor U50368 ( n49300,n49133,n28096 );
   not U50369 ( n49133,p1_uword_reg_9_ );
   nand U50370 ( n49304,n28364,p1_datao_reg_26_ );
   nor U50371 ( n49303,n49305,n49306 );
   nor U50372 ( n49306,n49307,n49257 );
   nor U50373 ( n49305,n49128,n28097 );
   not U50374 ( n49128,p1_uword_reg_10_ );
   nand U50375 ( n49309,n28364,p1_datao_reg_27_ );
   nor U50376 ( n49308,n49310,n49311 );
   nor U50377 ( n49311,n49312,n49257 );
   nor U50378 ( n49310,n49123,n28098 );
   not U50379 ( n49123,p1_uword_reg_11_ );
   nand U50380 ( n49314,n28364,p1_datao_reg_28_ );
   nor U50381 ( n49313,n49315,n49316 );
   nor U50382 ( n49316,n49317,n49257 );
   nor U50383 ( n49315,n49118,n28096 );
   not U50384 ( n49118,p1_uword_reg_12_ );
   nand U50385 ( n49319,n28364,p1_datao_reg_29_ );
   nor U50386 ( n49318,n49320,n49321 );
   nor U50387 ( n49321,n49322,n49257 );
   nor U50388 ( n49320,n49113,n28097 );
   not U50389 ( n49113,p1_uword_reg_13_ );
   nand U50390 ( n49324,n28364,p1_datao_reg_30_ );
   nor U50391 ( n49323,n49325,n49326 );
   nor U50392 ( n49326,n49327,n49257 );
   nand U50393 ( n49257,n49185,n47351 );
   nor U50394 ( n49185,n28095,n49176 );
   not U50395 ( n49176,n49328 );
   nor U50396 ( n49325,n49108,n28097 );
   not U50397 ( n49108,p1_uword_reg_14_ );
   nand U50398 ( n49328,n49329,n49330 );
   nand U50399 ( n49330,n49331,n45360 );
   nor U50400 ( n49331,n49332,n48283 );
   nor U50401 ( n49332,n45797,n45444 );
   not U50402 ( n45444,n45836 );
   nor U50403 ( n45797,n48912,n47433 );
   nand U50404 ( n49329,n45503,n28094 );
   nor U50405 ( n45503,n45432,n28375 );
   not U50406 ( n28479,p1_datao_reg_31_ );
   nand U50407 ( n49334,n49335,p1_eax_reg_0_ );
   nor U50408 ( n49333,n49336,n49337 );
   nor U50409 ( n49337,n48304,n49338 );
   nor U50410 ( n49336,n47359,n49339 );
   not U50411 ( n47359,n49340 );
   nand U50412 ( n49342,n28261,p1_eax_reg_1_ );
   nor U50413 ( n49341,n49343,n49344 );
   nor U50414 ( n49344,n48310,n49338 );
   nor U50415 ( n49343,n47341,n28224 );
   not U50416 ( n47341,n49345 );
   nand U50417 ( n49347,n28261,p1_eax_reg_2_ );
   nor U50418 ( n49346,n49348,n49349 );
   nor U50419 ( n49349,n49350,n28307 );
   nor U50420 ( n49348,n47325,n28224 );
   not U50421 ( n47325,n49351 );
   nand U50422 ( n49353,n49335,p1_eax_reg_3_ );
   nor U50423 ( n49352,n49354,n49355 );
   nor U50424 ( n49355,n49356,n49338 );
   nor U50425 ( n49354,n47310,n28224 );
   not U50426 ( n47310,n49357 );
   nand U50427 ( n49359,n49335,p1_eax_reg_4_ );
   nor U50428 ( n49358,n49360,n49361 );
   nor U50429 ( n49361,n49362,n49338 );
   nor U50430 ( n49360,n47294,n49339 );
   not U50431 ( n47294,n49363 );
   nand U50432 ( n49365,n28261,p1_eax_reg_5_ );
   nor U50433 ( n49364,n49366,n49367 );
   nor U50434 ( n49367,n49368,n28307 );
   nor U50435 ( n49366,n47278,n49339 );
   not U50436 ( n47278,n49369 );
   nand U50437 ( n49371,n49335,p1_eax_reg_6_ );
   nor U50438 ( n49370,n49372,n49373 );
   nor U50439 ( n49373,n49374,n28307 );
   nor U50440 ( n49372,n47262,n49339 );
   not U50441 ( n47262,n49375 );
   nand U50442 ( n49377,n49335,p1_eax_reg_7_ );
   nor U50443 ( n49376,n49378,n49379 );
   nor U50444 ( n49379,n49380,n49338 );
   nor U50445 ( n49378,n47246,n49339 );
   not U50446 ( n47246,n49381 );
   nand U50447 ( n49383,n28261,p1_eax_reg_8_ );
   nor U50448 ( n49382,n49384,n49385 );
   nor U50449 ( n49385,n49386,n49338 );
   nor U50450 ( n49384,n49137,n49339 );
   not U50451 ( n49137,n49387 );
   nand U50452 ( n49389,n49335,p1_eax_reg_9_ );
   nor U50453 ( n49388,n49390,n49391 );
   nor U50454 ( n49391,n49392,n49338 );
   nor U50455 ( n49390,n49132,n49339 );
   not U50456 ( n49132,n49393 );
   nand U50457 ( n49395,n49335,p1_eax_reg_10_ );
   nor U50458 ( n49394,n49396,n49397 );
   nor U50459 ( n49397,n49398,n49338 );
   nor U50460 ( n49396,n49127,n49339 );
   not U50461 ( n49127,n49399 );
   nand U50462 ( n49401,n49335,p1_eax_reg_11_ );
   nor U50463 ( n49400,n49402,n49403 );
   nor U50464 ( n49403,n49404,n49338 );
   nor U50465 ( n49402,n49122,n49339 );
   not U50466 ( n49122,n49405 );
   nand U50467 ( n49407,n28261,p1_eax_reg_12_ );
   nor U50468 ( n49406,n49408,n49409 );
   nor U50469 ( n49409,n49410,n49338 );
   nor U50470 ( n49408,n49117,n49339 );
   not U50471 ( n49117,n49411 );
   nand U50472 ( n49413,n28261,p1_eax_reg_13_ );
   nor U50473 ( n49412,n49414,n49415 );
   nor U50474 ( n49415,n49416,n49338 );
   nor U50475 ( n49414,n49112,n49339 );
   not U50476 ( n49112,n49417 );
   nand U50477 ( n49419,n49335,p1_eax_reg_14_ );
   nor U50478 ( n49418,n49420,n49421 );
   nor U50479 ( n49421,n49422,n49338 );
   nor U50480 ( n49420,n49107,n28224 );
   not U50481 ( n49107,n49423 );
   nand U50482 ( n49425,n49335,p1_eax_reg_15_ );
   nor U50483 ( n49424,n49426,n49427 );
   nor U50484 ( n49427,n49428,n49338 );
   nor U50485 ( n49426,n49027,n49339 );
   nand U50486 ( n49339,n49429,n28243 );
   nor U50487 ( n49429,n49431,n47426 );
   and U50488 ( n49027,n49432,n49433 );
   nand U50489 ( n49433,datai_15_,n28329 );
   nand U50490 ( n49432,buf1_reg_15_,n27894 );
   nor U50491 ( n49435,n49436,n49437 );
   nand U50492 ( n49437,n49438,n49439 );
   nand U50493 ( n49439,n49440,n49340 );
   nor U50494 ( n49340,n49441,n49442 );
   nor U50495 ( n49442,datai_0_,n27894 );
   nor U50496 ( n49441,buf1_reg_0_,n28765 );
   nand U50497 ( n49438,n49443,n48568 );
   nor U50498 ( n49436,n49444,n49445 );
   not U50499 ( n49444,datai_16_ );
   nor U50500 ( n49434,n49446,n49447 );
   nor U50501 ( n49447,n49256,n49430 );
   nor U50502 ( n49446,n28647,n49448 );
   not U50503 ( n28647,buf1_reg_16_ );
   nor U50504 ( n49450,n49451,n49452 );
   nand U50505 ( n49452,n49453,n49454 );
   nand U50506 ( n49454,n49440,n49345 );
   nor U50507 ( n49345,n49455,n49456 );
   nor U50508 ( n49456,datai_1_,n27894 );
   nor U50509 ( n49455,buf1_reg_1_,n28765 );
   nand U50510 ( n49453,n49443,n48583 );
   nor U50511 ( n49451,n49457,n28212 );
   not U50512 ( n49457,datai_17_ );
   nor U50513 ( n49449,n49458,n49459 );
   nor U50514 ( n49459,n49262,n49430 );
   nor U50515 ( n49458,n28653,n28223 );
   not U50516 ( n28653,buf1_reg_17_ );
   nor U50517 ( n49461,n49462,n49463 );
   nand U50518 ( n49463,n49464,n49465 );
   nand U50519 ( n49465,n49440,n49351 );
   nor U50520 ( n49351,n49466,n49467 );
   nor U50521 ( n49467,datai_2_,n27894 );
   nor U50522 ( n49466,buf1_reg_2_,n28329 );
   nand U50523 ( n49464,n49443,n48601 );
   nor U50524 ( n49462,n49468,n28212 );
   not U50525 ( n49468,datai_18_ );
   nor U50526 ( n49460,n49469,n49470 );
   nor U50527 ( n49470,n49267,n49430 );
   nor U50528 ( n49469,n28659,n28223 );
   not U50529 ( n28659,buf1_reg_18_ );
   nor U50530 ( n49472,n49473,n49474 );
   nand U50531 ( n49474,n49475,n49476 );
   nand U50532 ( n49476,n49440,n49357 );
   nor U50533 ( n49357,n49477,n49478 );
   nor U50534 ( n49478,datai_3_,n47355 );
   nor U50535 ( n49477,buf1_reg_3_,n28329 );
   nand U50536 ( n49475,n49443,n48616 );
   nor U50537 ( n49473,n49479,n28212 );
   not U50538 ( n49479,datai_19_ );
   nor U50539 ( n49471,n49480,n49481 );
   nor U50540 ( n49481,n49272,n49430 );
   nor U50541 ( n49480,n28665,n28223 );
   not U50542 ( n28665,buf1_reg_19_ );
   nor U50543 ( n49483,n49484,n49485 );
   nand U50544 ( n49485,n49486,n49487 );
   nand U50545 ( n49487,n49440,n49363 );
   nor U50546 ( n49363,n49488,n49489 );
   nor U50547 ( n49489,datai_4_,n47355 );
   nor U50548 ( n49488,buf1_reg_4_,n28765 );
   nand U50549 ( n49486,n49443,n48631 );
   nor U50550 ( n49484,n49490,n49445 );
   not U50551 ( n49490,datai_20_ );
   nor U50552 ( n49482,n49491,n49492 );
   nor U50553 ( n49492,n49277,n28243 );
   nor U50554 ( n49491,n28671,n49448 );
   not U50555 ( n28671,buf1_reg_20_ );
   nor U50556 ( n49494,n49495,n49496 );
   nand U50557 ( n49496,n49497,n49498 );
   nand U50558 ( n49498,n49440,n49369 );
   nor U50559 ( n49369,n49499,n49500 );
   nor U50560 ( n49500,datai_5_,n47355 );
   nor U50561 ( n49499,buf1_reg_5_,n28765 );
   nand U50562 ( n49497,n49443,n48651 );
   nor U50563 ( n49495,n49501,n49445 );
   not U50564 ( n49501,datai_21_ );
   nor U50565 ( n49493,n49502,n49503 );
   nor U50566 ( n49503,n49282,n28243 );
   nor U50567 ( n49502,n28677,n49448 );
   not U50568 ( n28677,buf1_reg_21_ );
   nor U50569 ( n49505,n49506,n49507 );
   nand U50570 ( n49507,n49508,n49509 );
   nand U50571 ( n49509,n49440,n49375 );
   nor U50572 ( n49375,n49510,n49511 );
   nor U50573 ( n49511,datai_6_,n47355 );
   nor U50574 ( n49510,buf1_reg_6_,n28765 );
   nand U50575 ( n49508,n49443,n48671 );
   nor U50576 ( n49506,n49512,n49445 );
   not U50577 ( n49512,datai_22_ );
   nor U50578 ( n49504,n49513,n49514 );
   nor U50579 ( n49514,n49287,n49430 );
   nor U50580 ( n49513,n28683,n49448 );
   not U50581 ( n28683,buf1_reg_22_ );
   nor U50582 ( n49516,n49517,n49518 );
   nand U50583 ( n49518,n49519,n49520 );
   nand U50584 ( n49520,n49440,n49381 );
   nor U50585 ( n49381,n49521,n49522 );
   nor U50586 ( n49522,datai_7_,n47355 );
   nor U50587 ( n49521,buf1_reg_7_,n28329 );
   nand U50588 ( n49519,n49443,n48690 );
   nor U50589 ( n49517,n49523,n49445 );
   not U50590 ( n49523,datai_23_ );
   nor U50591 ( n49515,n49524,n49525 );
   nor U50592 ( n49525,n49292,n49430 );
   nor U50593 ( n49524,n28689,n49448 );
   not U50594 ( n28689,buf1_reg_23_ );
   nor U50595 ( n49527,n49528,n49529 );
   nand U50596 ( n49529,n49530,n49531 );
   nand U50597 ( n49531,n49440,n49387 );
   nor U50598 ( n49387,n49532,n49533 );
   nor U50599 ( n49533,datai_8_,n47355 );
   nor U50600 ( n49532,buf1_reg_8_,n28765 );
   nand U50601 ( n49530,n49443,n48704 );
   nor U50602 ( n49528,n49534,n49445 );
   not U50603 ( n49534,datai_24_ );
   nor U50604 ( n49526,n49535,n49536 );
   nor U50605 ( n49536,n49297,n49430 );
   nor U50606 ( n49535,n28695,n49448 );
   not U50607 ( n28695,buf1_reg_24_ );
   nor U50608 ( n49538,n49539,n49540 );
   nand U50609 ( n49540,n49541,n49542 );
   nand U50610 ( n49542,n49440,n49393 );
   nor U50611 ( n49393,n49543,n49544 );
   nor U50612 ( n49544,datai_9_,n47355 );
   nor U50613 ( n49543,buf1_reg_9_,n28765 );
   nand U50614 ( n49541,n49443,n48723 );
   nor U50615 ( n49539,n49545,n49445 );
   not U50616 ( n49545,datai_25_ );
   nor U50617 ( n49537,n49546,n49547 );
   nor U50618 ( n49547,n49302,n49430 );
   not U50619 ( n49302,p1_eax_reg_25_ );
   nor U50620 ( n49546,n28701,n49448 );
   not U50621 ( n28701,buf1_reg_25_ );
   nor U50622 ( n49549,n49550,n49551 );
   nand U50623 ( n49551,n49552,n49553 );
   nand U50624 ( n49553,n49440,n49399 );
   nor U50625 ( n49399,n49554,n49555 );
   nor U50626 ( n49555,datai_10_,n47355 );
   nor U50627 ( n49554,buf1_reg_10_,n28765 );
   nand U50628 ( n49552,n49443,n48738 );
   nor U50629 ( n49550,n49556,n49445 );
   not U50630 ( n49556,datai_26_ );
   nor U50631 ( n49548,n49557,n49558 );
   nor U50632 ( n49558,n49307,n49430 );
   nor U50633 ( n49557,n28707,n49448 );
   not U50634 ( n28707,buf1_reg_26_ );
   nor U50635 ( n49560,n49561,n49562 );
   nand U50636 ( n49562,n49563,n49564 );
   nand U50637 ( n49564,n49440,n49405 );
   nor U50638 ( n49405,n49565,n49566 );
   nor U50639 ( n49566,datai_11_,n27894 );
   nor U50640 ( n49565,buf1_reg_11_,n28329 );
   nand U50641 ( n49563,n49443,n48761 );
   nor U50642 ( n49561,n49567,n49445 );
   not U50643 ( n49567,datai_27_ );
   nor U50644 ( n49559,n49568,n49569 );
   nor U50645 ( n49569,n49312,n49430 );
   not U50646 ( n49312,p1_eax_reg_27_ );
   nor U50647 ( n49568,n28713,n49448 );
   not U50648 ( n28713,buf1_reg_27_ );
   nor U50649 ( n49571,n49572,n49573 );
   nand U50650 ( n49573,n49574,n49575 );
   nand U50651 ( n49575,n49440,n49411 );
   nor U50652 ( n49411,n49576,n49577 );
   nor U50653 ( n49577,datai_12_,n47355 );
   nor U50654 ( n49576,buf1_reg_12_,n28765 );
   nand U50655 ( n49574,n49443,n48783 );
   nor U50656 ( n49572,n49578,n49445 );
   not U50657 ( n49578,datai_28_ );
   nor U50658 ( n49570,n49579,n49580 );
   nor U50659 ( n49580,n49317,n49430 );
   nor U50660 ( n49579,n28719,n49448 );
   not U50661 ( n28719,buf1_reg_28_ );
   nor U50662 ( n49582,n49583,n49584 );
   nand U50663 ( n49584,n49585,n49586 );
   nand U50664 ( n49586,n49440,n49417 );
   nor U50665 ( n49417,n49587,n49588 );
   nor U50666 ( n49588,datai_13_,n47355 );
   nor U50667 ( n49587,buf1_reg_13_,n28329 );
   nand U50668 ( n49585,n49443,n48798 );
   nor U50669 ( n49583,n49589,n49445 );
   not U50670 ( n49589,datai_29_ );
   nor U50671 ( n49581,n49590,n49591 );
   nor U50672 ( n49591,n49322,n49430 );
   nor U50673 ( n49590,n28725,n49448 );
   not U50674 ( n28725,buf1_reg_29_ );
   nor U50675 ( n49593,n49594,n49595 );
   nand U50676 ( n49595,n49596,n49597 );
   nand U50677 ( n49597,n49443,n48824 );
   not U50678 ( n49443,n49338 );
   nand U50679 ( n49338,n28243,n49598 );
   nand U50680 ( n49598,n47236,n48260 );
   nand U50681 ( n49596,n49440,n49423 );
   nor U50682 ( n49423,n49599,n49600 );
   nor U50683 ( n49600,datai_14_,n47355 );
   nor U50684 ( n49599,buf1_reg_14_,n28329 );
   and U50685 ( n49440,n49601,n49602 );
   nor U50686 ( n49601,n47426,n49335 );
   nor U50687 ( n49594,n49603,n28212 );
   not U50688 ( n49603,datai_30_ );
   nor U50689 ( n49592,n49604,n49605 );
   nor U50690 ( n49605,n49327,n49430 );
   nor U50691 ( n49604,n28731,n28223 );
   not U50692 ( n28731,buf1_reg_30_ );
   nor U50693 ( n49607,n49608,n49609 );
   and U50694 ( n49609,p1_eax_reg_31_,n28261 );
   nor U50695 ( n49608,n49335,n49610 );
   nand U50696 ( n49610,n47426,n48835 );
   nor U50697 ( n49606,n49611,n49612 );
   nor U50698 ( n49612,n28736,n49448 );
   nand U50699 ( n49448,n49613,n49614 );
   nor U50700 ( n49613,n49335,n28329 );
   not U50701 ( n28736,buf1_reg_31_ );
   nor U50702 ( n49611,n49615,n49445 );
   nand U50703 ( n49445,n49616,n49614 );
   nor U50704 ( n49616,n47355,n49335 );
   not U50705 ( n49335,n49430 );
   nand U50706 ( n49430,n49617,n49618 );
   nand U50707 ( n49618,n49619,n47457 );
   nor U50708 ( n47457,n47433,n49620 );
   nor U50709 ( n49619,n45701,n48283 );
   nand U50710 ( n49617,n49621,n49622 );
   nor U50711 ( n49621,n49623,n49624 );
   nor U50712 ( n49623,n49625,n49626 );
   nand U50713 ( n49626,n49627,n49628 );
   nand U50714 ( n49628,n49629,n45853 );
   nor U50715 ( n49629,n45880,n45877 );
   nand U50716 ( n49627,n47444,n49630 );
   nor U50717 ( n47444,n45701,n45865 );
   nor U50718 ( n49625,n49631,n49632 );
   not U50719 ( n47355,n28765 );
   nand U50720 ( n28765,p1_address_reg_29_,n49633 );
   nand U50721 ( n49633,n49634,n49635 );
   nor U50722 ( n49635,n49636,n49637 );
   nand U50723 ( n49637,n49638,n49639 );
   nor U50724 ( n49639,n49640,n49641 );
   or U50725 ( n49641,p1_address_reg_25_,p1_address_reg_26_ );
   or U50726 ( n49640,p1_address_reg_27_,p1_address_reg_28_ );
   nor U50727 ( n49638,p1_address_reg_22_,n49642 );
   or U50728 ( n49642,p1_address_reg_23_,p1_address_reg_24_ );
   nand U50729 ( n49636,n49643,n49644 );
   nor U50730 ( n49644,n49645,n49646 );
   or U50731 ( n49646,p1_address_reg_6_,p1_address_reg_7_ );
   or U50732 ( n49645,p1_address_reg_8_,p1_address_reg_9_ );
   nor U50733 ( n49643,n49647,n49648 );
   or U50734 ( n49648,p1_address_reg_2_,p1_address_reg_3_ );
   or U50735 ( n49647,p1_address_reg_4_,p1_address_reg_5_ );
   nor U50736 ( n49634,n49649,n49650 );
   nand U50737 ( n49650,n49651,n49652 );
   nor U50738 ( n49652,n49653,n49654 );
   or U50739 ( n49654,p1_address_reg_12_,p1_address_reg_13_ );
   or U50740 ( n49653,p1_address_reg_14_,p1_address_reg_15_ );
   nor U50741 ( n49651,p1_address_reg_0_,n49655 );
   or U50742 ( n49655,p1_address_reg_10_,p1_address_reg_11_ );
   nand U50743 ( n49649,n49656,n49657 );
   nor U50744 ( n49657,n49658,n49659 );
   or U50745 ( n49659,p1_address_reg_19_,p1_address_reg_1_ );
   or U50746 ( n49658,p1_address_reg_20_,p1_address_reg_21_ );
   nor U50747 ( n49656,p1_address_reg_16_,n49660 );
   or U50748 ( n49660,p1_address_reg_17_,p1_address_reg_18_ );
   not U50749 ( n49615,datai_31_ );
   nand U50750 ( n49662,p1_ebx_reg_0_,n28348 );
   nor U50751 ( n49661,n49664,n49665 );
   nor U50752 ( n49665,n47475,n28102 );
   not U50753 ( n47475,n49667 );
   nor U50754 ( n49664,n48304,n28110 );
   nand U50755 ( n49669,p1_ebx_reg_1_,n28348 );
   nor U50756 ( n49668,n49670,n49671 );
   nor U50757 ( n49671,n47492,n28103 );
   not U50758 ( n47492,n49672 );
   nor U50759 ( n49670,n48310,n28110 );
   nand U50760 ( n49674,p1_ebx_reg_2_,n49663 );
   nor U50761 ( n49673,n49675,n49676 );
   nor U50762 ( n49676,n47521,n28103 );
   not U50763 ( n47521,n49677 );
   nor U50764 ( n49675,n49350,n28108 );
   not U50765 ( n49350,n48329 );
   nand U50766 ( n49679,p1_ebx_reg_3_,n28348 );
   nor U50767 ( n49678,n49680,n49681 );
   nor U50768 ( n49681,n47541,n28102 );
   not U50769 ( n47541,n49682 );
   nor U50770 ( n49680,n49356,n28108 );
   not U50771 ( n49356,n48345 );
   nand U50772 ( n49684,p1_ebx_reg_4_,n49663 );
   nor U50773 ( n49683,n49685,n49686 );
   nor U50774 ( n49686,n47567,n49666 );
   nor U50775 ( n49685,n49362,n28109 );
   not U50776 ( n49362,n48359 );
   nand U50777 ( n49688,p1_ebx_reg_5_,n49663 );
   nor U50778 ( n49687,n49689,n49690 );
   nor U50779 ( n49690,n47586,n28103 );
   not U50780 ( n47586,n49691 );
   nor U50781 ( n49689,n49368,n28109 );
   not U50782 ( n49368,n48373 );
   nand U50783 ( n49693,p1_ebx_reg_6_,n49663 );
   nor U50784 ( n49692,n49694,n49695 );
   nor U50785 ( n49695,n47614,n28102 );
   nor U50786 ( n49694,n49374,n28110 );
   not U50787 ( n49374,n48387 );
   nand U50788 ( n49697,p1_ebx_reg_7_,n49663 );
   nor U50789 ( n49696,n49698,n49699 );
   nor U50790 ( n49699,n47633,n49666 );
   not U50791 ( n47633,n49700 );
   nor U50792 ( n49698,n49380,n28110 );
   not U50793 ( n49380,n48407 );
   nand U50794 ( n49702,p1_ebx_reg_8_,n49663 );
   nor U50795 ( n49701,n49703,n49704 );
   nor U50796 ( n49704,n47660,n28103 );
   nor U50797 ( n49703,n49386,n28108 );
   not U50798 ( n49386,n48423 );
   nand U50799 ( n49706,p1_ebx_reg_9_,n49663 );
   nor U50800 ( n49705,n49707,n49708 );
   nor U50801 ( n49708,n47679,n28102 );
   not U50802 ( n47679,n49709 );
   nor U50803 ( n49707,n49392,n28108 );
   not U50804 ( n49392,n48441 );
   nand U50805 ( n49711,p1_ebx_reg_10_,n49663 );
   nor U50806 ( n49710,n49712,n49713 );
   nor U50807 ( n49713,n47706,n49666 );
   nor U50808 ( n49712,n49398,n28109 );
   not U50809 ( n49398,n48456 );
   nand U50810 ( n49715,p1_ebx_reg_11_,n49663 );
   nor U50811 ( n49714,n49716,n49717 );
   nor U50812 ( n49717,n47727,n28103 );
   not U50813 ( n47727,n49718 );
   nor U50814 ( n49716,n49404,n28109 );
   nand U50815 ( n49720,p1_ebx_reg_12_,n49663 );
   nor U50816 ( n49719,n49721,n49722 );
   nor U50817 ( n49722,n47754,n28102 );
   nor U50818 ( n49721,n49410,n28109 );
   not U50819 ( n49410,n48492 );
   nand U50820 ( n49724,p1_ebx_reg_13_,n49663 );
   nor U50821 ( n49723,n49725,n49726 );
   nor U50822 ( n49726,n47773,n49666 );
   not U50823 ( n47773,n49727 );
   nor U50824 ( n49725,n49416,n28110 );
   not U50825 ( n49416,n48507 );
   nand U50826 ( n49729,p1_ebx_reg_14_,n49663 );
   nor U50827 ( n49728,n49730,n49731 );
   nor U50828 ( n49731,n47800,n49666 );
   nor U50829 ( n49730,n49422,n28110 );
   not U50830 ( n49422,n48522 );
   nand U50831 ( n49733,p1_ebx_reg_15_,n49663 );
   nor U50832 ( n49732,n49734,n49735 );
   nor U50833 ( n49735,n47821,n28102 );
   not U50834 ( n47821,n49736 );
   nor U50835 ( n49734,n49428,n28109 );
   not U50836 ( n49428,n48547 );
   nand U50837 ( n49738,p1_ebx_reg_16_,n49663 );
   nor U50838 ( n49737,n49739,n49740 );
   nor U50839 ( n49740,n47848,n28103 );
   nor U50840 ( n49739,n49741,n28109 );
   nand U50841 ( n49743,p1_ebx_reg_17_,n49663 );
   nor U50842 ( n49742,n49744,n49745 );
   nor U50843 ( n49745,n47867,n49666 );
   not U50844 ( n47867,n49746 );
   nor U50845 ( n49744,n49747,n28108 );
   not U50846 ( n49747,n48583 );
   nand U50847 ( n49749,p1_ebx_reg_18_,n28348 );
   nor U50848 ( n49748,n49750,n49751 );
   nor U50849 ( n49751,n47894,n28102 );
   nor U50850 ( n49750,n49752,n28108 );
   not U50851 ( n49752,n48601 );
   nand U50852 ( n49754,p1_ebx_reg_19_,n28348 );
   nor U50853 ( n49753,n49755,n49756 );
   nor U50854 ( n49756,n47913,n49666 );
   not U50855 ( n47913,n49757 );
   nor U50856 ( n49755,n49758,n28108 );
   not U50857 ( n49758,n48616 );
   nand U50858 ( n49760,p1_ebx_reg_20_,n28348 );
   nor U50859 ( n49759,n49761,n49762 );
   nor U50860 ( n49762,n47940,n28103 );
   nor U50861 ( n49761,n49763,n28109 );
   not U50862 ( n49763,n48631 );
   nand U50863 ( n49765,p1_ebx_reg_21_,n28348 );
   nor U50864 ( n49764,n49766,n49767 );
   nor U50865 ( n49767,n47959,n28102 );
   not U50866 ( n47959,n49768 );
   nor U50867 ( n49766,n49769,n28109 );
   not U50868 ( n49769,n48651 );
   nand U50869 ( n49771,p1_ebx_reg_22_,n28348 );
   nor U50870 ( n49770,n49772,n49773 );
   nor U50871 ( n49773,n47986,n49666 );
   nor U50872 ( n49772,n49774,n28110 );
   nand U50873 ( n49776,p1_ebx_reg_23_,n28348 );
   nor U50874 ( n49775,n49777,n49778 );
   nor U50875 ( n49778,n48005,n28103 );
   not U50876 ( n48005,n49779 );
   nor U50877 ( n49777,n49780,n28110 );
   not U50878 ( n49780,n48690 );
   nand U50879 ( n49782,p1_ebx_reg_24_,n28348 );
   nor U50880 ( n49781,n49783,n49784 );
   nor U50881 ( n49784,n48032,n28102 );
   nor U50882 ( n49783,n49785,n28108 );
   not U50883 ( n49785,n48704 );
   nand U50884 ( n49787,p1_ebx_reg_25_,n28348 );
   nor U50885 ( n49786,n49788,n49789 );
   nor U50886 ( n49789,n48051,n49666 );
   not U50887 ( n48051,n49790 );
   nor U50888 ( n49788,n49791,n28108 );
   not U50889 ( n49791,n48723 );
   nand U50890 ( n49793,p1_ebx_reg_26_,n28348 );
   nor U50891 ( n49792,n49794,n49795 );
   nor U50892 ( n49795,n48081,n28103 );
   nor U50893 ( n49794,n49796,n28109 );
   nand U50894 ( n49798,p1_ebx_reg_27_,n28348 );
   nor U50895 ( n49797,n49799,n49800 );
   nor U50896 ( n49800,n48100,n28102 );
   not U50897 ( n48100,n49801 );
   nor U50898 ( n49799,n49802,n28109 );
   nand U50899 ( n49804,p1_ebx_reg_28_,n28348 );
   nor U50900 ( n49803,n49805,n49806 );
   nor U50901 ( n49806,n48124,n49666 );
   nor U50902 ( n49805,n49807,n28110 );
   not U50903 ( n49807,n48783 );
   nand U50904 ( n49809,p1_ebx_reg_29_,n28348 );
   nor U50905 ( n49808,n49810,n49811 );
   nor U50906 ( n49811,n48137,n28103 );
   not U50907 ( n48137,n49812 );
   nor U50908 ( n49810,n49813,n28110 );
   not U50909 ( n49813,n48798 );
   nand U50910 ( n49815,p1_ebx_reg_30_,n28348 );
   nor U50911 ( n49814,n49816,n49817 );
   nor U50912 ( n49817,n48150,n28102 );
   not U50913 ( n49666,n49818 );
   not U50914 ( n48150,n49819 );
   nor U50915 ( n49816,n49820,n28108 );
   not U50916 ( n49820,n48824 );
   nand U50917 ( n49822,n49818,n49823 );
   nor U50918 ( n49818,n49663,n47236 );
   nand U50919 ( n49821,p1_ebx_reg_31_,n28348 );
   nand U50920 ( n49663,n45771,n49824 );
   nand U50921 ( n49824,n47450,n49825 );
   nand U50922 ( n49825,n49826,n49827 );
   nor U50923 ( n49826,n49620,n49631 );
   nand U50924 ( n49631,n49828,n49829 );
   nor U50925 ( n49828,n47287,n47236 );
   nand U50926 ( n47450,n47416,n45880 );
   nor U50927 ( n49831,n49832,n49833 );
   nand U50928 ( n49833,n49834,n49835 );
   nand U50929 ( n49835,p1_phyaddrpointer_reg_0_,n49836 );
   nand U50930 ( n49836,n49837,n28279 );
   nand U50931 ( n49834,p1_reip_reg_0_,n49839 );
   nand U50932 ( n49839,n49840,n28250 );
   nor U50933 ( n49832,n49842,n48304 );
   xor U50934 ( n48304,n28407,n49844 );
   nand U50935 ( n49844,n49845,n49846 );
   nor U50936 ( n49830,n49847,n49848 );
   nand U50937 ( n49848,n49849,n49850 );
   nand U50938 ( n49850,n28286,n49667 );
   xor U50939 ( n49667,n49852,n49853 );
   nand U50940 ( n49849,n49854,n45834 );
   nor U50941 ( n49847,n49855,n49856 );
   nor U50942 ( n49858,n49859,n49860 );
   nand U50943 ( n49860,n49861,n49862 );
   or U50944 ( n49862,n48310,n49842 );
   not U50945 ( n49842,n49863 );
   xor U50946 ( n48310,n49864,n49865 );
   nand U50947 ( n49865,n49866,n49867 );
   nand U50948 ( n49861,n49851,n49672 );
   xor U50949 ( n49672,n49868,n49869 );
   xor U50950 ( n49869,n49870,n49871 );
   nor U50951 ( n49859,n45404,n49872 );
   nor U50952 ( n49857,n49873,n49874 );
   nand U50953 ( n49874,n49875,n49876 );
   nand U50954 ( n49876,n28354,p1_ebx_reg_1_ );
   nor U50955 ( n49875,n49878,n49879 );
   nor U50956 ( n49879,n45674,n49840 );
   nor U50957 ( n49878,p1_reip_reg_1_,n28250 );
   nand U50958 ( n49873,n49880,n49881 );
   nand U50959 ( n49881,n49882,n48317 );
   nand U50960 ( n49880,n28358,p1_phyaddrpointer_reg_1_ );
   nor U50961 ( n49885,n49886,n49887 );
   nand U50962 ( n49887,n49888,n49889 );
   nand U50963 ( n49889,n49854,n46612 );
   nand U50964 ( n49888,n49882,n49890 );
   nand U50965 ( n49886,n49891,n49892 );
   nand U50966 ( n49892,n49863,n48329 );
   nand U50967 ( n48329,n49893,n49894 );
   nand U50968 ( n49894,n49895,n49896 );
   nand U50969 ( n49895,n49897,n49898 );
   or U50970 ( n49893,n49899,n49900 );
   nand U50971 ( n49891,n49851,n49677 );
   xor U50972 ( n49677,n49901,n49902 );
   nor U50973 ( n49884,n49903,n49904 );
   nand U50974 ( n49904,n49905,n49906 );
   nand U50975 ( n49906,n28358,p1_phyaddrpointer_reg_2_ );
   nand U50976 ( n49905,n49877,p1_ebx_reg_2_ );
   nand U50977 ( n49903,n49907,n49908 );
   nand U50978 ( n49908,p1_reip_reg_2_,n49909 );
   nand U50979 ( n49907,n49910,n45669 );
   nor U50980 ( n49910,n45674,n28250 );
   nor U50981 ( n49912,n49913,n49914 );
   nand U50982 ( n49914,n49915,n49916 );
   nand U50983 ( n49916,n49854,n46954 );
   nand U50984 ( n49915,n49882,n48346 );
   nand U50985 ( n49913,n49917,n49918 );
   nand U50986 ( n49918,n48345,n49863 );
   xor U50987 ( n48345,n49919,n49899 );
   nand U50988 ( n49899,n49898,n49920 );
   nand U50989 ( n49920,n49896,n49897 );
   nand U50990 ( n49896,n49866,n49921 );
   nand U50991 ( n49921,n49864,n49867 );
   nand U50992 ( n49864,n49846,n49922 );
   nand U50993 ( n49922,n49843,n49845 );
   nor U50994 ( n49919,n49923,n49924 );
   not U50995 ( n49923,n49925 );
   nand U50996 ( n49917,n49851,n49682 );
   xor U50997 ( n49682,n49926,n49927 );
   nor U50998 ( n49911,n49928,n49929 );
   nand U50999 ( n49929,n49930,n49931 );
   nand U51000 ( n49931,n49883,p1_phyaddrpointer_reg_3_ );
   nand U51001 ( n49930,n28354,p1_ebx_reg_3_ );
   nand U51002 ( n49928,n49932,n49933 );
   nand U51003 ( n49933,p1_reip_reg_3_,n49934 );
   nand U51004 ( n49934,n49935,n49936 );
   nand U51005 ( n49936,n28141,n45669 );
   not U51006 ( n45669,p1_reip_reg_2_ );
   not U51007 ( n49935,n49909 );
   nand U51008 ( n49909,n49840,n49937 );
   nand U51009 ( n49937,n28139,n45674 );
   nand U51010 ( n49932,n49938,n45664 );
   nor U51011 ( n49938,n49841,n49939 );
   nand U51012 ( n49939,p1_reip_reg_2_,p1_reip_reg_1_ );
   nor U51013 ( n49941,n49942,n49943 );
   nand U51014 ( n49943,n49944,n49945 );
   nand U51015 ( n49945,n49851,n49946 );
   not U51016 ( n49946,n47567 );
   nand U51017 ( n47567,n49947,n49948 );
   nand U51018 ( n49947,n49949,n49950 );
   nand U51019 ( n49944,n49854,n47458 );
   not U51020 ( n49854,n49872 );
   nand U51021 ( n49872,n49951,n49952 );
   nand U51022 ( n49942,n49953,n49954 );
   nand U51023 ( n49953,n48359,n49863 );
   xor U51024 ( n48359,n49955,n49956 );
   and U51025 ( n49955,n49957,n49958 );
   nor U51026 ( n49940,n49959,n49960 );
   nand U51027 ( n49960,n49961,n49962 );
   nand U51028 ( n49962,n28354,p1_ebx_reg_4_ );
   nor U51029 ( n49961,n49963,n49964 );
   nor U51030 ( n49964,p1_reip_reg_4_,n49965 );
   nand U51031 ( n49965,n49966,n28141 );
   nor U51032 ( n49963,n49967,n45659 );
   nand U51033 ( n49959,n49968,n49969 );
   nand U51034 ( n49969,n49882,n49970 );
   nand U51035 ( n49968,n49883,p1_phyaddrpointer_reg_4_ );
   nor U51036 ( n49972,n49973,n49974 );
   nand U51037 ( n49974,n49975,n49976 );
   nand U51038 ( n49976,n49851,n49691 );
   xor U51039 ( n49691,n49948,n49977 );
   nand U51040 ( n49975,n49882,n48374 );
   nand U51041 ( n49973,n49978,n49954 );
   nand U51042 ( n49978,n48373,n49863 );
   nand U51043 ( n49863,n49979,n49980 );
   nand U51044 ( n49980,n49952,n45328 );
   xor U51045 ( n48373,n49981,n49982 );
   and U51046 ( n49981,n49983,n49984 );
   nor U51047 ( n49971,n49985,n49986 );
   nand U51048 ( n49986,n49987,n49988 );
   nand U51049 ( n49988,n49883,p1_phyaddrpointer_reg_5_ );
   nand U51050 ( n49987,n28354,p1_ebx_reg_5_ );
   nand U51051 ( n49985,n49989,n49990 );
   nand U51052 ( n49990,p1_reip_reg_5_,n49991 );
   nand U51053 ( n49991,n49967,n49992 );
   nand U51054 ( n49992,n28141,n45659 );
   and U51055 ( n49967,n28220,n49993 );
   nand U51056 ( n49993,n28140,n49994 );
   nand U51057 ( n49989,n49995,n45654 );
   nor U51058 ( n49995,n49994,n49996 );
   nand U51059 ( n49996,n28140,p1_reip_reg_4_ );
   nor U51060 ( n49998,n49999,n50000 );
   nand U51061 ( n50000,n50001,n50002 );
   nand U51062 ( n50002,n49851,n50003 );
   not U51063 ( n50003,n47614 );
   nand U51064 ( n47614,n50004,n50005 );
   nand U51065 ( n50004,n50006,n50007 );
   nand U51066 ( n50001,n49882,n50008 );
   nand U51067 ( n49999,n50009,n49954 );
   nand U51068 ( n50009,n28334,n48387 );
   nand U51069 ( n48387,n50011,n50012 );
   nand U51070 ( n50012,n50013,n50014 );
   or U51071 ( n50011,n50015,n50013 );
   nor U51072 ( n49997,n50016,n50017 );
   nand U51073 ( n50017,n50018,n50019 );
   nand U51074 ( n50019,n49883,p1_phyaddrpointer_reg_6_ );
   nand U51075 ( n50018,n28354,p1_ebx_reg_6_ );
   nand U51076 ( n50016,n50020,n50021 );
   nand U51077 ( n50021,p1_reip_reg_6_,n50022 );
   nand U51078 ( n50020,n50023,n45649 );
   nor U51079 ( n50023,n28250,n50024 );
   nor U51080 ( n50026,n50027,n50028 );
   nand U51081 ( n50028,n50029,n50030 );
   nand U51082 ( n50030,n49851,n49700 );
   xor U51083 ( n49700,n50005,n50031 );
   nand U51084 ( n50029,n49882,n48408 );
   nand U51085 ( n50027,n50032,n49954 );
   nand U51086 ( n50032,n50010,n48407 );
   xor U51087 ( n48407,n50015,n50033 );
   nor U51088 ( n50025,n50034,n50035 );
   nand U51089 ( n50035,n50036,n50037 );
   nand U51090 ( n50037,n49883,p1_phyaddrpointer_reg_7_ );
   nand U51091 ( n50036,n28354,p1_ebx_reg_7_ );
   nand U51092 ( n50034,n50038,n50039 );
   nand U51093 ( n50039,p1_reip_reg_7_,n50040 );
   nand U51094 ( n50040,n50041,n50042 );
   nand U51095 ( n50042,n28139,n45649 );
   not U51096 ( n45649,p1_reip_reg_6_ );
   not U51097 ( n50041,n50022 );
   nand U51098 ( n50022,n49840,n50043 );
   nand U51099 ( n50043,n28139,n50024 );
   nand U51100 ( n50038,n50044,n45644 );
   not U51101 ( n45644,p1_reip_reg_7_ );
   nor U51102 ( n50044,n50024,n50045 );
   nand U51103 ( n50045,n28141,p1_reip_reg_6_ );
   nor U51104 ( n50047,n50048,n50049 );
   nand U51105 ( n50049,n50050,n50051 );
   nand U51106 ( n50051,n49851,n50052 );
   not U51107 ( n50052,n47660 );
   nand U51108 ( n47660,n50053,n50054 );
   nand U51109 ( n50053,n50055,n50056 );
   nand U51110 ( n50050,n49882,n50057 );
   nand U51111 ( n50048,n50058,n49954 );
   nand U51112 ( n50058,n28334,n48423 );
   xor U51113 ( n48423,n50059,n50060 );
   nor U51114 ( n50046,n50061,n50062 );
   nand U51115 ( n50062,n50063,n50064 );
   nand U51116 ( n50064,n49883,p1_phyaddrpointer_reg_8_ );
   nand U51117 ( n50063,n28354,p1_ebx_reg_8_ );
   nand U51118 ( n50061,n50065,n50066 );
   nand U51119 ( n50066,p1_reip_reg_8_,n50067 );
   nand U51120 ( n50065,n50068,n45639 );
   nor U51121 ( n50068,n49841,n50069 );
   nor U51122 ( n50071,n50072,n50073 );
   nand U51123 ( n50073,n50074,n50075 );
   nand U51124 ( n50075,n49851,n49709 );
   xor U51125 ( n49709,n50076,n50054 );
   nand U51126 ( n50074,n49882,n48442 );
   nand U51127 ( n50072,n50077,n49954 );
   nand U51128 ( n50077,n28334,n48441 );
   xor U51129 ( n48441,n50078,n50079 );
   nor U51130 ( n50070,n50080,n50081 );
   nand U51131 ( n50081,n50082,n50083 );
   nand U51132 ( n50083,n49883,p1_phyaddrpointer_reg_9_ );
   nand U51133 ( n50082,n28354,p1_ebx_reg_9_ );
   nand U51134 ( n50080,n50084,n50085 );
   nand U51135 ( n50085,p1_reip_reg_9_,n50086 );
   nand U51136 ( n50086,n50087,n50088 );
   nand U51137 ( n50088,n28141,n45639 );
   not U51138 ( n50087,n50067 );
   nand U51139 ( n50067,n49840,n50089 );
   nand U51140 ( n50089,n28140,n50069 );
   nand U51141 ( n50084,n50090,n45634 );
   nor U51142 ( n50090,n50069,n50091 );
   nand U51143 ( n50091,n28140,p1_reip_reg_8_ );
   not U51144 ( n50069,n50092 );
   nor U51145 ( n50094,n50095,n50096 );
   nand U51146 ( n50096,n50097,n50098 );
   nand U51147 ( n50098,n49851,n50099 );
   not U51148 ( n50099,n47706 );
   nand U51149 ( n47706,n50100,n50101 );
   nand U51150 ( n50100,n50102,n50103 );
   or U51151 ( n50097,n49838,n48457 );
   nand U51152 ( n50095,n50104,n49954 );
   nand U51153 ( n50104,n28334,n48456 );
   nand U51154 ( n48456,n50105,n50106 );
   or U51155 ( n50106,n50107,n50108 );
   nand U51156 ( n50105,n50108,n50109 );
   nor U51157 ( n50093,n50110,n50111 );
   nand U51158 ( n50111,n50112,n50113 );
   nand U51159 ( n50113,n49883,p1_phyaddrpointer_reg_10_ );
   nand U51160 ( n50112,n28354,p1_ebx_reg_10_ );
   nand U51161 ( n50110,n50114,n50115 );
   nand U51162 ( n50115,p1_reip_reg_10_,n50116 );
   nand U51163 ( n50114,n50117,n45629 );
   nor U51164 ( n50117,n28250,n50118 );
   nor U51165 ( n50120,n50121,n50122 );
   nand U51166 ( n50122,n50123,n50124 );
   nand U51167 ( n50124,n49851,n49718 );
   xor U51168 ( n49718,n50125,n50101 );
   nand U51169 ( n50123,n49882,n48478 );
   nand U51170 ( n50121,n50126,n49954 );
   nand U51171 ( n50126,n28334,n48477 );
   not U51172 ( n48477,n49404 );
   xor U51173 ( n49404,n50127,n50107 );
   nand U51174 ( n50107,n50128,n50129 );
   nand U51175 ( n50128,n50130,n50109 );
   nand U51176 ( n50109,n50131,n50132 );
   nand U51177 ( n50132,n50079,n50078 );
   nor U51178 ( n50119,n50133,n50134 );
   nand U51179 ( n50134,n50135,n50136 );
   nand U51180 ( n50136,n49883,p1_phyaddrpointer_reg_11_ );
   nand U51181 ( n50135,n28354,p1_ebx_reg_11_ );
   nand U51182 ( n50133,n50137,n50138 );
   nand U51183 ( n50138,p1_reip_reg_11_,n50139 );
   nand U51184 ( n50139,n50140,n50141 );
   nand U51185 ( n50141,n28139,n45629 );
   not U51186 ( n45629,p1_reip_reg_10_ );
   not U51187 ( n50140,n50116 );
   nand U51188 ( n50116,n49840,n50142 );
   nand U51189 ( n50142,n28139,n50118 );
   nand U51190 ( n50137,n50143,n45624 );
   not U51191 ( n45624,p1_reip_reg_11_ );
   nor U51192 ( n50143,n50118,n50144 );
   nand U51193 ( n50144,n28141,p1_reip_reg_10_ );
   nor U51194 ( n50146,n50147,n50148 );
   nand U51195 ( n50148,n50149,n50150 );
   nand U51196 ( n50150,n49851,n50151 );
   not U51197 ( n50151,n47754 );
   nand U51198 ( n47754,n50152,n50153 );
   nand U51199 ( n50152,n50154,n50155 );
   nand U51200 ( n50149,n49882,n50156 );
   nand U51201 ( n50147,n50157,n49954 );
   nand U51202 ( n50157,n28334,n48492 );
   xor U51203 ( n48492,n50158,n50159 );
   nor U51204 ( n50145,n50160,n50161 );
   nand U51205 ( n50161,n50162,n50163 );
   nand U51206 ( n50163,n49883,p1_phyaddrpointer_reg_12_ );
   nand U51207 ( n50162,n28354,p1_ebx_reg_12_ );
   nand U51208 ( n50160,n50164,n50165 );
   nand U51209 ( n50165,p1_reip_reg_12_,n50166 );
   nand U51210 ( n50164,n50167,n45619 );
   nor U51211 ( n50167,n28250,n50168 );
   nor U51212 ( n50170,n50171,n50172 );
   nand U51213 ( n50172,n50173,n50174 );
   nand U51214 ( n50174,n49851,n49727 );
   xor U51215 ( n49727,n50175,n50153 );
   nand U51216 ( n50173,n49882,n48508 );
   not U51217 ( n49882,n49838 );
   nand U51218 ( n50171,n50176,n49954 );
   nand U51219 ( n50176,n28334,n48507 );
   xor U51220 ( n48507,n50177,n50178 );
   nor U51221 ( n50169,n50179,n50180 );
   nand U51222 ( n50180,n50181,n50182 );
   nand U51223 ( n50182,n49883,p1_phyaddrpointer_reg_13_ );
   nand U51224 ( n50181,n28354,p1_ebx_reg_13_ );
   nand U51225 ( n50179,n50183,n50184 );
   nand U51226 ( n50184,p1_reip_reg_13_,n50185 );
   nand U51227 ( n50185,n50186,n50187 );
   nand U51228 ( n50187,n28141,n45619 );
   not U51229 ( n50186,n50166 );
   nand U51230 ( n50166,n49840,n50188 );
   nand U51231 ( n50188,n28140,n50168 );
   nand U51232 ( n50183,n50189,n45614 );
   nor U51233 ( n50189,n50168,n50190 );
   nand U51234 ( n50190,n28140,p1_reip_reg_12_ );
   not U51235 ( n50168,n50191 );
   nor U51236 ( n50193,n50194,n50195 );
   nand U51237 ( n50195,n50196,n50197 );
   nand U51238 ( n50197,n49851,n50198 );
   not U51239 ( n50198,n47800 );
   nand U51240 ( n47800,n50199,n50200 );
   nand U51241 ( n50199,n50201,n50202 );
   or U51242 ( n50196,n49838,n48523 );
   nand U51243 ( n50194,n50203,n49954 );
   nand U51244 ( n50203,n28334,n48522 );
   nand U51245 ( n48522,n50204,n50205 );
   nand U51246 ( n50205,n50206,n50207 );
   or U51247 ( n50204,n50208,n50206 );
   not U51248 ( n50206,n50209 );
   nor U51249 ( n50192,n50210,n50211 );
   nand U51250 ( n50211,n50212,n50213 );
   nand U51251 ( n50213,n49883,p1_phyaddrpointer_reg_14_ );
   nand U51252 ( n50212,n28354,p1_ebx_reg_14_ );
   nand U51253 ( n50210,n50214,n50215 );
   nand U51254 ( n50215,p1_reip_reg_14_,n50216 );
   nand U51255 ( n50214,n50217,n45609 );
   nor U51256 ( n50217,n49841,n50218 );
   nor U51257 ( n50220,n50221,n50222 );
   nand U51258 ( n50222,n50223,n50224 );
   nand U51259 ( n50224,n49851,n49736 );
   xor U51260 ( n49736,n50225,n50200 );
   or U51261 ( n50223,n49838,n48548 );
   nand U51262 ( n50221,n50226,n49954 );
   nand U51263 ( n50226,n50010,n48547 );
   xor U51264 ( n48547,n50227,n50208 );
   nor U51265 ( n50219,n50228,n50229 );
   nand U51266 ( n50229,n50230,n50231 );
   nand U51267 ( n50231,n49883,p1_phyaddrpointer_reg_15_ );
   nand U51268 ( n50230,n28354,p1_ebx_reg_15_ );
   nand U51269 ( n50228,n50232,n50233 );
   nand U51270 ( n50233,p1_reip_reg_15_,n50234 );
   nand U51271 ( n50234,n50235,n50236 );
   nand U51272 ( n50236,n28139,n45609 );
   not U51273 ( n45609,p1_reip_reg_14_ );
   not U51274 ( n50235,n50216 );
   nand U51275 ( n50216,n49840,n50237 );
   nand U51276 ( n50237,n28139,n50218 );
   nand U51277 ( n50232,n50238,n45604 );
   not U51278 ( n45604,p1_reip_reg_15_ );
   nor U51279 ( n50238,n50218,n50239 );
   nand U51280 ( n50239,n28140,p1_reip_reg_14_ );
   nor U51281 ( n50241,n50242,n50243 );
   nand U51282 ( n50243,n50244,n50245 );
   nand U51283 ( n50245,n28286,n50246 );
   not U51284 ( n50246,n47848 );
   nand U51285 ( n47848,n50247,n50248 );
   nand U51286 ( n50247,n50249,n50250 );
   or U51287 ( n50244,n49838,n48569 );
   nand U51288 ( n50242,n50251,n49954 );
   nand U51289 ( n50251,n50010,n48568 );
   not U51290 ( n48568,n49741 );
   nand U51291 ( n49741,n50252,n50253 );
   nand U51292 ( n50253,n50254,n50255 );
   nor U51293 ( n50240,n50256,n50257 );
   nand U51294 ( n50257,n50258,n50259 );
   nand U51295 ( n50259,n49883,p1_phyaddrpointer_reg_16_ );
   nand U51296 ( n50258,n49877,p1_ebx_reg_16_ );
   nand U51297 ( n50256,n50260,n50261 );
   nand U51298 ( n50261,p1_reip_reg_16_,n50262 );
   nand U51299 ( n50260,n50263,n45599 );
   nor U51300 ( n50263,n28250,n50264 );
   nor U51301 ( n50266,n50267,n50268 );
   nand U51302 ( n50268,n50269,n50270 );
   nand U51303 ( n50270,n28286,n49746 );
   xor U51304 ( n49746,n50271,n50248 );
   or U51305 ( n50269,n49838,n48584 );
   nand U51306 ( n50267,n50272,n49954 );
   nand U51307 ( n50272,n50010,n48583 );
   xor U51308 ( n48583,n50273,n50274 );
   nor U51309 ( n50265,n50275,n50276 );
   nand U51310 ( n50276,n50277,n50278 );
   nand U51311 ( n50278,n49883,p1_phyaddrpointer_reg_17_ );
   nand U51312 ( n50277,n49877,p1_ebx_reg_17_ );
   nand U51313 ( n50275,n50279,n50280 );
   nand U51314 ( n50280,p1_reip_reg_17_,n50281 );
   nand U51315 ( n50281,n50282,n50283 );
   nand U51316 ( n50283,n28140,n45599 );
   not U51317 ( n50282,n50262 );
   nand U51318 ( n50262,n49840,n50284 );
   nand U51319 ( n50284,n28139,n50264 );
   nand U51320 ( n50279,n50285,n45594 );
   nor U51321 ( n50285,n50264,n50286 );
   nand U51322 ( n50286,n28141,p1_reip_reg_16_ );
   not U51323 ( n50264,n50287 );
   nor U51324 ( n50289,n50290,n50291 );
   nand U51325 ( n50291,n50292,n50293 );
   nand U51326 ( n50293,n28286,n50294 );
   not U51327 ( n50294,n47894 );
   nand U51328 ( n47894,n50295,n50296 );
   nand U51329 ( n50295,n50297,n50298 );
   or U51330 ( n50292,n49838,n48602 );
   nand U51331 ( n50290,n50299,n49954 );
   nand U51332 ( n50299,n50010,n48601 );
   xor U51333 ( n48601,n50300,n50301 );
   nor U51334 ( n50288,n50302,n50303 );
   nand U51335 ( n50303,n50304,n50305 );
   nand U51336 ( n50305,n28358,p1_phyaddrpointer_reg_18_ );
   nand U51337 ( n50304,n49877,p1_ebx_reg_18_ );
   nand U51338 ( n50302,n50306,n50307 );
   nand U51339 ( n50307,p1_reip_reg_18_,n50308 );
   nand U51340 ( n50306,n50309,n45589 );
   nor U51341 ( n50309,n28250,n50310 );
   nor U51342 ( n50312,n50313,n50314 );
   nand U51343 ( n50314,n50315,n50316 );
   nand U51344 ( n50316,n28286,n49757 );
   xor U51345 ( n49757,n50317,n50296 );
   or U51346 ( n50315,n49838,n48617 );
   nand U51347 ( n50313,n50318,n49954 );
   nand U51348 ( n49954,n45326,n49840 );
   nand U51349 ( n50318,n50010,n48616 );
   xor U51350 ( n48616,n50319,n50320 );
   nor U51351 ( n50311,n50321,n50322 );
   nand U51352 ( n50322,n50323,n50324 );
   nand U51353 ( n50324,n28358,p1_phyaddrpointer_reg_19_ );
   nand U51354 ( n50323,n49877,p1_ebx_reg_19_ );
   nand U51355 ( n50321,n50325,n50326 );
   nand U51356 ( n50326,p1_reip_reg_19_,n50327 );
   nand U51357 ( n50327,n50328,n50329 );
   nand U51358 ( n50329,n28139,n45589 );
   not U51359 ( n45589,p1_reip_reg_18_ );
   not U51360 ( n50328,n50308 );
   nand U51361 ( n50308,n49840,n50330 );
   nand U51362 ( n50330,n28139,n50310 );
   nand U51363 ( n50325,n50331,n45584 );
   not U51364 ( n45584,p1_reip_reg_19_ );
   nor U51365 ( n50331,n50310,n50332 );
   nand U51366 ( n50332,n28140,p1_reip_reg_18_ );
   nor U51367 ( n50334,n50335,n50336 );
   nand U51368 ( n50336,n50337,n50338 );
   nand U51369 ( n50338,n50010,n48631 );
   xor U51370 ( n48631,n50339,n50340 );
   nand U51371 ( n50337,n28286,n50341 );
   not U51372 ( n50341,n47940 );
   nand U51373 ( n47940,n50342,n50343 );
   nand U51374 ( n50342,n50344,n50345 );
   nor U51375 ( n50335,n48632,n28279 );
   nor U51376 ( n50333,n50346,n50347 );
   nand U51377 ( n50347,n50348,n50349 );
   nand U51378 ( n50349,n28358,p1_phyaddrpointer_reg_20_ );
   nand U51379 ( n50348,n49877,p1_ebx_reg_20_ );
   nand U51380 ( n50346,n50350,n50351 );
   nand U51381 ( n50351,p1_reip_reg_20_,n50352 );
   nand U51382 ( n50350,n50353,n45579 );
   nor U51383 ( n50353,n49841,n50354 );
   nor U51384 ( n50356,n50357,n50358 );
   nand U51385 ( n50358,n50359,n50360 );
   nand U51386 ( n50360,n50010,n48651 );
   xor U51387 ( n48651,n50361,n50362 );
   nand U51388 ( n50359,n28286,n49768 );
   xor U51389 ( n49768,n50363,n50343 );
   nor U51390 ( n50357,n48652,n28279 );
   nor U51391 ( n50355,n50364,n50365 );
   nand U51392 ( n50365,n50366,n50367 );
   nand U51393 ( n50367,n28358,p1_phyaddrpointer_reg_21_ );
   nand U51394 ( n50366,n49877,p1_ebx_reg_21_ );
   nand U51395 ( n50364,n50368,n50369 );
   nand U51396 ( n50369,p1_reip_reg_21_,n50370 );
   nand U51397 ( n50370,n50371,n50372 );
   nand U51398 ( n50372,n28140,n45579 );
   not U51399 ( n50371,n50352 );
   nand U51400 ( n50352,n49840,n50373 );
   nand U51401 ( n50373,n28141,n50354 );
   nand U51402 ( n50368,n50374,n45574 );
   nor U51403 ( n50374,n50354,n50375 );
   nand U51404 ( n50375,n28141,p1_reip_reg_20_ );
   not U51405 ( n50354,n50376 );
   nor U51406 ( n50378,n50379,n50380 );
   nand U51407 ( n50380,n50381,n50382 );
   nand U51408 ( n50382,n50010,n48671 );
   not U51409 ( n48671,n49774 );
   xor U51410 ( n49774,n50383,n50384 );
   nand U51411 ( n50384,n50385,n50386 );
   nor U51412 ( n50383,n50387,n50388 );
   nor U51413 ( n50387,n50361,n50362 );
   and U51414 ( n50361,n50389,n50386 );
   nand U51415 ( n50381,n28286,n50390 );
   not U51416 ( n50390,n47986 );
   nand U51417 ( n47986,n50391,n50392 );
   nand U51418 ( n50391,n50393,n50394 );
   nor U51419 ( n50379,n48672,n28279 );
   nor U51420 ( n50377,n50395,n50396 );
   nand U51421 ( n50396,n50397,n50398 );
   nand U51422 ( n50398,n28358,p1_phyaddrpointer_reg_22_ );
   nand U51423 ( n50397,n49877,p1_ebx_reg_22_ );
   nand U51424 ( n50395,n50399,n50400 );
   nand U51425 ( n50400,p1_reip_reg_22_,n50401 );
   nand U51426 ( n50399,n50402,n45569 );
   nor U51427 ( n50402,n49841,n50403 );
   nor U51428 ( n50405,n50406,n50407 );
   nand U51429 ( n50407,n50408,n50409 );
   nand U51430 ( n50409,n50010,n48690 );
   xor U51431 ( n48690,n50410,n50411 );
   nand U51432 ( n50408,n28286,n49779 );
   xor U51433 ( n49779,n50412,n50392 );
   nor U51434 ( n50406,n48691,n28279 );
   nor U51435 ( n50404,n50413,n50414 );
   nand U51436 ( n50414,n50415,n50416 );
   nand U51437 ( n50416,n28358,p1_phyaddrpointer_reg_23_ );
   nand U51438 ( n50415,n49877,p1_ebx_reg_23_ );
   nand U51439 ( n50413,n50417,n50418 );
   nand U51440 ( n50418,p1_reip_reg_23_,n50419 );
   nand U51441 ( n50419,n50420,n50421 );
   nand U51442 ( n50421,n28139,n45569 );
   not U51443 ( n45569,p1_reip_reg_22_ );
   not U51444 ( n50420,n50401 );
   nand U51445 ( n50401,n49840,n50422 );
   nand U51446 ( n50422,n28139,n50403 );
   nand U51447 ( n50417,n50423,n45564 );
   not U51448 ( n45564,p1_reip_reg_23_ );
   nor U51449 ( n50423,n50403,n50424 );
   nand U51450 ( n50424,n28141,p1_reip_reg_22_ );
   nor U51451 ( n50426,n50427,n50428 );
   nand U51452 ( n50428,n50429,n50430 );
   nand U51453 ( n50430,n50010,n48704 );
   xor U51454 ( n48704,n50431,n50432 );
   nand U51455 ( n50429,n28286,n50433 );
   not U51456 ( n50433,n48032 );
   nand U51457 ( n48032,n50434,n50435 );
   nand U51458 ( n50434,n50436,n50437 );
   nor U51459 ( n50427,n48705,n28279 );
   nor U51460 ( n50425,n50438,n50439 );
   nand U51461 ( n50439,n50440,n50441 );
   nand U51462 ( n50441,n28358,p1_phyaddrpointer_reg_24_ );
   nand U51463 ( n50440,n49877,p1_ebx_reg_24_ );
   nand U51464 ( n50438,n50442,n50443 );
   nand U51465 ( n50443,p1_reip_reg_24_,n50444 );
   nand U51466 ( n50442,n50445,n45559 );
   nor U51467 ( n50445,n49841,n50446 );
   nor U51468 ( n50448,n50449,n50450 );
   nand U51469 ( n50450,n50451,n50452 );
   nand U51470 ( n50452,n50010,n48723 );
   xor U51471 ( n48723,n50453,n50454 );
   nand U51472 ( n50451,n28286,n49790 );
   xor U51473 ( n49790,n50455,n50435 );
   nor U51474 ( n50449,n48724,n28279 );
   nor U51475 ( n50447,n50456,n50457 );
   nand U51476 ( n50457,n50458,n50459 );
   nand U51477 ( n50459,n28358,p1_phyaddrpointer_reg_25_ );
   nand U51478 ( n50458,n49877,p1_ebx_reg_25_ );
   nand U51479 ( n50456,n50460,n50461 );
   nand U51480 ( n50461,p1_reip_reg_25_,n50462 );
   nand U51481 ( n50462,n50463,n50464 );
   nand U51482 ( n50464,n28140,n45559 );
   not U51483 ( n50463,n50444 );
   nand U51484 ( n50444,n49840,n50465 );
   nand U51485 ( n50465,n28141,n50446 );
   nand U51486 ( n50460,n50466,n45554 );
   nor U51487 ( n50466,n50446,n50467 );
   nand U51488 ( n50467,n28141,p1_reip_reg_24_ );
   not U51489 ( n50446,n50468 );
   nor U51490 ( n50470,n50471,n50472 );
   nand U51491 ( n50472,n50473,n50474 );
   nand U51492 ( n50474,n50010,n48738 );
   not U51493 ( n48738,n49796 );
   xor U51494 ( n49796,n50475,n50476 );
   nand U51495 ( n50476,n50477,n50386 );
   nor U51496 ( n50475,n50478,n50479 );
   nor U51497 ( n50478,n50453,n50454 );
   nand U51498 ( n50473,n28286,n50480 );
   not U51499 ( n50480,n48081 );
   nand U51500 ( n48081,n50481,n50482 );
   nand U51501 ( n50481,n50483,n50484 );
   nor U51502 ( n50471,n48739,n49838 );
   nor U51503 ( n50469,n50485,n50486 );
   nand U51504 ( n50486,n50487,n50488 );
   nand U51505 ( n50488,n28358,p1_phyaddrpointer_reg_26_ );
   nand U51506 ( n50487,n49877,p1_ebx_reg_26_ );
   nand U51507 ( n50485,n50489,n50490 );
   nand U51508 ( n50490,p1_reip_reg_26_,n50491 );
   nand U51509 ( n50489,n50492,n45549 );
   nor U51510 ( n50492,n28250,n50493 );
   nor U51511 ( n50495,n50496,n50497 );
   nand U51512 ( n50497,n50498,n50499 );
   nand U51513 ( n50499,n50010,n48761 );
   not U51514 ( n48761,n49802 );
   xor U51515 ( n49802,n50500,n50501 );
   nor U51516 ( n50500,n50479,n50502 );
   nand U51517 ( n50498,n28286,n49801 );
   xor U51518 ( n49801,n50503,n50482 );
   nor U51519 ( n50496,n48762,n28279 );
   nor U51520 ( n50494,n50504,n50505 );
   nand U51521 ( n50505,n50506,n50507 );
   nand U51522 ( n50507,n28358,p1_phyaddrpointer_reg_27_ );
   nand U51523 ( n50506,n49877,p1_ebx_reg_27_ );
   nand U51524 ( n50504,n50508,n50509 );
   nand U51525 ( n50509,p1_reip_reg_27_,n50510 );
   nand U51526 ( n50510,n50511,n50512 );
   nand U51527 ( n50512,n28139,n45549 );
   not U51528 ( n45549,p1_reip_reg_26_ );
   not U51529 ( n50511,n50491 );
   nand U51530 ( n50491,n49840,n50513 );
   nand U51531 ( n50513,n28139,n50493 );
   nand U51532 ( n50508,n50514,n45544 );
   not U51533 ( n45544,p1_reip_reg_27_ );
   nor U51534 ( n50514,n50493,n50515 );
   nand U51535 ( n50515,n28140,p1_reip_reg_26_ );
   nor U51536 ( n50517,n50518,n50519 );
   nand U51537 ( n50519,n50520,n50521 );
   nand U51538 ( n50521,n50010,n48783 );
   xor U51539 ( n48783,n50522,n50523 );
   nand U51540 ( n50520,n28286,n50524 );
   not U51541 ( n50524,n48124 );
   nand U51542 ( n48124,n50525,n50526 );
   nand U51543 ( n50525,n50527,n50528 );
   nor U51544 ( n50518,n48784,n28279 );
   nor U51545 ( n50516,n50529,n50530 );
   nand U51546 ( n50530,n50531,n50532 );
   nand U51547 ( n50532,n28358,p1_phyaddrpointer_reg_28_ );
   nand U51548 ( n50531,n49877,p1_ebx_reg_28_ );
   nand U51549 ( n50529,n50533,n50534 );
   nand U51550 ( n50534,p1_reip_reg_28_,n50535 );
   nand U51551 ( n50533,n50536,n45539 );
   nor U51552 ( n50536,n49841,n50537 );
   nor U51553 ( n50539,n50540,n50541 );
   nand U51554 ( n50541,n50542,n50543 );
   nand U51555 ( n50543,n50010,n48798 );
   xor U51556 ( n48798,n50544,n50545 );
   nand U51557 ( n50542,n28286,n49812 );
   xor U51558 ( n49812,n50546,n50526 );
   nor U51559 ( n50540,n48799,n28279 );
   nor U51560 ( n50538,n50547,n50548 );
   nand U51561 ( n50548,n50549,n50550 );
   nand U51562 ( n50550,n28358,p1_phyaddrpointer_reg_29_ );
   nand U51563 ( n50549,n49877,p1_ebx_reg_29_ );
   nand U51564 ( n50547,n50551,n50552 );
   or U51565 ( n50552,n50553,p1_reip_reg_29_ );
   or U51566 ( n50551,n45534,n50554 );
   nor U51567 ( n50556,n50557,n50558 );
   nand U51568 ( n50558,n50559,n50560 );
   nand U51569 ( n50560,n50010,n48824 );
   xor U51570 ( n48824,n50561,n50562 );
   nand U51571 ( n50559,n28286,n49819 );
   xor U51572 ( n49819,n50563,n50564 );
   nor U51573 ( n50557,n48825,n28279 );
   nand U51574 ( n49838,n50565,n49010 );
   nor U51575 ( n50565,n50566,n45432 );
   nor U51576 ( n50555,n50567,n50568 );
   nand U51577 ( n50568,n50569,n50570 );
   nand U51578 ( n50570,n28358,p1_phyaddrpointer_reg_30_ );
   nand U51579 ( n50569,n28354,p1_ebx_reg_30_ );
   not U51580 ( n49877,n49856 );
   nand U51581 ( n50567,n50571,n50572 );
   nand U51582 ( n50572,p1_reip_reg_30_,n50573 );
   nand U51583 ( n50571,n50574,n45529 );
   nor U51584 ( n50574,n45534,n50553 );
   nor U51585 ( n50576,n50577,n50578 );
   nand U51586 ( n50578,n50579,n50580 );
   nand U51587 ( n50580,n28334,n48835 );
   and U51588 ( n48835,n50581,n50582 );
   nand U51589 ( n50582,n50583,n50584 );
   nand U51590 ( n50584,n50562,n50561 );
   nand U51591 ( n50562,n50585,n50586 );
   nand U51592 ( n50585,n50587,n50588 );
   not U51593 ( n50583,n50589 );
   nand U51594 ( n50581,n50590,n50589 );
   nand U51595 ( n50589,n50591,n50592 );
   nand U51596 ( n50592,p1_phyaddrpointer_reg_31_,n49013 );
   nand U51597 ( n50591,p1_eax_reg_31_,n50593 );
   nor U51598 ( n50590,n50594,n50586 );
   nand U51599 ( n50586,n50545,n50544 );
   nand U51600 ( n50544,n50595,n50386 );
   xor U51601 ( n50595,n50587,n28184 );
   nand U51602 ( n50587,n50596,n50597 );
   nor U51603 ( n50597,n50598,n50599 );
   nor U51604 ( n50599,n28182,n48799 );
   nand U51605 ( n48799,n50600,n50601 );
   nand U51606 ( n50601,n50602,n48802 );
   nor U51607 ( n50598,n50603,n28241 );
   xor U51608 ( n50603,n50605,n50606 );
   nor U51609 ( n50596,n50607,n50608 );
   nor U51610 ( n50608,n28288,n49322 );
   not U51611 ( n49322,p1_eax_reg_29_ );
   nor U51612 ( n50607,n28251,n48802 );
   nand U51613 ( n50545,n50611,n50612 );
   nand U51614 ( n50612,n50522,n50523 );
   nand U51615 ( n50523,n50613,n50386 );
   xor U51616 ( n50613,n50614,n28184 );
   nand U51617 ( n50522,n50615,n50616 );
   nand U51618 ( n50616,n50502,n50501 );
   nand U51619 ( n50501,n50617,n50386 );
   nor U51620 ( n50502,n50618,n50454 );
   nand U51621 ( n50454,n50431,n50432 );
   nand U51622 ( n50432,n50619,n50386 );
   not U51623 ( n50619,n50620 );
   and U51624 ( n50431,n50410,n50411 );
   nand U51625 ( n50411,n50621,n50622 );
   nand U51626 ( n50622,n50623,n50588 );
   nand U51627 ( n50623,n50385,n50362 );
   nor U51628 ( n50621,n50388,n50624 );
   nor U51629 ( n50624,n50389,n50625 );
   or U51630 ( n50625,n50385,n50362 );
   nand U51631 ( n50362,n50339,n50340 );
   nand U51632 ( n50340,n50626,n50386 );
   and U51633 ( n50339,n50320,n50319 );
   nand U51634 ( n50319,n50627,n50628 );
   nand U51635 ( n50628,n50629,n50588 );
   nand U51636 ( n50629,n50630,n50631 );
   nand U51637 ( n50627,n50301,n50300 );
   nand U51638 ( n50300,n50630,n50386 );
   xor U51639 ( n50630,n28183,n50632 );
   nand U51640 ( n50632,n50633,n50634 );
   nor U51641 ( n50634,n50635,n50636 );
   nor U51642 ( n50636,n28182,n48602 );
   nand U51643 ( n48602,n50637,n50638 );
   nand U51644 ( n50637,n48605,n50639 );
   nand U51645 ( n50639,n50640,p1_phyaddrpointer_reg_17_ );
   nor U51646 ( n50635,n50641,n50642 );
   nor U51647 ( n50641,n50643,n50644 );
   nand U51648 ( n50644,n50645,n50646 );
   nor U51649 ( n50646,n50647,n50648 );
   nand U51650 ( n50648,n50649,n50650 );
   nand U51651 ( n50650,n50651,p1_instqueue_reg_7__2_ );
   nand U51652 ( n50649,n50652,p1_instqueue_reg_6__2_ );
   nand U51653 ( n50647,n50653,n50654 );
   nand U51654 ( n50654,n50655,p1_instqueue_reg_5__2_ );
   nand U51655 ( n50653,n50656,p1_instqueue_reg_4__2_ );
   nor U51656 ( n50645,n50657,n50658 );
   nand U51657 ( n50658,n50659,n50660 );
   nand U51658 ( n50660,n50661,p1_instqueue_reg_3__2_ );
   nand U51659 ( n50659,n50662,p1_instqueue_reg_2__2_ );
   nand U51660 ( n50657,n50663,n50664 );
   nand U51661 ( n50664,n50665,p1_instqueue_reg_1__2_ );
   nand U51662 ( n50663,n50666,p1_instqueue_reg_0__2_ );
   nand U51663 ( n50643,n50667,n50668 );
   nor U51664 ( n50668,n50669,n50670 );
   nand U51665 ( n50670,n50671,n50672 );
   nand U51666 ( n50672,n50673,p1_instqueue_reg_15__2_ );
   nand U51667 ( n50671,n50674,p1_instqueue_reg_14__2_ );
   nand U51668 ( n50669,n50675,n50676 );
   nand U51669 ( n50676,n50677,p1_instqueue_reg_13__2_ );
   nand U51670 ( n50675,n50678,p1_instqueue_reg_12__2_ );
   nor U51671 ( n50667,n50679,n50680 );
   nand U51672 ( n50680,n50681,n50682 );
   nand U51673 ( n50682,n50683,p1_instqueue_reg_11__2_ );
   nand U51674 ( n50681,n50684,p1_instqueue_reg_10__2_ );
   nand U51675 ( n50679,n50685,n50686 );
   nand U51676 ( n50686,n50687,p1_instqueue_reg_9__2_ );
   nand U51677 ( n50685,n50688,p1_instqueue_reg_8__2_ );
   nor U51678 ( n50633,n50689,n50690 );
   nor U51679 ( n50690,n50609,n49267 );
   not U51680 ( n49267,p1_eax_reg_18_ );
   nor U51681 ( n50689,n50610,n48605 );
   not U51682 ( n48605,p1_phyaddrpointer_reg_18_ );
   and U51683 ( n50301,n50274,n50273 );
   nand U51684 ( n50273,n50631,n50386 );
   xor U51685 ( n50631,n28183,n50691 );
   nand U51686 ( n50691,n50692,n50693 );
   nor U51687 ( n50693,n50694,n50695 );
   nor U51688 ( n50695,n48584,n28182 );
   xor U51689 ( n48584,n48587,n50640 );
   nor U51690 ( n50694,n50696,n50642 );
   nor U51691 ( n50696,n50697,n50698 );
   nand U51692 ( n50698,n50699,n50700 );
   nor U51693 ( n50700,n50701,n50702 );
   nand U51694 ( n50702,n50703,n50704 );
   nand U51695 ( n50704,n50651,p1_instqueue_reg_7__1_ );
   nand U51696 ( n50703,n50652,p1_instqueue_reg_6__1_ );
   nand U51697 ( n50701,n50705,n50706 );
   nand U51698 ( n50706,n50655,p1_instqueue_reg_5__1_ );
   nand U51699 ( n50705,n50656,p1_instqueue_reg_4__1_ );
   nor U51700 ( n50699,n50707,n50708 );
   nand U51701 ( n50708,n50709,n50710 );
   nand U51702 ( n50710,n50661,p1_instqueue_reg_3__1_ );
   nand U51703 ( n50709,n50662,p1_instqueue_reg_2__1_ );
   nand U51704 ( n50707,n50711,n50712 );
   nand U51705 ( n50712,n50665,p1_instqueue_reg_1__1_ );
   nand U51706 ( n50711,n50666,p1_instqueue_reg_0__1_ );
   nand U51707 ( n50697,n50713,n50714 );
   nor U51708 ( n50714,n50715,n50716 );
   nand U51709 ( n50716,n50717,n50718 );
   nand U51710 ( n50718,n50673,p1_instqueue_reg_15__1_ );
   nand U51711 ( n50717,n50674,p1_instqueue_reg_14__1_ );
   nand U51712 ( n50715,n50719,n50720 );
   nand U51713 ( n50720,n50677,p1_instqueue_reg_13__1_ );
   nand U51714 ( n50719,n50678,p1_instqueue_reg_12__1_ );
   nor U51715 ( n50713,n50721,n50722 );
   nand U51716 ( n50722,n50723,n50724 );
   nand U51717 ( n50724,n50683,p1_instqueue_reg_11__1_ );
   nand U51718 ( n50723,n50684,p1_instqueue_reg_10__1_ );
   nand U51719 ( n50721,n50725,n50726 );
   nand U51720 ( n50726,n50687,p1_instqueue_reg_9__1_ );
   nand U51721 ( n50725,n50688,p1_instqueue_reg_8__1_ );
   nor U51722 ( n50692,n50727,n50728 );
   nor U51723 ( n50728,n28288,n49262 );
   not U51724 ( n49262,p1_eax_reg_17_ );
   nor U51725 ( n50727,n28252,n48587 );
   nand U51726 ( n50274,n50729,n50252 );
   or U51727 ( n50252,n50255,n50254 );
   and U51728 ( n50254,n50730,n50731 );
   nand U51729 ( n50731,n50732,n50733 );
   not U51730 ( n50732,n50734 );
   nand U51731 ( n50730,n50208,n50227 );
   nand U51732 ( n50227,n50735,n50734 );
   nand U51733 ( n50734,n50736,n28262 );
   xor U51734 ( n50736,n48875,n48876 );
   xor U51735 ( n50735,n50733,n28185 );
   nand U51736 ( n50733,n50738,n50739 );
   nand U51737 ( n50739,p1_eax_reg_15_,n50593 );
   nor U51738 ( n50738,n50740,n50741 );
   nor U51739 ( n50741,n28252,n48551 );
   nor U51740 ( n50740,n28185,n48548 );
   nand U51741 ( n48548,n50742,n50743 );
   nand U51742 ( n50743,n50744,n48551 );
   nand U51743 ( n50208,n50745,n50746 );
   nand U51744 ( n50746,n50747,n28262 );
   nor U51745 ( n50747,n50748,n50749 );
   not U51746 ( n50749,n48877 );
   nand U51747 ( n50745,n50207,n50209 );
   nand U51748 ( n50209,n50750,n50751 );
   nand U51749 ( n50751,n50737,n48877 );
   nor U51750 ( n48877,n48875,n50752 );
   and U51751 ( n50752,n50753,n50754 );
   xor U51752 ( n50750,n50748,n49843 );
   and U51753 ( n50748,n50755,n50756 );
   nand U51754 ( n50756,p1_eax_reg_14_,n50593 );
   nor U51755 ( n50755,n50757,n50758 );
   nor U51756 ( n50758,n28252,n48526 );
   nor U51757 ( n50757,n28184,n48523 );
   nand U51758 ( n48523,n50744,n50759 );
   nand U51759 ( n50759,n50760,n48526 );
   not U51760 ( n48526,p1_phyaddrpointer_reg_14_ );
   or U51761 ( n50760,n50761,n48511 );
   nand U51762 ( n50207,n50762,n50763 );
   nand U51763 ( n50763,n50764,n50765 );
   nand U51764 ( n50762,n50178,n50177 );
   or U51765 ( n50177,n50765,n50764 );
   and U51766 ( n50764,n50737,n48869 );
   and U51767 ( n48869,n50754,n50766 );
   nand U51768 ( n50766,n50767,n50768 );
   xor U51769 ( n50765,n50769,n28182 );
   nor U51770 ( n50769,n50770,n50771 );
   nand U51771 ( n50771,n50772,n50773 );
   nand U51772 ( n50773,n28408,n48508 );
   xor U51773 ( n48508,n48511,n50761 );
   nand U51774 ( n50772,p1_phyaddrpointer_reg_13_,n49013 );
   nor U51775 ( n50770,n28287,n49243 );
   not U51776 ( n49243,p1_eax_reg_13_ );
   nand U51777 ( n50178,n50774,n50775 );
   nand U51778 ( n50775,n50776,n50777 );
   not U51779 ( n50777,n50778 );
   nor U51780 ( n50776,n48864,n50604 );
   nand U51781 ( n50774,n50158,n50159 );
   nand U51782 ( n50159,n50778,n50779 );
   nand U51783 ( n50779,n50737,n48985 );
   not U51784 ( n48985,n48864 );
   nand U51785 ( n48864,n50780,n50768 );
   nand U51786 ( n50780,n50781,n50782 );
   nand U51787 ( n50782,n50783,n50784 );
   xor U51788 ( n50778,n50785,n49843 );
   nor U51789 ( n50785,n50786,n50787 );
   nand U51790 ( n50787,n50788,n50789 );
   nand U51791 ( n50789,n50156,n49843 );
   not U51792 ( n50156,n48493 );
   nand U51793 ( n48493,n50790,n50761 );
   nand U51794 ( n50790,n48496,n50791 );
   or U51795 ( n50791,n50792,n48481 );
   not U51796 ( n48496,p1_phyaddrpointer_reg_12_ );
   nand U51797 ( n50788,p1_phyaddrpointer_reg_12_,n49013 );
   nor U51798 ( n50786,n50609,n49238 );
   not U51799 ( n49238,p1_eax_reg_12_ );
   nand U51800 ( n50158,n50793,n50794 );
   nand U51801 ( n50794,n50795,n50796 );
   nand U51802 ( n50796,n50129,n50797 );
   nand U51803 ( n50797,n50798,n50078 );
   nand U51804 ( n50078,n50799,n50800 );
   nand U51805 ( n50800,n28262,n48885 );
   nand U51806 ( n50798,n50801,n50131 );
   nand U51807 ( n50131,n50802,n50803 );
   not U51808 ( n50803,n50799 );
   xor U51809 ( n50799,n50804,n49843 );
   nor U51810 ( n50804,n50805,n50806 );
   nand U51811 ( n50806,n50807,n50808 );
   nand U51812 ( n50808,n28407,n48442 );
   xor U51813 ( n48442,n48445,n50809 );
   nand U51814 ( n50807,p1_phyaddrpointer_reg_9_,n49013 );
   nor U51815 ( n50805,n28288,n49224 );
   not U51816 ( n49224,p1_eax_reg_9_ );
   nor U51817 ( n50802,n50604,n48888 );
   not U51818 ( n48888,n48885 );
   xor U51819 ( n48885,n50810,n50811 );
   not U51820 ( n50801,n50079 );
   nand U51821 ( n50079,n50812,n50813 );
   nand U51822 ( n50813,n50814,n50815 );
   nand U51823 ( n50812,n50060,n50059 );
   or U51824 ( n50059,n50815,n50814 );
   and U51825 ( n50814,n50816,n28262 );
   nor U51826 ( n50816,n50811,n50817 );
   nor U51827 ( n50817,n48970,n48969 );
   xor U51828 ( n50815,n50818,n28185 );
   nor U51829 ( n50818,n50819,n50820 );
   nand U51830 ( n50820,n50821,n50822 );
   nand U51831 ( n50822,n50057,n28408 );
   not U51832 ( n50057,n48424 );
   nand U51833 ( n48424,n50823,n50809 );
   nand U51834 ( n50823,n48427,n50824 );
   or U51835 ( n50824,n50825,n48411 );
   not U51836 ( n48427,p1_phyaddrpointer_reg_8_ );
   nand U51837 ( n50821,p1_phyaddrpointer_reg_8_,n49013 );
   nor U51838 ( n50819,n28287,n49219 );
   not U51839 ( n49219,p1_eax_reg_8_ );
   nand U51840 ( n50060,n50826,n50827 );
   nand U51841 ( n50827,n50015,n50033 );
   nand U51842 ( n50033,n50828,n50829 );
   nor U51843 ( n50015,n50013,n50830 );
   nor U51844 ( n50830,n50014,n50831 );
   and U51845 ( n50831,n50832,n28262 );
   and U51846 ( n50832,n50833,n48956 );
   nand U51847 ( n50014,n49983,n50834 );
   nand U51848 ( n50834,n49984,n49982 );
   nand U51849 ( n49982,n49957,n50835 );
   nand U51850 ( n50835,n49958,n49956 );
   nand U51851 ( n49956,n49925,n50836 );
   nand U51852 ( n50836,n50837,n50838 );
   nand U51853 ( n50838,n50839,n50840 );
   nand U51854 ( n50840,n50841,n50842 );
   nand U51855 ( n50842,n28185,n49846 );
   nand U51856 ( n49846,n50843,n50844 );
   and U51857 ( n50841,n49845,n49867 );
   nand U51858 ( n49867,n50845,n50846 );
   or U51859 ( n49845,n50844,n50843 );
   and U51860 ( n50843,p1_state2_reg_2_,n50847 );
   nand U51861 ( n50847,n47130,n48218 );
   not U51862 ( n47130,n45389 );
   nand U51863 ( n45389,n50848,n50849 );
   nand U51864 ( n50849,n48996,n50850 );
   nand U51865 ( n50848,n50851,n50852 );
   nand U51866 ( n50852,n50853,n50854 );
   nor U51867 ( n50854,n50855,n50856 );
   nor U51868 ( n50855,n47364,n48270 );
   nor U51869 ( n50853,n28094,n50857 );
   xor U51870 ( n50844,n28408,n50858 );
   nand U51871 ( n50858,n50859,n50860 );
   nor U51872 ( n50860,n50861,n50862 );
   nor U51873 ( n50862,n28287,n49179 );
   not U51874 ( n49179,p1_eax_reg_0_ );
   nor U51875 ( n50861,n45394,n50604 );
   nor U51876 ( n50859,n50863,n50864 );
   nor U51877 ( n50864,n50865,n48295 );
   not U51878 ( n48295,p1_phyaddrpointer_reg_0_ );
   nor U51879 ( n50865,n28407,n49013 );
   nor U51880 ( n50863,n45451,n50866 );
   and U51881 ( n50839,n49866,n49898 );
   nand U51882 ( n49898,n50867,n50868 );
   nand U51883 ( n50868,n50869,n28251 );
   nand U51884 ( n50869,n28262,n45414 );
   or U51885 ( n49866,n50846,n50845 );
   xor U51886 ( n50845,n50870,n28407 );
   nor U51887 ( n50870,n50871,n50872 );
   nand U51888 ( n50872,n50873,n50874 );
   nand U51889 ( n50874,n48249,p1_instqueuerd_addr_reg_1_ );
   nor U51890 ( n50873,n50875,n50876 );
   nor U51891 ( n50876,n28251,n48317 );
   nor U51892 ( n50875,p1_phyaddrpointer_reg_1_,n28185 );
   nand U51893 ( n50871,n50877,n50878 );
   nand U51894 ( n50878,n50737,n46090 );
   nand U51895 ( n50877,p1_eax_reg_1_,n50593 );
   nand U51896 ( n50846,n50737,n45401 );
   xor U51897 ( n45401,n50851,n50879 );
   nand U51898 ( n50879,n50880,n50881 );
   nor U51899 ( n50837,n49924,n49900 );
   not U51900 ( n49900,n49897 );
   nand U51901 ( n49897,n50882,n50883 );
   xor U51902 ( n50883,n50867,n28184 );
   nand U51903 ( n50867,n50884,n50885 );
   nor U51904 ( n50885,n50886,n50887 );
   nand U51905 ( n50887,n50888,n50889 );
   nand U51906 ( n50889,n49890,n49843 );
   not U51907 ( n49890,n48331 );
   nand U51908 ( n48331,n50890,n50891 );
   nand U51909 ( n50891,n48317,n48335 );
   not U51910 ( n48317,p1_phyaddrpointer_reg_1_ );
   nand U51911 ( n50888,n50737,n46612 );
   nor U51912 ( n50886,n28252,n48335 );
   not U51913 ( n48335,p1_phyaddrpointer_reg_2_ );
   nor U51914 ( n50884,n50892,n50893 );
   nor U51915 ( n50893,n47402,n50866 );
   nor U51916 ( n50892,n50609,n49190 );
   not U51917 ( n49190,p1_eax_reg_2_ );
   nor U51918 ( n50882,n49013,n50894 );
   nor U51919 ( n50894,n46269,n28241 );
   not U51920 ( n46269,n45414 );
   nand U51921 ( n45414,n50895,n50896 );
   nand U51922 ( n50896,n50897,n50898 );
   nand U51923 ( n50898,n50899,n50900 );
   nand U51924 ( n50895,n50901,n50899 );
   nor U51925 ( n49924,n50902,n50903 );
   xor U51926 ( n50902,n50904,n28407 );
   nand U51927 ( n49925,n50903,n50904 );
   nand U51928 ( n50904,n50905,n50906 );
   nor U51929 ( n50906,n50907,n50908 );
   nand U51930 ( n50908,n50909,n50910 );
   nand U51931 ( n50910,n28408,n48346 );
   xor U51932 ( n48346,n48349,n50890 );
   nand U51933 ( n50909,n50737,n46954 );
   nor U51934 ( n50907,n28251,n48349 );
   nor U51935 ( n50905,n50911,n50912 );
   nor U51936 ( n50912,n50913,n50866 );
   not U51937 ( n50866,n48249 );
   nor U51938 ( n50911,n28288,n49195 );
   not U51939 ( n49195,p1_eax_reg_3_ );
   nor U51940 ( n50903,n50604,n46268 );
   not U51941 ( n46268,n45428 );
   xor U51942 ( n45428,n50914,n50915 );
   nand U51943 ( n50915,n50916,n50917 );
   nor U51944 ( n50914,n50918,n50919 );
   nor U51945 ( n50918,n50920,n50921 );
   nand U51946 ( n49958,n50922,n50923 );
   or U51947 ( n49957,n50923,n50922 );
   xor U51948 ( n50922,n28183,n50924 );
   nand U51949 ( n50924,n50925,n50926 );
   nor U51950 ( n50926,n50927,n50928 );
   nand U51951 ( n50928,n50929,n50930 );
   nand U51952 ( n50930,n49970,n28407 );
   not U51953 ( n49970,n48360 );
   nand U51954 ( n48360,n50931,n50932 );
   nand U51955 ( n50931,n48363,n50933 );
   or U51956 ( n50933,n50890,n48349 );
   nand U51957 ( n50929,n50737,n47458 );
   xor U51958 ( n47458,n50934,n50935 );
   nand U51959 ( n50935,n50936,n50937 );
   nor U51960 ( n50927,n50610,n48363 );
   not U51961 ( n48363,p1_phyaddrpointer_reg_4_ );
   nor U51962 ( n50925,n50938,n50939 );
   and U51963 ( n50939,p1_instqueuerd_addr_reg_4_,n48249 );
   nor U51964 ( n50938,n28287,n49200 );
   not U51965 ( n49200,p1_eax_reg_4_ );
   nand U51966 ( n50923,n50737,n48917 );
   xor U51967 ( n48917,n50940,n50941 );
   nand U51968 ( n50941,n50942,n50943 );
   not U51969 ( n50940,n50944 );
   nand U51970 ( n49984,n50945,n50946 );
   or U51971 ( n49983,n50946,n50945 );
   xor U51972 ( n50945,n50947,n28408 );
   nor U51973 ( n50947,n50948,n50949 );
   nand U51974 ( n50949,n50950,n50951 );
   nand U51975 ( n50951,p1_phyaddrpointer_reg_5_,n49013 );
   nand U51976 ( n50950,p1_eax_reg_5_,n50593 );
   nand U51977 ( n50948,n50952,n50953 );
   nand U51978 ( n50953,n50954,n50955 );
   and U51979 ( n50955,n50937,n50936 );
   nor U51980 ( n50954,n50934,n28241 );
   nand U51981 ( n50934,p1_instqueuerd_addr_reg_4_,n50956 );
   nand U51982 ( n50956,n45836,n47429 );
   nand U51983 ( n50952,n28407,n48374 );
   xor U51984 ( n48374,n48377,n50932 );
   nand U51985 ( n50946,n50737,n48905 );
   nand U51986 ( n48905,n50957,n50958 );
   nand U51987 ( n50958,n50959,n50960 );
   nand U51988 ( n50959,n50961,n50962 );
   nand U51989 ( n50957,n50963,n50961 );
   and U51990 ( n50013,n50964,n50965 );
   nand U51991 ( n50965,n50737,n48956 );
   xor U51992 ( n48956,n50966,n50967 );
   and U51993 ( n50966,n50968,n50969 );
   xor U51994 ( n50964,n50833,n28182 );
   nand U51995 ( n50833,n50970,n50971 );
   nand U51996 ( n50971,n50008,n28408 );
   not U51997 ( n50008,n48388 );
   nand U51998 ( n48388,n50825,n50972 );
   nand U51999 ( n50972,n50973,n48391 );
   or U52000 ( n50973,n50932,n48377 );
   nor U52001 ( n50970,n50974,n50975 );
   nor U52002 ( n50975,n28251,n48391 );
   not U52003 ( n48391,p1_phyaddrpointer_reg_6_ );
   nor U52004 ( n50974,n50609,n49209 );
   not U52005 ( n49209,p1_eax_reg_6_ );
   or U52006 ( n50826,n50829,n50828 );
   xor U52007 ( n50828,n50976,n28408 );
   nor U52008 ( n50976,n50977,n50978 );
   nand U52009 ( n50978,n50979,n50980 );
   nand U52010 ( n50980,n28408,n48408 );
   xor U52011 ( n48408,n48411,n50825 );
   nand U52012 ( n50979,p1_phyaddrpointer_reg_7_,n49013 );
   nor U52013 ( n50977,n28288,n49214 );
   not U52014 ( n49214,p1_eax_reg_7_ );
   nand U52015 ( n50829,n50981,n48974 );
   nor U52016 ( n48974,n50982,n50983 );
   nor U52017 ( n50983,n50969,n50984 );
   and U52018 ( n50982,n50985,n50986 );
   and U52019 ( n50986,n50968,n50961 );
   nor U52020 ( n50985,n50963,n50984 );
   nor U52021 ( n50963,n50960,n50987 );
   nor U52022 ( n50981,n48975,n28241 );
   nand U52023 ( n48975,n50988,n50989 );
   nand U52024 ( n50989,n50990,n50991 );
   not U52025 ( n50991,n50967 );
   and U52026 ( n50990,n50969,n50984 );
   nand U52027 ( n50988,n50992,n50984 );
   nand U52028 ( n50984,n50993,n50994 );
   nand U52029 ( n50129,n50995,n28262 );
   nor U52030 ( n50995,n50996,n48882 );
   nor U52031 ( n50795,n50108,n50127 );
   nor U52032 ( n50127,n50997,n50998 );
   not U52033 ( n50108,n50130 );
   nand U52034 ( n50130,n50999,n51000 );
   or U52035 ( n51000,n50604,n48882 );
   nand U52036 ( n48882,n51001,n51002 );
   nand U52037 ( n51002,n51003,n51004 );
   not U52038 ( n51001,n50783 );
   xor U52039 ( n50999,n28407,n50996 );
   and U52040 ( n50996,n51005,n51006 );
   nand U52041 ( n51006,p1_eax_reg_10_,n50593 );
   nor U52042 ( n51005,n51007,n51008 );
   nor U52043 ( n51008,n50610,n48460 );
   nor U52044 ( n51007,n28185,n48457 );
   nand U52045 ( n48457,n50792,n51009 );
   nand U52046 ( n51009,n51010,n48460 );
   not U52047 ( n48460,p1_phyaddrpointer_reg_10_ );
   or U52048 ( n51010,n50809,n48445 );
   nand U52049 ( n50793,n50998,n50997 );
   xor U52050 ( n50997,n51011,n28182 );
   nor U52051 ( n51011,n51012,n51013 );
   nand U52052 ( n51013,n51014,n51015 );
   nand U52053 ( n51015,n49843,n48478 );
   xor U52054 ( n48478,n48481,n50792 );
   nand U52055 ( n51014,p1_phyaddrpointer_reg_11_,n49013 );
   nor U52056 ( n51012,n28287,n49233 );
   not U52057 ( n49233,p1_eax_reg_11_ );
   nor U52058 ( n50998,n50604,n48983 );
   xor U52059 ( n48983,n51016,n50783 );
   nor U52060 ( n50255,n51017,n50588 );
   nand U52061 ( n50729,n51017,n50588 );
   xor U52062 ( n51017,n49843,n51018 );
   nand U52063 ( n51018,n51019,n51020 );
   nor U52064 ( n51020,n51021,n51022 );
   nor U52065 ( n51022,n28184,n48569 );
   nand U52066 ( n48569,n51023,n51024 );
   nand U52067 ( n51023,n48572,n50742 );
   nor U52068 ( n51021,n51025,n50642 );
   nor U52069 ( n51025,n51026,n51027 );
   nand U52070 ( n51027,n51028,n51029 );
   nor U52071 ( n51029,n51030,n51031 );
   nand U52072 ( n51031,n51032,n51033 );
   nand U52073 ( n51033,n50651,p1_instqueue_reg_7__0_ );
   nand U52074 ( n51032,n50652,p1_instqueue_reg_6__0_ );
   nand U52075 ( n51030,n51034,n51035 );
   nand U52076 ( n51035,n50655,p1_instqueue_reg_5__0_ );
   nand U52077 ( n51034,n50656,p1_instqueue_reg_4__0_ );
   nor U52078 ( n51028,n51036,n51037 );
   nand U52079 ( n51037,n51038,n51039 );
   nand U52080 ( n51039,n50661,p1_instqueue_reg_3__0_ );
   nand U52081 ( n51038,n50662,p1_instqueue_reg_2__0_ );
   nand U52082 ( n51036,n51040,n51041 );
   nand U52083 ( n51041,n50665,p1_instqueue_reg_1__0_ );
   nand U52084 ( n51040,n50666,p1_instqueue_reg_0__0_ );
   nand U52085 ( n51026,n51042,n51043 );
   nor U52086 ( n51043,n51044,n51045 );
   nand U52087 ( n51045,n51046,n51047 );
   nand U52088 ( n51047,n50673,p1_instqueue_reg_15__0_ );
   nand U52089 ( n51046,n50674,p1_instqueue_reg_14__0_ );
   nand U52090 ( n51044,n51048,n51049 );
   nand U52091 ( n51049,n50677,p1_instqueue_reg_13__0_ );
   nand U52092 ( n51048,n50678,p1_instqueue_reg_12__0_ );
   nor U52093 ( n51042,n51050,n51051 );
   nand U52094 ( n51051,n51052,n51053 );
   nand U52095 ( n51053,n50683,p1_instqueue_reg_11__0_ );
   nand U52096 ( n51052,n50684,p1_instqueue_reg_10__0_ );
   nand U52097 ( n51050,n51054,n51055 );
   nand U52098 ( n51055,n50687,p1_instqueue_reg_9__0_ );
   nand U52099 ( n51054,n50688,p1_instqueue_reg_8__0_ );
   nor U52100 ( n51019,n51056,n51057 );
   nor U52101 ( n51057,n50609,n49256 );
   not U52102 ( n49256,p1_eax_reg_16_ );
   nor U52103 ( n51056,n28251,n48572 );
   nand U52104 ( n50320,n51058,n50386 );
   xor U52105 ( n51058,n51059,n28407 );
   xor U52106 ( n50385,n28183,n51060 );
   nand U52107 ( n51060,n51061,n51062 );
   nor U52108 ( n51062,n51063,n51064 );
   nor U52109 ( n51064,n28185,n48672 );
   nand U52110 ( n48672,n51065,n51066 );
   nand U52111 ( n51065,n48675,n51067 );
   nand U52112 ( n51067,n51068,p1_phyaddrpointer_reg_21_ );
   nor U52113 ( n51063,n51069,n50642 );
   nor U52114 ( n51069,n51070,n51071 );
   nand U52115 ( n51071,n51072,n51073 );
   nor U52116 ( n51073,n51074,n51075 );
   nand U52117 ( n51075,n51076,n51077 );
   nand U52118 ( n51077,n50651,p1_instqueue_reg_7__6_ );
   nand U52119 ( n51076,n50652,p1_instqueue_reg_6__6_ );
   nand U52120 ( n51074,n51078,n51079 );
   nand U52121 ( n51079,n50655,p1_instqueue_reg_5__6_ );
   nand U52122 ( n51078,n50656,p1_instqueue_reg_4__6_ );
   nor U52123 ( n51072,n51080,n51081 );
   nand U52124 ( n51081,n51082,n51083 );
   nand U52125 ( n51083,n50661,p1_instqueue_reg_3__6_ );
   nand U52126 ( n51082,n50662,p1_instqueue_reg_2__6_ );
   nand U52127 ( n51080,n51084,n51085 );
   nand U52128 ( n51085,n50665,p1_instqueue_reg_1__6_ );
   nand U52129 ( n51084,n50666,p1_instqueue_reg_0__6_ );
   nand U52130 ( n51070,n51086,n51087 );
   nor U52131 ( n51087,n51088,n51089 );
   nand U52132 ( n51089,n51090,n51091 );
   nand U52133 ( n51091,n50673,p1_instqueue_reg_15__6_ );
   nand U52134 ( n51090,n50674,p1_instqueue_reg_14__6_ );
   nand U52135 ( n51088,n51092,n51093 );
   nand U52136 ( n51093,n50677,p1_instqueue_reg_13__6_ );
   nand U52137 ( n51092,n50678,p1_instqueue_reg_12__6_ );
   nor U52138 ( n51086,n51094,n51095 );
   nand U52139 ( n51095,n51096,n51097 );
   nand U52140 ( n51097,n50683,p1_instqueue_reg_11__6_ );
   nand U52141 ( n51096,n50684,p1_instqueue_reg_10__6_ );
   nand U52142 ( n51094,n51098,n51099 );
   nand U52143 ( n51099,n50687,p1_instqueue_reg_9__6_ );
   nand U52144 ( n51098,n50688,p1_instqueue_reg_8__6_ );
   nor U52145 ( n51061,n51100,n51101 );
   nor U52146 ( n51101,n28287,n49287 );
   not U52147 ( n49287,p1_eax_reg_22_ );
   nor U52148 ( n51100,n28252,n48675 );
   not U52149 ( n48675,p1_phyaddrpointer_reg_22_ );
   and U52150 ( n50388,n51102,n50588 );
   nand U52151 ( n51102,n51103,n51059 );
   and U52152 ( n51059,n51104,n51105 );
   nor U52153 ( n51105,n51106,n51107 );
   nor U52154 ( n51107,n28288,n49272 );
   not U52155 ( n49272,p1_eax_reg_19_ );
   nor U52156 ( n51106,n28182,n48617 );
   nand U52157 ( n48617,n51108,n51109 );
   nand U52158 ( n51109,n50638,n48620 );
   nor U52159 ( n51104,n51110,n51111 );
   nor U52160 ( n51111,n50610,n48620 );
   nor U52161 ( n51110,n51112,n50642 );
   nor U52162 ( n51112,n51113,n51114 );
   nand U52163 ( n51114,n51115,n51116 );
   nor U52164 ( n51116,n51117,n51118 );
   nand U52165 ( n51118,n51119,n51120 );
   nand U52166 ( n51120,n50673,p1_instqueue_reg_15__3_ );
   nand U52167 ( n51119,n50683,p1_instqueue_reg_11__3_ );
   nand U52168 ( n51117,n51121,n51122 );
   nand U52169 ( n51122,n50651,p1_instqueue_reg_7__3_ );
   nand U52170 ( n51121,n50661,p1_instqueue_reg_3__3_ );
   nor U52171 ( n51115,n51123,n51124 );
   nand U52172 ( n51124,n51125,n51126 );
   nand U52173 ( n51126,n50687,p1_instqueue_reg_9__3_ );
   nand U52174 ( n51125,n50688,p1_instqueue_reg_8__3_ );
   nand U52175 ( n51123,n51127,n51128 );
   nand U52176 ( n51128,n50678,p1_instqueue_reg_12__3_ );
   nand U52177 ( n51127,n50684,p1_instqueue_reg_10__3_ );
   nand U52178 ( n51113,n51129,n51130 );
   nor U52179 ( n51130,n51131,n51132 );
   nand U52180 ( n51132,n51133,n51134 );
   nand U52181 ( n51134,n50677,p1_instqueue_reg_13__3_ );
   nand U52182 ( n51133,n50674,p1_instqueue_reg_14__3_ );
   nand U52183 ( n51131,n51135,n51136 );
   nand U52184 ( n51136,n50665,p1_instqueue_reg_1__3_ );
   nand U52185 ( n51135,n50666,p1_instqueue_reg_0__3_ );
   nor U52186 ( n51129,n51137,n51138 );
   nand U52187 ( n51138,n51139,n51140 );
   nand U52188 ( n51140,n50656,p1_instqueue_reg_4__3_ );
   nand U52189 ( n51139,n50662,p1_instqueue_reg_2__3_ );
   nand U52190 ( n51137,n51141,n51142 );
   nand U52191 ( n51142,n50655,p1_instqueue_reg_5__3_ );
   nand U52192 ( n51141,n50652,p1_instqueue_reg_6__3_ );
   and U52193 ( n51103,n50626,n50389 );
   xor U52194 ( n50389,n28183,n51143 );
   nand U52195 ( n51143,n51144,n51145 );
   nor U52196 ( n51145,n51146,n51147 );
   nor U52197 ( n51147,n48652,n28184 );
   xor U52198 ( n48652,n48655,n51068 );
   nor U52199 ( n51146,n51148,n50642 );
   nor U52200 ( n51148,n51149,n51150 );
   nand U52201 ( n51150,n51151,n51152 );
   nor U52202 ( n51152,n51153,n51154 );
   nand U52203 ( n51154,n51155,n51156 );
   nand U52204 ( n51156,n50651,p1_instqueue_reg_7__5_ );
   nand U52205 ( n51155,n50652,p1_instqueue_reg_6__5_ );
   nand U52206 ( n51153,n51157,n51158 );
   nand U52207 ( n51158,n50655,p1_instqueue_reg_5__5_ );
   nand U52208 ( n51157,n50656,p1_instqueue_reg_4__5_ );
   nor U52209 ( n51151,n51159,n51160 );
   nand U52210 ( n51160,n51161,n51162 );
   nand U52211 ( n51162,n50661,p1_instqueue_reg_3__5_ );
   nand U52212 ( n51161,n50662,p1_instqueue_reg_2__5_ );
   nand U52213 ( n51159,n51163,n51164 );
   nand U52214 ( n51164,n50665,p1_instqueue_reg_1__5_ );
   nand U52215 ( n51163,n50666,p1_instqueue_reg_0__5_ );
   nand U52216 ( n51149,n51165,n51166 );
   nor U52217 ( n51166,n51167,n51168 );
   nand U52218 ( n51168,n51169,n51170 );
   nand U52219 ( n51170,n50673,p1_instqueue_reg_15__5_ );
   nand U52220 ( n51169,n50674,p1_instqueue_reg_14__5_ );
   nand U52221 ( n51167,n51171,n51172 );
   nand U52222 ( n51172,n50677,p1_instqueue_reg_13__5_ );
   nand U52223 ( n51171,n50678,p1_instqueue_reg_12__5_ );
   nor U52224 ( n51165,n51173,n51174 );
   nand U52225 ( n51174,n51175,n51176 );
   nand U52226 ( n51176,n50683,p1_instqueue_reg_11__5_ );
   nand U52227 ( n51175,n50684,p1_instqueue_reg_10__5_ );
   nand U52228 ( n51173,n51177,n51178 );
   nand U52229 ( n51178,n50687,p1_instqueue_reg_9__5_ );
   nand U52230 ( n51177,n50688,p1_instqueue_reg_8__5_ );
   nor U52231 ( n51144,n51179,n51180 );
   nor U52232 ( n51180,n50609,n49282 );
   not U52233 ( n49282,p1_eax_reg_21_ );
   nor U52234 ( n51179,n28251,n48655 );
   xor U52235 ( n50626,n28183,n51181 );
   nand U52236 ( n51181,n51182,n51183 );
   nor U52237 ( n51183,n51184,n51185 );
   nor U52238 ( n51185,n28182,n48632 );
   nand U52239 ( n48632,n51186,n51187 );
   nand U52240 ( n51186,n48635,n51108 );
   nor U52241 ( n51184,n51188,n50642 );
   nand U52242 ( n50642,n50737,n51189 );
   nor U52243 ( n51188,n51190,n51191 );
   nand U52244 ( n51191,n51192,n51193 );
   nor U52245 ( n51193,n51194,n51195 );
   nand U52246 ( n51195,n51196,n51197 );
   nand U52247 ( n51197,n50651,p1_instqueue_reg_7__4_ );
   not U52248 ( n50651,n51198 );
   nand U52249 ( n51196,n50652,p1_instqueue_reg_6__4_ );
   not U52250 ( n50652,n51199 );
   nand U52251 ( n51194,n51200,n51201 );
   nand U52252 ( n51201,n50655,p1_instqueue_reg_5__4_ );
   not U52253 ( n50655,n51202 );
   nand U52254 ( n51200,n50656,p1_instqueue_reg_4__4_ );
   not U52255 ( n50656,n51203 );
   nor U52256 ( n51192,n51204,n51205 );
   nand U52257 ( n51205,n51206,n51207 );
   nand U52258 ( n51207,n50661,p1_instqueue_reg_3__4_ );
   not U52259 ( n50661,n51208 );
   nand U52260 ( n51206,n50662,p1_instqueue_reg_2__4_ );
   not U52261 ( n50662,n51209 );
   nand U52262 ( n51204,n51210,n51211 );
   nand U52263 ( n51211,n50665,p1_instqueue_reg_1__4_ );
   not U52264 ( n50665,n51212 );
   nand U52265 ( n51210,n50666,p1_instqueue_reg_0__4_ );
   not U52266 ( n50666,n51213 );
   nand U52267 ( n51190,n51214,n51215 );
   nor U52268 ( n51215,n51216,n51217 );
   nand U52269 ( n51217,n51218,n51219 );
   nand U52270 ( n51219,n50673,p1_instqueue_reg_15__4_ );
   not U52271 ( n50673,n51220 );
   nand U52272 ( n51218,n50674,p1_instqueue_reg_14__4_ );
   not U52273 ( n50674,n51221 );
   nand U52274 ( n51216,n51222,n51223 );
   nand U52275 ( n51223,n50677,p1_instqueue_reg_13__4_ );
   not U52276 ( n50677,n51224 );
   nand U52277 ( n51222,n50678,p1_instqueue_reg_12__4_ );
   not U52278 ( n50678,n51225 );
   nor U52279 ( n51214,n51226,n51227 );
   nand U52280 ( n51227,n51228,n51229 );
   nand U52281 ( n51229,n50683,p1_instqueue_reg_11__4_ );
   not U52282 ( n50683,n51230 );
   nand U52283 ( n51228,n50684,p1_instqueue_reg_10__4_ );
   not U52284 ( n50684,n51231 );
   nand U52285 ( n51226,n51232,n51233 );
   nand U52286 ( n51233,n50687,p1_instqueue_reg_9__4_ );
   not U52287 ( n50687,n51234 );
   nand U52288 ( n51232,n50688,p1_instqueue_reg_8__4_ );
   not U52289 ( n50688,n51235 );
   nor U52290 ( n51182,n51236,n51237 );
   nor U52291 ( n51237,n28287,n49277 );
   not U52292 ( n49277,p1_eax_reg_20_ );
   nor U52293 ( n51236,n28252,n48635 );
   nand U52294 ( n50410,n51238,n50386 );
   xor U52295 ( n51238,n51239,n28408 );
   or U52296 ( n50618,n50453,n51240 );
   and U52297 ( n51240,n50386,n50477 );
   nor U52298 ( n50453,n51241,n50588 );
   nor U52299 ( n50615,n50479,n51242 );
   nor U52300 ( n51242,n50386,n51243 );
   and U52301 ( n51243,n50477,n50617 );
   xor U52302 ( n50617,n51244,n28408 );
   nor U52303 ( n51244,n51245,n51246 );
   nand U52304 ( n51246,n51247,n51248 );
   nand U52305 ( n51248,p1_phyaddrpointer_reg_27_,n49013 );
   nand U52306 ( n51247,p1_eax_reg_27_,n50593 );
   nand U52307 ( n51245,n51249,n51250 );
   nand U52308 ( n51250,n50737,n51251 );
   xor U52309 ( n51251,n51252,n51253 );
   or U52310 ( n51249,n28184,n48762 );
   xor U52311 ( n48762,p1_phyaddrpointer_reg_27_,n51254 );
   xor U52312 ( n50477,n28183,n51255 );
   nand U52313 ( n51255,n51256,n51257 );
   nor U52314 ( n51257,n51258,n51259 );
   nor U52315 ( n51259,n28182,n48739 );
   nand U52316 ( n48739,n51260,n51254 );
   nand U52317 ( n51260,n48742,n51261 );
   nand U52318 ( n51261,n51262,p1_phyaddrpointer_reg_25_ );
   nor U52319 ( n51258,n50604,n51263 );
   nand U52320 ( n51263,n51264,n51253 );
   nand U52321 ( n51264,n51265,n51266 );
   nor U52322 ( n51256,n51267,n51268 );
   nor U52323 ( n51268,n28288,n49307 );
   not U52324 ( n49307,p1_eax_reg_26_ );
   nor U52325 ( n51267,n50610,n48742 );
   not U52326 ( n48742,p1_phyaddrpointer_reg_26_ );
   and U52327 ( n50479,n51269,n50588 );
   nand U52328 ( n51269,n51270,n51239 );
   and U52329 ( n51239,n51271,n51272 );
   nor U52330 ( n51272,n51273,n51274 );
   nor U52331 ( n51274,n28184,n48691 );
   nand U52332 ( n48691,n51275,n51276 );
   nand U52333 ( n51276,n51066,n48694 );
   and U52334 ( n51273,n51277,n28262 );
   xor U52335 ( n51277,n51278,n51279 );
   nor U52336 ( n51271,n51280,n51281 );
   nor U52337 ( n51281,n28251,n48694 );
   nor U52338 ( n51280,n50609,n49292 );
   not U52339 ( n49292,p1_eax_reg_23_ );
   nor U52340 ( n51270,n50620,n51241 );
   xor U52341 ( n51241,n51282,n28182 );
   nor U52342 ( n51282,n51283,n51284 );
   nand U52343 ( n51284,n51285,n51286 );
   nand U52344 ( n51286,p1_phyaddrpointer_reg_25_,n49013 );
   nand U52345 ( n51285,p1_eax_reg_25_,n50593 );
   nand U52346 ( n51283,n51287,n51288 );
   nand U52347 ( n51288,n50737,n51289 );
   xor U52348 ( n51289,n51290,n51291 );
   or U52349 ( n51287,n28185,n48724 );
   xor U52350 ( n48724,n48727,n51262 );
   xor U52351 ( n50620,n49843,n51292 );
   nand U52352 ( n51292,n51293,n51294 );
   nor U52353 ( n51294,n51295,n51296 );
   nor U52354 ( n51296,n28184,n48705 );
   nand U52355 ( n48705,n51297,n51298 );
   nand U52356 ( n51297,n48708,n51275 );
   nor U52357 ( n51295,n50604,n51299 );
   nand U52358 ( n51299,n51300,n51291 );
   nand U52359 ( n51300,n51301,n51302 );
   nor U52360 ( n51293,n51303,n51304 );
   nor U52361 ( n51304,n28287,n49297 );
   not U52362 ( n49297,p1_eax_reg_24_ );
   nor U52363 ( n51303,n28252,n48708 );
   nand U52364 ( n50611,n50614,n50588 );
   not U52365 ( n50588,n50386 );
   nand U52366 ( n50614,n51305,n51306 );
   nor U52367 ( n51306,n51307,n51308 );
   nor U52368 ( n51308,n28185,n48784 );
   nand U52369 ( n48784,n50602,n51309 );
   nand U52370 ( n51309,n51310,n48787 );
   nor U52371 ( n51307,n50604,n51311 );
   nand U52372 ( n51311,n51312,n51313 );
   nand U52373 ( n51312,n51314,n51315 );
   nor U52374 ( n51305,n51316,n51317 );
   nor U52375 ( n51317,n28288,n49317 );
   not U52376 ( n49317,p1_eax_reg_28_ );
   nor U52377 ( n51316,n50610,n48787 );
   not U52378 ( n50594,n50561 );
   nand U52379 ( n50561,n51318,n50386 );
   nand U52380 ( n50386,n50737,n49009 );
   nor U52381 ( n49009,n51319,n48873 );
   and U52382 ( n48873,n48875,n48876 );
   nand U52383 ( n48876,n51320,n51321 );
   nor U52384 ( n51320,n51322,n51323 );
   nor U52385 ( n51323,n28327,n51324 );
   nor U52386 ( n51322,n51325,n51326 );
   not U52387 ( n51325,n51324 );
   nand U52388 ( n51324,n51327,n51328 );
   nor U52389 ( n51328,n51329,n51330 );
   nand U52390 ( n51330,n51331,n51332 );
   nor U52391 ( n51332,n51333,n51334 );
   nor U52392 ( n51334,n51335,n51336 );
   nor U52393 ( n51333,n51337,n51338 );
   nor U52394 ( n51331,n51339,n51340 );
   nor U52395 ( n51340,n51341,n51342 );
   nor U52396 ( n51339,n51343,n51344 );
   nand U52397 ( n51329,n51345,n51346 );
   nor U52398 ( n51346,n51347,n51348 );
   nor U52399 ( n51348,n51349,n51350 );
   nor U52400 ( n51347,n51351,n51352 );
   nor U52401 ( n51345,n51353,n51354 );
   nor U52402 ( n51354,n51355,n51356 );
   nor U52403 ( n51353,n51357,n51358 );
   nor U52404 ( n51327,n51359,n51360 );
   nand U52405 ( n51360,n51361,n51362 );
   nor U52406 ( n51362,n51363,n51364 );
   nor U52407 ( n51364,n51365,n51366 );
   nor U52408 ( n51363,n51367,n51368 );
   nor U52409 ( n51361,n51369,n51370 );
   nor U52410 ( n51370,n51371,n51372 );
   nor U52411 ( n51369,n51373,n51374 );
   nand U52412 ( n51359,n51375,n51376 );
   nor U52413 ( n51376,n51377,n51378 );
   nor U52414 ( n51378,n51379,n51380 );
   nor U52415 ( n51377,n51381,n51382 );
   nor U52416 ( n51375,n51383,n51384 );
   nor U52417 ( n51384,n47243,n51385 );
   nor U52418 ( n51383,n51386,n51387 );
   nor U52419 ( n48875,n50754,n50753 );
   xor U52420 ( n50753,n48996,n51388 );
   nand U52421 ( n51388,n51389,n51390 );
   nand U52422 ( n51390,n51391,n51392 );
   nor U52423 ( n51392,n51393,n51394 );
   nand U52424 ( n51394,n51395,n51396 );
   nor U52425 ( n51396,n51397,n51398 );
   nor U52426 ( n51398,n51399,n51336 );
   nor U52427 ( n51397,n51400,n51338 );
   nor U52428 ( n51395,n51401,n51402 );
   nor U52429 ( n51402,n51403,n51342 );
   nor U52430 ( n51401,n51404,n51344 );
   nand U52431 ( n51393,n51405,n51406 );
   nor U52432 ( n51406,n51407,n51408 );
   nor U52433 ( n51408,n51409,n51350 );
   nor U52434 ( n51407,n51410,n51352 );
   nor U52435 ( n51405,n51411,n51412 );
   nor U52436 ( n51412,n51413,n51356 );
   nor U52437 ( n51411,n51414,n51358 );
   nor U52438 ( n51391,n51415,n51416 );
   nand U52439 ( n51416,n51417,n51418 );
   nor U52440 ( n51418,n51419,n51420 );
   nor U52441 ( n51420,n51421,n51366 );
   nor U52442 ( n51419,n51422,n51368 );
   nor U52443 ( n51417,n51423,n51424 );
   nor U52444 ( n51424,n51425,n51372 );
   nor U52445 ( n51423,n51426,n51374 );
   nand U52446 ( n51415,n51427,n51428 );
   nor U52447 ( n51428,n51429,n51430 );
   nor U52448 ( n51430,n51431,n51380 );
   nor U52449 ( n51429,n51432,n51382 );
   nor U52450 ( n51427,n51433,n51434 );
   nor U52451 ( n51434,n47260,n51385 );
   nor U52452 ( n51433,n51435,n51387 );
   or U52453 ( n50754,n50768,n50767 );
   and U52454 ( n50767,n51436,n51321 );
   nor U52455 ( n51436,n51437,n51438 );
   nor U52456 ( n51438,n28327,n51439 );
   nor U52457 ( n51437,n51440,n51326 );
   not U52458 ( n51440,n51439 );
   nand U52459 ( n51439,n51441,n51442 );
   nor U52460 ( n51442,n51443,n51444 );
   nand U52461 ( n51444,n51445,n51446 );
   nor U52462 ( n51446,n51447,n51448 );
   nor U52463 ( n51448,n51449,n51336 );
   nor U52464 ( n51447,n51450,n51338 );
   nor U52465 ( n51445,n51451,n51452 );
   nor U52466 ( n51452,n51453,n51342 );
   nor U52467 ( n51451,n51454,n51344 );
   nand U52468 ( n51443,n51455,n51456 );
   nor U52469 ( n51456,n51457,n51458 );
   nor U52470 ( n51458,n51459,n51350 );
   nor U52471 ( n51457,n51460,n51352 );
   nor U52472 ( n51455,n51461,n51462 );
   nor U52473 ( n51462,n51463,n51356 );
   nor U52474 ( n51461,n51464,n51358 );
   nor U52475 ( n51441,n51465,n51466 );
   nand U52476 ( n51466,n51467,n51468 );
   nor U52477 ( n51468,n51469,n51470 );
   nor U52478 ( n51470,n51471,n51366 );
   nor U52479 ( n51469,n51472,n51368 );
   nor U52480 ( n51467,n51473,n51474 );
   nor U52481 ( n51474,n51475,n51372 );
   nor U52482 ( n51473,n51476,n51374 );
   nand U52483 ( n51465,n51477,n51478 );
   nor U52484 ( n51478,n51479,n51480 );
   nor U52485 ( n51480,n51481,n51380 );
   nor U52486 ( n51479,n51482,n51382 );
   nor U52487 ( n51477,n51483,n51484 );
   nor U52488 ( n51484,n47276,n51385 );
   nor U52489 ( n51483,n51485,n51387 );
   nand U52490 ( n50768,n51486,n50783 );
   nor U52491 ( n50783,n51004,n51003 );
   and U52492 ( n51003,n51487,n51321 );
   nor U52493 ( n51487,n51488,n51489 );
   nor U52494 ( n51489,n51319,n51490 );
   nor U52495 ( n51488,n51491,n51326 );
   not U52496 ( n51491,n51490 );
   nand U52497 ( n51490,n51492,n51493 );
   nor U52498 ( n51493,n51494,n51495 );
   nand U52499 ( n51495,n51496,n51497 );
   nor U52500 ( n51497,n51498,n51499 );
   nor U52501 ( n51499,n51500,n51336 );
   nor U52502 ( n51498,n51501,n51338 );
   nor U52503 ( n51496,n51502,n51503 );
   nor U52504 ( n51503,n51504,n51342 );
   nor U52505 ( n51502,n51505,n51344 );
   nand U52506 ( n51494,n51506,n51507 );
   nor U52507 ( n51507,n51508,n51509 );
   nor U52508 ( n51509,n51510,n51350 );
   nor U52509 ( n51508,n51511,n51352 );
   nor U52510 ( n51506,n51512,n51513 );
   nor U52511 ( n51513,n51514,n51356 );
   nor U52512 ( n51512,n51515,n51358 );
   nor U52513 ( n51492,n51516,n51517 );
   nand U52514 ( n51517,n51518,n51519 );
   nor U52515 ( n51519,n51520,n51521 );
   nor U52516 ( n51521,n51522,n51366 );
   nor U52517 ( n51520,n51523,n51368 );
   nor U52518 ( n51518,n51524,n51525 );
   nor U52519 ( n51525,n51526,n51372 );
   nor U52520 ( n51524,n51527,n51374 );
   nand U52521 ( n51516,n51528,n51529 );
   nor U52522 ( n51529,n51530,n51531 );
   nor U52523 ( n51531,n51532,n51380 );
   nor U52524 ( n51530,n51533,n51382 );
   nor U52525 ( n51528,n51534,n51535 );
   nor U52526 ( n51535,n47323,n51385 );
   nor U52527 ( n51534,n51536,n51387 );
   nand U52528 ( n51004,n50811,n50810 );
   nand U52529 ( n50810,n51537,n51321 );
   nor U52530 ( n51537,n51538,n51539 );
   nor U52531 ( n51539,n51319,n51540 );
   nor U52532 ( n51538,n51541,n51326 );
   not U52533 ( n51541,n51540 );
   nand U52534 ( n51540,n51542,n51543 );
   nor U52535 ( n51543,n51544,n51545 );
   nand U52536 ( n51545,n51546,n51547 );
   nor U52537 ( n51547,n51548,n51549 );
   nor U52538 ( n51549,n51550,n51336 );
   nor U52539 ( n51548,n51551,n51338 );
   nor U52540 ( n51546,n51552,n51553 );
   nor U52541 ( n51553,n51554,n51342 );
   nor U52542 ( n51552,n51555,n51344 );
   nand U52543 ( n51544,n51556,n51557 );
   nor U52544 ( n51557,n51558,n51559 );
   nor U52545 ( n51559,n51560,n51350 );
   nor U52546 ( n51558,n51561,n51352 );
   nor U52547 ( n51556,n51562,n51563 );
   nor U52548 ( n51563,n51564,n51356 );
   nor U52549 ( n51562,n51565,n51358 );
   nor U52550 ( n51542,n51566,n51567 );
   nand U52551 ( n51567,n51568,n51569 );
   nor U52552 ( n51569,n51570,n51571 );
   nor U52553 ( n51571,n51572,n51366 );
   nor U52554 ( n51570,n51573,n51368 );
   nor U52555 ( n51568,n51574,n51575 );
   nor U52556 ( n51575,n51576,n51372 );
   nor U52557 ( n51574,n51577,n51374 );
   nand U52558 ( n51566,n51578,n51579 );
   nor U52559 ( n51579,n51580,n51581 );
   nor U52560 ( n51581,n51582,n51380 );
   nor U52561 ( n51580,n51583,n51382 );
   nor U52562 ( n51578,n51584,n51585 );
   nor U52563 ( n51585,n47339,n51385 );
   nor U52564 ( n51584,n51586,n51387 );
   and U52565 ( n50811,n48969,n48970 );
   nand U52566 ( n48970,n51587,n51321 );
   nor U52567 ( n51587,n51588,n51589 );
   nor U52568 ( n51589,n51319,n51590 );
   nor U52569 ( n51588,n51591,n51326 );
   not U52570 ( n51591,n51590 );
   nand U52571 ( n51590,n51592,n51593 );
   nor U52572 ( n51593,n51594,n51595 );
   nand U52573 ( n51595,n51596,n51597 );
   nor U52574 ( n51597,n51598,n51599 );
   nor U52575 ( n51599,n51600,n51336 );
   nor U52576 ( n51598,n51601,n51338 );
   nor U52577 ( n51596,n51602,n51603 );
   nor U52578 ( n51603,n51604,n51342 );
   nor U52579 ( n51602,n51605,n51344 );
   nand U52580 ( n51594,n51606,n51607 );
   nor U52581 ( n51607,n51608,n51609 );
   nor U52582 ( n51609,n51610,n51350 );
   nor U52583 ( n51608,n51611,n51352 );
   nor U52584 ( n51606,n51612,n51613 );
   nor U52585 ( n51613,n51614,n51356 );
   nor U52586 ( n51612,n51615,n51358 );
   nor U52587 ( n51592,n51616,n51617 );
   nand U52588 ( n51617,n51618,n51619 );
   nor U52589 ( n51619,n51620,n51621 );
   nor U52590 ( n51621,n51622,n51366 );
   nor U52591 ( n51620,n51623,n51368 );
   nor U52592 ( n51618,n51624,n51625 );
   nor U52593 ( n51625,n51626,n51372 );
   nor U52594 ( n51624,n51627,n51374 );
   nand U52595 ( n51616,n51628,n51629 );
   nor U52596 ( n51629,n51630,n51631 );
   nor U52597 ( n51631,n51632,n51380 );
   nor U52598 ( n51630,n51633,n51382 );
   nor U52599 ( n51628,n51634,n51635 );
   nor U52600 ( n51635,n47364,n51385 );
   nor U52601 ( n51634,n51636,n51387 );
   nand U52602 ( n48969,n50994,n51637 );
   nand U52603 ( n51637,n51638,n50993 );
   or U52604 ( n50993,n51639,n48996 );
   nand U52605 ( n51638,n50969,n51640 );
   nand U52606 ( n51640,n50967,n50968 );
   not U52607 ( n50968,n50992 );
   nor U52608 ( n50992,n51641,n51642 );
   nand U52609 ( n50967,n50962,n51643 );
   nand U52610 ( n51643,n50960,n50961 );
   nand U52611 ( n50961,n51644,n51645 );
   nand U52612 ( n50960,n50943,n51646 );
   nand U52613 ( n51646,n50944,n50942 );
   or U52614 ( n50942,n51647,n51648 );
   nand U52615 ( n50944,n50916,n51649 );
   nand U52616 ( n51649,n51650,n50917 );
   nand U52617 ( n50917,n51651,n51652 );
   nor U52618 ( n51650,n50920,n50901 );
   nor U52619 ( n50901,n50897,n50919 );
   not U52620 ( n50919,n50900 );
   nand U52621 ( n50900,n51653,n51654 );
   or U52622 ( n51654,n51655,n48996 );
   nor U52623 ( n51653,n51656,n48980 );
   not U52624 ( n50897,n50921 );
   nand U52625 ( n50921,n50881,n51657 );
   nand U52626 ( n51657,n50851,n50880 );
   or U52627 ( n50880,n51658,n51659 );
   nor U52628 ( n50851,n50850,n48996 );
   and U52629 ( n50850,n51660,n51661 );
   or U52630 ( n51661,n50857,n28095 );
   nand U52631 ( n50857,n51662,n51663 );
   nand U52632 ( n51663,n51664,n48950 );
   nand U52633 ( n51662,n48247,n48978 );
   xor U52634 ( n51660,n50856,n48996 );
   nand U52635 ( n50856,n51665,n51666 );
   nand U52636 ( n51666,n45834,n28095 );
   not U52637 ( n45834,n45394 );
   nand U52638 ( n45394,n51667,n51668 );
   nand U52639 ( n51668,n51669,n51670 );
   nor U52640 ( n51665,n51671,n51672 );
   nor U52641 ( n51672,n48950,n28327 );
   nor U52642 ( n51671,n48933,n51673 );
   not U52643 ( n48933,n48950 );
   nand U52644 ( n48950,n51674,n51675 );
   nor U52645 ( n51675,n51676,n51677 );
   nand U52646 ( n51677,n51678,n51679 );
   nor U52647 ( n51679,n51680,n51681 );
   nor U52648 ( n51681,n51636,n51682 );
   nor U52649 ( n51680,n51632,n51683 );
   nor U52650 ( n51678,n51684,n51685 );
   nor U52651 ( n51685,n51633,n51686 );
   nor U52652 ( n51684,n51627,n51687 );
   nand U52653 ( n51676,n51688,n51689 );
   nor U52654 ( n51689,n51690,n51691 );
   nor U52655 ( n51691,n51622,n51692 );
   nor U52656 ( n51690,n51623,n51693 );
   nor U52657 ( n51688,n51694,n51695 );
   nor U52658 ( n51695,n51615,n51696 );
   nor U52659 ( n51694,n51610,n51697 );
   nor U52660 ( n51674,n51698,n51699 );
   nand U52661 ( n51699,n51700,n51701 );
   nor U52662 ( n51701,n51702,n51703 );
   nor U52663 ( n51703,n51611,n51704 );
   nor U52664 ( n51702,n51605,n51705 );
   nor U52665 ( n51700,n51706,n51707 );
   nor U52666 ( n51707,n51600,n51708 );
   nor U52667 ( n51706,n51601,n51709 );
   nand U52668 ( n51698,n51710,n51711 );
   nor U52669 ( n51711,n51712,n51713 );
   nor U52670 ( n51713,n47364,n51714 );
   nor U52671 ( n51712,n51626,n51715 );
   nor U52672 ( n51710,n51716,n51717 );
   nor U52673 ( n51717,n51614,n51718 );
   nor U52674 ( n51716,n51604,n51719 );
   nand U52675 ( n50881,n51659,n51658 );
   xor U52676 ( n51658,n51319,n51720 );
   nand U52677 ( n51720,n51721,n51722 );
   nand U52678 ( n51722,n46090,n45347 );
   not U52679 ( n46090,n45404 );
   xor U52680 ( n45404,n51723,n51724 );
   xor U52681 ( n51723,n51725,n51667 );
   nor U52682 ( n51721,n51726,n51727 );
   nor U52683 ( n51727,n28327,n48982 );
   nor U52684 ( n51726,n48934,n51673 );
   and U52685 ( n51659,n51728,n51729 );
   nand U52686 ( n51729,n51730,p1_instqueue_reg_0__1_ );
   nor U52687 ( n51728,n51731,n51732 );
   nor U52688 ( n51732,n48934,n51733 );
   not U52689 ( n48934,n48982 );
   nand U52690 ( n48982,n51734,n51735 );
   nor U52691 ( n51735,n51736,n51737 );
   nand U52692 ( n51737,n51738,n51739 );
   nor U52693 ( n51739,n51740,n51741 );
   nor U52694 ( n51741,n51586,n51682 );
   nor U52695 ( n51740,n51582,n51683 );
   nor U52696 ( n51738,n51742,n51743 );
   nor U52697 ( n51743,n51583,n51686 );
   nor U52698 ( n51742,n51577,n51687 );
   nand U52699 ( n51736,n51744,n51745 );
   nor U52700 ( n51745,n51746,n51747 );
   nor U52701 ( n51747,n51572,n51692 );
   nor U52702 ( n51746,n51573,n51693 );
   nor U52703 ( n51744,n51748,n51749 );
   nor U52704 ( n51749,n51565,n51696 );
   nor U52705 ( n51748,n51560,n51697 );
   nor U52706 ( n51734,n51750,n51751 );
   nand U52707 ( n51751,n51752,n51753 );
   nor U52708 ( n51753,n51754,n51755 );
   nor U52709 ( n51755,n51561,n51704 );
   nor U52710 ( n51754,n51555,n51705 );
   nor U52711 ( n51752,n51756,n51757 );
   nor U52712 ( n51757,n51550,n51708 );
   nor U52713 ( n51756,n51551,n51709 );
   nand U52714 ( n51750,n51758,n51759 );
   nor U52715 ( n51759,n51760,n51761 );
   nor U52716 ( n51761,n47339,n51714 );
   nor U52717 ( n51760,n51576,n51715 );
   nor U52718 ( n51758,n51762,n51763 );
   nor U52719 ( n51763,n51564,n51718 );
   nor U52720 ( n51762,n51554,n51719 );
   not U52721 ( n50920,n50899 );
   nand U52722 ( n50899,n51764,n51765 );
   xor U52723 ( n51765,n51655,n51319 );
   nand U52724 ( n51655,n51766,n51767 );
   nand U52725 ( n51767,n46612,n28094 );
   not U52726 ( n46612,n45417 );
   xor U52727 ( n45417,n51768,n51769 );
   nor U52728 ( n51768,n51770,n51771 );
   nor U52729 ( n51766,n51772,n51773 );
   nor U52730 ( n51773,n51319,n48932 );
   nor U52731 ( n51772,n48980,n51673 );
   nor U52732 ( n51764,n51774,n51775 );
   nor U52733 ( n51775,n48270,n47323 );
   nor U52734 ( n51774,n48980,n51733 );
   not U52735 ( n48980,n48932 );
   nand U52736 ( n48932,n51776,n51777 );
   nor U52737 ( n51777,n51778,n51779 );
   nand U52738 ( n51779,n51780,n51781 );
   nor U52739 ( n51781,n51782,n51783 );
   nor U52740 ( n51783,n51536,n51682 );
   nor U52741 ( n51782,n51532,n51683 );
   nor U52742 ( n51780,n51784,n51785 );
   nor U52743 ( n51785,n51533,n51686 );
   nor U52744 ( n51784,n51527,n51687 );
   nand U52745 ( n51778,n51786,n51787 );
   nor U52746 ( n51787,n51788,n51789 );
   nor U52747 ( n51789,n51522,n51692 );
   nor U52748 ( n51788,n51523,n51693 );
   nor U52749 ( n51786,n51790,n51791 );
   nor U52750 ( n51791,n51515,n51696 );
   nor U52751 ( n51790,n51510,n51697 );
   nor U52752 ( n51776,n51792,n51793 );
   nand U52753 ( n51793,n51794,n51795 );
   nor U52754 ( n51795,n51796,n51797 );
   nor U52755 ( n51797,n51511,n51704 );
   nor U52756 ( n51796,n51505,n51705 );
   nor U52757 ( n51794,n51798,n51799 );
   nor U52758 ( n51799,n51500,n51708 );
   nor U52759 ( n51798,n51501,n51709 );
   nand U52760 ( n51792,n51800,n51801 );
   nor U52761 ( n51801,n51802,n51803 );
   nor U52762 ( n51803,n47323,n51714 );
   nor U52763 ( n51802,n51526,n51715 );
   nor U52764 ( n51800,n51804,n51805 );
   nor U52765 ( n51805,n51514,n51718 );
   nor U52766 ( n51804,n51504,n51719 );
   or U52767 ( n50916,n51652,n51651 );
   and U52768 ( n51651,n51806,n51807 );
   nand U52769 ( n51807,n51664,n48915 );
   nand U52770 ( n51806,p1_instqueue_reg_0__3_,n51730 );
   xor U52771 ( n51652,n51319,n51808 );
   nand U52772 ( n51808,n51809,n51810 );
   nand U52773 ( n51810,n46954,n28095 );
   xor U52774 ( n46954,n50937,n50936 );
   nor U52775 ( n50936,n51811,n51769 );
   nand U52776 ( n51769,n51812,n51813 );
   nand U52777 ( n51813,n51814,n51667 );
   or U52778 ( n51667,n51670,n51669 );
   and U52779 ( n51669,n51815,n51816 );
   nor U52780 ( n51816,n51817,n51818 );
   nand U52781 ( n51818,n51819,n48206 );
   nand U52782 ( n48206,n51820,n45876 );
   nor U52783 ( n51820,n51821,n51822 );
   nor U52784 ( n51822,n47287,n48863 );
   not U52785 ( n48863,n48870 );
   nor U52786 ( n51821,n51823,n51824 );
   nand U52787 ( n51824,n51825,n48289 );
   nor U52788 ( n51825,n51826,n51827 );
   nor U52789 ( n51827,n47446,n51828 );
   nor U52790 ( n51828,n47287,n51829 );
   nand U52791 ( n51829,n47255,n49632 );
   nor U52792 ( n51826,n45878,n51830 );
   nand U52793 ( n51830,n51831,n49632 );
   not U52794 ( n49632,n49827 );
   nand U52795 ( n51831,n48218,n47287 );
   nand U52796 ( n51823,n47236,n51832 );
   nand U52797 ( n51819,n51833,n47334 );
   nand U52798 ( n51833,n51834,n51835 );
   nor U52799 ( n51835,n45876,n48209 );
   nor U52800 ( n48209,n49431,n48247 );
   nor U52801 ( n51834,n45877,n48266 );
   nor U52802 ( n51817,n51836,n51837 );
   nor U52803 ( n51837,n45358,n48200 );
   nor U52804 ( n48200,n47255,n48216 );
   nor U52805 ( n51836,n51838,n51839 );
   nand U52806 ( n51839,n48259,n48247 );
   nand U52807 ( n51838,n47303,n48260 );
   nor U52808 ( n51815,n51840,n45772 );
   nand U52809 ( n45772,n45443,p1_state2_reg_0_ );
   nor U52810 ( n51840,n45876,n47446 );
   nand U52811 ( n51670,n51841,n51842 );
   nand U52812 ( n51842,n51843,n51844 );
   nand U52813 ( n51844,p1_instqueuerd_addr_reg_0_,n51845 );
   nor U52814 ( n51843,p1_instqueuewr_addr_reg_0_,n45342 );
   nand U52815 ( n51841,n45759,n51846 );
   nand U52816 ( n51846,n51847,n51848 );
   nand U52817 ( n51848,n51849,p1_instqueuewr_addr_reg_0_ );
   nand U52818 ( n51847,n49019,n45451 );
   nand U52819 ( n51814,n51725,n51724 );
   or U52820 ( n51812,n51725,n51724 );
   nand U52821 ( n51724,n51850,n51851 );
   nand U52822 ( n51851,p1_instqueuerd_addr_reg_1_,n51845 );
   nor U52823 ( n51850,n51852,n51853 );
   nor U52824 ( n51853,n45759,n45842 );
   nor U52825 ( n51852,n46447,n49019 );
   nor U52826 ( n46447,n46185,n46098 );
   nor U52827 ( n46098,n45842,p1_instqueuewr_addr_reg_0_ );
   nor U52828 ( n46185,n51854,p1_instqueuewr_addr_reg_1_ );
   nand U52829 ( n51725,n51855,n51856 );
   nand U52830 ( n51856,n51857,n51858 );
   nor U52831 ( n51858,n47271,n51859 );
   nand U52832 ( n51859,n48289,p1_state2_reg_0_ );
   nor U52833 ( n51857,n48286,n48216 );
   nand U52834 ( n48216,n49829,n45876 );
   nor U52835 ( n49829,n47303,n45878 );
   nor U52836 ( n51855,n51860,n51861 );
   not U52837 ( n51861,n51862 );
   or U52838 ( n51811,n51771,n51770 );
   and U52839 ( n51770,n51863,n47402 );
   and U52840 ( n51771,n51863,n51849 );
   and U52841 ( n51863,n51864,n51865 );
   nand U52842 ( n51865,n45342,n46445 );
   xor U52843 ( n46445,p1_instqueuewr_addr_reg_2_,n46008 );
   nand U52844 ( n51864,p1_instqueuewr_addr_reg_2_,n49624 );
   nand U52845 ( n50937,n51866,n51867 );
   nand U52846 ( n51867,p1_instqueuewr_addr_reg_3_,n49624 );
   nor U52847 ( n51866,n51868,n51869 );
   nor U52848 ( n51869,n51849,n50913 );
   not U52849 ( n51849,n51845 );
   nand U52850 ( n51845,n51870,n51871 );
   nor U52851 ( n51871,n51872,n51873 );
   nand U52852 ( n51873,n51862,n51874 );
   nand U52853 ( n51874,n51730,n48260 );
   not U52854 ( n48260,n49431 );
   nand U52855 ( n51862,n51875,n51876 );
   nor U52856 ( n51875,n51877,n45347 );
   nor U52857 ( n51877,n51878,n51879 );
   nor U52858 ( n51879,n51880,n48912 );
   nand U52859 ( n51872,n51881,n51882 );
   not U52860 ( n51882,n45350 );
   nand U52861 ( n51881,n51883,n45329 );
   nor U52862 ( n51883,n48219,n28095 );
   not U52863 ( n48219,n48266 );
   nand U52864 ( n48266,n48259,n51884 );
   nand U52865 ( n51884,n49431,n48247 );
   nor U52866 ( n51870,n51885,n51886 );
   nand U52867 ( n51886,n51887,n51888 );
   nand U52868 ( n51888,n48210,p1_state2_reg_0_ );
   nand U52869 ( n51887,n49622,n51889 );
   nand U52870 ( n51889,n47303,n51832 );
   nand U52871 ( n51832,n47303,n47420 );
   nor U52872 ( n51885,n51890,n28095 );
   nor U52873 ( n51890,n48220,n51891 );
   nand U52874 ( n51891,n47446,n51892 );
   nand U52875 ( n51892,n45358,n51893 );
   nand U52876 ( n51893,n48259,n51894 );
   nand U52877 ( n51894,n48218,n51895 );
   nor U52878 ( n48259,n47426,n49827 );
   nor U52879 ( n49827,n47271,n48218 );
   nor U52880 ( n48220,n28404,n45879 );
   nor U52881 ( n51868,n46446,n49019 );
   not U52882 ( n46446,n47127 );
   nand U52883 ( n47127,n51896,n51897 );
   nand U52884 ( n51897,p1_instqueuewr_addr_reg_3_,n45820 );
   not U52885 ( n45820,n46008 );
   nor U52886 ( n51896,n46363,n46702 );
   not U52887 ( n46702,n46629 );
   nand U52888 ( n46629,n46790,n46008 );
   nor U52889 ( n46008,n51854,n45842 );
   not U52890 ( n51854,p1_instqueuewr_addr_reg_0_ );
   nor U52891 ( n46790,n45840,p1_instqueuewr_addr_reg_3_ );
   nor U52892 ( n46363,n46275,p1_instqueuewr_addr_reg_2_ );
   nor U52893 ( n51809,n51898,n51899 );
   nor U52894 ( n51899,n51319,n48915 );
   and U52895 ( n51898,n48915,n51731 );
   nand U52896 ( n48915,n51900,n51901 );
   nor U52897 ( n51901,n51902,n51903 );
   nand U52898 ( n51903,n51904,n51905 );
   nor U52899 ( n51905,n51906,n51907 );
   nor U52900 ( n51907,n51908,n51682 );
   nor U52901 ( n51906,n51909,n51683 );
   nor U52902 ( n51904,n51910,n51911 );
   nor U52903 ( n51911,n51912,n51686 );
   nor U52904 ( n51910,n51913,n51687 );
   nand U52905 ( n51902,n51914,n51915 );
   nor U52906 ( n51915,n51916,n51917 );
   nor U52907 ( n51917,n51918,n51692 );
   nor U52908 ( n51916,n51919,n51693 );
   nor U52909 ( n51914,n51920,n51921 );
   nor U52910 ( n51921,n51922,n51696 );
   nor U52911 ( n51920,n51923,n51697 );
   nor U52912 ( n51900,n51924,n51925 );
   nand U52913 ( n51925,n51926,n51927 );
   nor U52914 ( n51927,n51928,n51929 );
   nor U52915 ( n51929,n51930,n51704 );
   nor U52916 ( n51928,n51931,n51705 );
   nor U52917 ( n51926,n51932,n51933 );
   nor U52918 ( n51933,n51934,n51708 );
   nor U52919 ( n51932,n51935,n51709 );
   nand U52920 ( n51924,n51936,n51937 );
   nor U52921 ( n51937,n51938,n51939 );
   nor U52922 ( n51939,n47308,n51714 );
   nor U52923 ( n51938,n51940,n51715 );
   nor U52924 ( n51936,n51941,n51942 );
   nor U52925 ( n51942,n51943,n51718 );
   nor U52926 ( n51941,n51944,n51719 );
   nand U52927 ( n50943,n51648,n51647 );
   nand U52928 ( n51647,n51945,n51946 );
   nand U52929 ( n51946,n51664,n48913 );
   nand U52930 ( n51945,n51730,p1_instqueue_reg_0__4_ );
   and U52931 ( n51648,n51947,n48913 );
   nand U52932 ( n48913,n51948,n51949 );
   nor U52933 ( n51949,n51950,n51951 );
   nand U52934 ( n51951,n51952,n51953 );
   nor U52935 ( n51953,n51954,n51955 );
   nor U52936 ( n51955,n51956,n51682 );
   nor U52937 ( n51954,n51957,n51683 );
   nor U52938 ( n51952,n51958,n51959 );
   nor U52939 ( n51959,n51960,n51686 );
   nor U52940 ( n51958,n51961,n51687 );
   nand U52941 ( n51950,n51962,n51963 );
   nor U52942 ( n51963,n51964,n51965 );
   nor U52943 ( n51965,n51966,n51692 );
   nor U52944 ( n51964,n51967,n51693 );
   nor U52945 ( n51962,n51968,n51969 );
   nor U52946 ( n51969,n51970,n51696 );
   nor U52947 ( n51968,n51971,n51697 );
   nor U52948 ( n51948,n51972,n51973 );
   nand U52949 ( n51973,n51974,n51975 );
   nor U52950 ( n51975,n51976,n51977 );
   nor U52951 ( n51977,n51978,n51704 );
   nor U52952 ( n51976,n51979,n51705 );
   nor U52953 ( n51974,n51980,n51981 );
   nor U52954 ( n51981,n51982,n51708 );
   nor U52955 ( n51980,n51983,n51709 );
   nand U52956 ( n51972,n51984,n51985 );
   nor U52957 ( n51985,n51986,n51987 );
   nor U52958 ( n51987,n47292,n51714 );
   nor U52959 ( n51986,n51988,n51715 );
   nor U52960 ( n51984,n51989,n51990 );
   nor U52961 ( n51990,n51991,n51718 );
   nor U52962 ( n51989,n51992,n51719 );
   not U52963 ( n50962,n50987 );
   nor U52964 ( n50987,n51645,n51644 );
   and U52965 ( n51644,n51993,n51994 );
   nand U52966 ( n51994,n51664,n48904 );
   nand U52967 ( n51993,n51730,p1_instqueue_reg_0__5_ );
   nand U52968 ( n51645,n51947,n48904 );
   nand U52969 ( n48904,n51995,n51996 );
   nor U52970 ( n51996,n51997,n51998 );
   nand U52971 ( n51998,n51999,n52000 );
   nor U52972 ( n52000,n52001,n52002 );
   nor U52973 ( n52002,n51485,n51682 );
   nor U52974 ( n52001,n51481,n51683 );
   nor U52975 ( n51999,n52003,n52004 );
   nor U52976 ( n52004,n51482,n51686 );
   nor U52977 ( n52003,n51476,n51687 );
   nand U52978 ( n51997,n52005,n52006 );
   nor U52979 ( n52006,n52007,n52008 );
   nor U52980 ( n52008,n51471,n51692 );
   nor U52981 ( n52007,n51472,n51693 );
   nor U52982 ( n52005,n52009,n52010 );
   nor U52983 ( n52010,n51464,n51696 );
   nor U52984 ( n52009,n51459,n51697 );
   nor U52985 ( n51995,n52011,n52012 );
   nand U52986 ( n52012,n52013,n52014 );
   nor U52987 ( n52014,n52015,n52016 );
   nor U52988 ( n52016,n51460,n51704 );
   nor U52989 ( n52015,n51454,n51705 );
   nor U52990 ( n52013,n52017,n52018 );
   nor U52991 ( n52018,n51449,n51708 );
   nor U52992 ( n52017,n51450,n51709 );
   nand U52993 ( n52011,n52019,n52020 );
   nor U52994 ( n52020,n52021,n52022 );
   nor U52995 ( n52022,n47276,n51714 );
   nor U52996 ( n52021,n51475,n51715 );
   nor U52997 ( n52019,n52023,n52024 );
   nor U52998 ( n52024,n51463,n51718 );
   nor U52999 ( n52023,n51453,n51719 );
   nand U53000 ( n50969,n51642,n51641 );
   nand U53001 ( n51641,n52025,n52026 );
   nand U53002 ( n52026,n51664,n48954 );
   nand U53003 ( n52025,p1_instqueue_reg_0__6_,n51730 );
   and U53004 ( n51642,n51947,n48954 );
   nand U53005 ( n48954,n52027,n52028 );
   nor U53006 ( n52028,n52029,n52030 );
   nand U53007 ( n52030,n52031,n52032 );
   nor U53008 ( n52032,n52033,n52034 );
   nor U53009 ( n52034,n51435,n51682 );
   nor U53010 ( n52033,n51431,n51683 );
   nor U53011 ( n52031,n52035,n52036 );
   nor U53012 ( n52036,n51432,n51686 );
   nor U53013 ( n52035,n51426,n51687 );
   nand U53014 ( n52029,n52037,n52038 );
   nor U53015 ( n52038,n52039,n52040 );
   nor U53016 ( n52040,n51421,n51692 );
   nor U53017 ( n52039,n51422,n51693 );
   nor U53018 ( n52037,n52041,n52042 );
   nor U53019 ( n52042,n51414,n51696 );
   nor U53020 ( n52041,n51409,n51697 );
   nor U53021 ( n52027,n52043,n52044 );
   nand U53022 ( n52044,n52045,n52046 );
   nor U53023 ( n52046,n52047,n52048 );
   nor U53024 ( n52048,n51410,n51704 );
   nor U53025 ( n52047,n51404,n51705 );
   nor U53026 ( n52045,n52049,n52050 );
   nor U53027 ( n52050,n51399,n51708 );
   nor U53028 ( n52049,n51400,n51709 );
   nand U53029 ( n52043,n52051,n52052 );
   nor U53030 ( n52052,n52053,n52054 );
   nor U53031 ( n52054,n47260,n51714 );
   nor U53032 ( n52053,n51425,n51715 );
   nor U53033 ( n52051,n52055,n52056 );
   nor U53034 ( n52056,n51413,n51718 );
   nor U53035 ( n52055,n51403,n51719 );
   nand U53036 ( n51947,n28327,n51673 );
   not U53037 ( n51673,n51731 );
   nor U53038 ( n51731,n48978,n52057 );
   nand U53039 ( n50994,n48996,n51639 );
   nand U53040 ( n51639,n52058,n52059 );
   nand U53041 ( n52059,n51664,n48978 );
   nand U53042 ( n52058,p1_instqueue_reg_0__7_,n51730 );
   nor U53043 ( n51486,n51016,n50781 );
   xor U53044 ( n50781,n48996,n52060 );
   nand U53045 ( n52060,n51389,n52061 );
   nand U53046 ( n52061,n52062,n52063 );
   nor U53047 ( n52063,n52064,n52065 );
   nand U53048 ( n52065,n52066,n52067 );
   nor U53049 ( n52067,n52068,n52069 );
   nor U53050 ( n52069,n51982,n51336 );
   nor U53051 ( n52068,n51983,n51338 );
   nor U53052 ( n52066,n52070,n52071 );
   nor U53053 ( n52071,n51992,n51342 );
   nor U53054 ( n52070,n51979,n51344 );
   nand U53055 ( n52064,n52072,n52073 );
   nor U53056 ( n52073,n52074,n52075 );
   nor U53057 ( n52075,n51971,n51350 );
   nor U53058 ( n52074,n51978,n51352 );
   nor U53059 ( n52072,n52076,n52077 );
   nor U53060 ( n52077,n51991,n51356 );
   nor U53061 ( n52076,n51970,n51358 );
   nor U53062 ( n52062,n52078,n52079 );
   nand U53063 ( n52079,n52080,n52081 );
   nor U53064 ( n52081,n52082,n52083 );
   nor U53065 ( n52083,n51966,n51366 );
   nor U53066 ( n52082,n51967,n51368 );
   nor U53067 ( n52080,n52084,n52085 );
   nor U53068 ( n52085,n51988,n51372 );
   nor U53069 ( n52084,n51961,n51374 );
   nand U53070 ( n52078,n52086,n52087 );
   nor U53071 ( n52087,n52088,n52089 );
   nor U53072 ( n52089,n51957,n51380 );
   nor U53073 ( n52088,n51960,n51382 );
   nor U53074 ( n52086,n52090,n52091 );
   nor U53075 ( n52091,n47292,n51385 );
   nor U53076 ( n52090,n51956,n51387 );
   not U53077 ( n51016,n50784 );
   nand U53078 ( n50784,n52092,n51321 );
   nand U53079 ( n51321,n51656,n48996 );
   nor U53080 ( n52092,n52093,n52094 );
   nor U53081 ( n52094,n28327,n52095 );
   nor U53082 ( n52093,n52096,n51326 );
   nand U53083 ( n51326,n28327,n51389 );
   not U53084 ( n51389,n51656 );
   nor U53085 ( n51656,n51730,n51664 );
   not U53086 ( n52096,n52095 );
   nand U53087 ( n52095,n52097,n52098 );
   nor U53088 ( n52098,n52099,n52100 );
   nand U53089 ( n52100,n52101,n52102 );
   nor U53090 ( n52102,n52103,n52104 );
   nor U53091 ( n52104,n51934,n51336 );
   nand U53092 ( n51336,n52105,n52106 );
   nor U53093 ( n52103,n51935,n51338 );
   nand U53094 ( n51338,n52105,n52107 );
   nor U53095 ( n52101,n52108,n52109 );
   nor U53096 ( n52109,n51944,n51342 );
   nand U53097 ( n51342,n52105,n52110 );
   nor U53098 ( n52108,n51931,n51344 );
   nand U53099 ( n51344,n52105,n47399 );
   nor U53100 ( n52105,n47406,n47423 );
   nand U53101 ( n52099,n52111,n52112 );
   nor U53102 ( n52112,n52113,n52114 );
   nor U53103 ( n52114,n51923,n51350 );
   nand U53104 ( n51350,n52115,n52106 );
   nor U53105 ( n52113,n51930,n51352 );
   nand U53106 ( n51352,n52115,n52107 );
   nor U53107 ( n52111,n52116,n52117 );
   nor U53108 ( n52117,n51943,n51356 );
   nand U53109 ( n51356,n52115,n52110 );
   nor U53110 ( n52116,n51922,n51358 );
   nand U53111 ( n51358,n52115,n47399 );
   nor U53112 ( n52115,n52118,n47406 );
   nor U53113 ( n52097,n52119,n52120 );
   nand U53114 ( n52120,n52121,n52122 );
   nor U53115 ( n52122,n52123,n52124 );
   nor U53116 ( n52124,n51918,n51366 );
   nand U53117 ( n51366,n52125,n52106 );
   nor U53118 ( n52123,n51919,n51368 );
   nand U53119 ( n51368,n52125,n52107 );
   nor U53120 ( n52121,n52126,n52127 );
   nor U53121 ( n52127,n51940,n51372 );
   nand U53122 ( n51372,n52125,n52110 );
   nor U53123 ( n52126,n51913,n51374 );
   nand U53124 ( n51374,n52125,n47399 );
   nor U53125 ( n52125,n52128,n47423 );
   not U53126 ( n47423,n52118 );
   nand U53127 ( n52119,n52129,n52130 );
   nor U53128 ( n52130,n52131,n52132 );
   nor U53129 ( n52132,n51909,n51380 );
   nand U53130 ( n51380,n52133,n52106 );
   nor U53131 ( n52131,n51912,n51382 );
   nand U53132 ( n51382,n52133,n52107 );
   nor U53133 ( n52129,n52134,n52135 );
   nor U53134 ( n52135,n47308,n51385 );
   nand U53135 ( n51385,n52133,n52110 );
   nor U53136 ( n52134,n51908,n51387 );
   nand U53137 ( n51387,n52133,n47399 );
   nor U53138 ( n52133,n52118,n52128 );
   not U53139 ( n52128,n47406 );
   nand U53140 ( n47406,n52136,n52137 );
   nand U53141 ( n52137,n52138,p1_instqueuerd_addr_reg_2_ );
   nor U53142 ( n52138,n52139,n45825 );
   nand U53143 ( n52136,n52140,n50913 );
   nand U53144 ( n52140,n52139,p1_instqueuerd_addr_reg_1_ );
   xor U53145 ( n52118,p1_instqueuerd_addr_reg_2_,p1_instqueuerd_addr_reg_1_ );
   not U53146 ( n51319,n48996 );
   nor U53147 ( n48996,n52057,n48966 );
   not U53148 ( n48966,n48978 );
   nand U53149 ( n48978,n52141,n52142 );
   nor U53150 ( n52142,n52143,n52144 );
   nand U53151 ( n52144,n52145,n52146 );
   nor U53152 ( n52146,n52147,n52148 );
   nor U53153 ( n52148,n51386,n51682 );
   nand U53154 ( n51682,n52149,n52150 );
   nor U53155 ( n52147,n51379,n51683 );
   nand U53156 ( n51683,n52149,n52151 );
   nor U53157 ( n52145,n52152,n52153 );
   nor U53158 ( n52153,n51381,n51686 );
   nand U53159 ( n51686,n52149,n52154 );
   nor U53160 ( n52152,n51373,n51687 );
   nand U53161 ( n51687,n52150,n52155 );
   nand U53162 ( n52143,n52156,n52157 );
   nor U53163 ( n52157,n52158,n52159 );
   nor U53164 ( n52159,n51365,n51692 );
   nand U53165 ( n51692,n52151,n52155 );
   nor U53166 ( n52158,n51367,n51693 );
   nand U53167 ( n51693,n52154,n52155 );
   nor U53168 ( n52156,n52160,n52161 );
   nor U53169 ( n52161,n51357,n51696 );
   nand U53170 ( n51696,n52150,n52162 );
   nor U53171 ( n52160,n51349,n51697 );
   nand U53172 ( n51697,n52162,n52151 );
   nor U53173 ( n52141,n52163,n52164 );
   nand U53174 ( n52164,n52165,n52166 );
   nor U53175 ( n52166,n52167,n52168 );
   nor U53176 ( n52168,n51351,n51704 );
   nand U53177 ( n51704,n52162,n52154 );
   nor U53178 ( n52167,n51343,n51705 );
   nand U53179 ( n51705,n52169,n52150 );
   nor U53180 ( n52165,n52170,n52171 );
   nor U53181 ( n52171,n51335,n51708 );
   nand U53182 ( n51708,n52169,n52151 );
   nor U53183 ( n52170,n51337,n51709 );
   nand U53184 ( n51709,n52169,n52154 );
   nand U53185 ( n52163,n52172,n52173 );
   nor U53186 ( n52173,n52174,n52175 );
   nor U53187 ( n52175,n47243,n51714 );
   nand U53188 ( n51714,n52176,n52149 );
   nor U53189 ( n52149,n45488,n45472 );
   nor U53190 ( n52174,n51371,n51715 );
   nand U53191 ( n51715,n52176,n52155 );
   nor U53192 ( n52155,n45488,n47417 );
   nor U53193 ( n52172,n52177,n52178 );
   nor U53194 ( n52178,n51355,n51718 );
   nand U53195 ( n51718,n52176,n52162 );
   nor U53196 ( n52162,n45472,n47392 );
   not U53197 ( n45472,n47417 );
   nor U53198 ( n52177,n51341,n51719 );
   nand U53199 ( n51719,n52169,n52176 );
   nor U53200 ( n52169,n47417,n47392 );
   not U53201 ( n47392,n45488 );
   nand U53202 ( n45488,n52179,n52180 );
   or U53203 ( n52180,n50913,n52181 );
   nor U53204 ( n47417,n52182,n52183 );
   nor U53205 ( n52182,n47402,n47399 );
   not U53206 ( n50737,n50604 );
   xor U53207 ( n51318,n52184,n28185 );
   nand U53208 ( n52184,n52185,n52186 );
   nor U53209 ( n52186,n52187,n52188 );
   nor U53210 ( n52188,n28184,n48825 );
   nand U53211 ( n48825,n52189,n52190 );
   nand U53212 ( n52190,n50600,n48828 );
   not U53213 ( n50600,n52191 );
   nor U53214 ( n52187,n50604,n52192 );
   nand U53215 ( n52192,n52193,n52194 );
   nand U53216 ( n52194,n52195,n52196 );
   or U53217 ( n52195,n50605,n51313 );
   nand U53218 ( n52193,n52197,n52198 );
   not U53219 ( n52198,n52196 );
   nand U53220 ( n52196,n51189,n52199 );
   nand U53221 ( n52199,n52200,n52201 );
   nor U53222 ( n52201,n52202,n52203 );
   nand U53223 ( n52203,n52204,n52205 );
   nor U53224 ( n52205,n52206,n52207 );
   nor U53225 ( n52207,n51371,n52208 );
   nor U53226 ( n52206,n51373,n52209 );
   nor U53227 ( n52204,n52210,n52211 );
   nor U53228 ( n52211,n51365,n52212 );
   nor U53229 ( n52210,n51367,n52213 );
   nand U53230 ( n52202,n52214,n52215 );
   nor U53231 ( n52215,n52216,n52217 );
   nor U53232 ( n52217,n47243,n52218 );
   nor U53233 ( n52216,n51386,n52219 );
   nor U53234 ( n52214,n52220,n52221 );
   nor U53235 ( n52221,n51379,n52222 );
   nor U53236 ( n52220,n51381,n52223 );
   nor U53237 ( n52200,n52224,n52225 );
   nand U53238 ( n52225,n52226,n52227 );
   nor U53239 ( n52227,n52228,n52229 );
   nor U53240 ( n52229,n51341,n52230 );
   nor U53241 ( n52228,n51343,n52231 );
   nor U53242 ( n52226,n52232,n52233 );
   nor U53243 ( n52233,n51335,n52234 );
   nor U53244 ( n52232,n51337,n52235 );
   nand U53245 ( n52224,n52236,n52237 );
   nor U53246 ( n52237,n52238,n52239 );
   nor U53247 ( n52239,n51355,n52240 );
   nor U53248 ( n52238,n51357,n52241 );
   nor U53249 ( n52236,n52242,n52243 );
   nor U53250 ( n52243,n51349,n52244 );
   nor U53251 ( n52242,n51351,n52245 );
   nor U53252 ( n52197,n51313,n50605 );
   nand U53253 ( n50605,n51189,n52246 );
   nand U53254 ( n52246,n52247,n52248 );
   nor U53255 ( n52248,n52249,n52250 );
   nand U53256 ( n52250,n52251,n52252 );
   nor U53257 ( n52252,n52253,n52254 );
   nor U53258 ( n52254,n51425,n52208 );
   nor U53259 ( n52253,n51426,n52209 );
   nor U53260 ( n52251,n52255,n52256 );
   nor U53261 ( n52256,n51421,n52212 );
   nor U53262 ( n52255,n51422,n52213 );
   nand U53263 ( n52249,n52257,n52258 );
   nor U53264 ( n52258,n52259,n52260 );
   nor U53265 ( n52260,n47260,n52218 );
   nor U53266 ( n52259,n51435,n52219 );
   nor U53267 ( n52257,n52261,n52262 );
   nor U53268 ( n52262,n51431,n52222 );
   nor U53269 ( n52261,n51432,n52223 );
   nor U53270 ( n52247,n52263,n52264 );
   nand U53271 ( n52264,n52265,n52266 );
   nor U53272 ( n52266,n52267,n52268 );
   nor U53273 ( n52268,n51403,n52230 );
   nor U53274 ( n52267,n51404,n52231 );
   nor U53275 ( n52265,n52269,n52270 );
   nor U53276 ( n52270,n51399,n52234 );
   nor U53277 ( n52269,n51400,n52235 );
   nand U53278 ( n52263,n52271,n52272 );
   nor U53279 ( n52272,n52273,n52274 );
   nor U53280 ( n52274,n51413,n52240 );
   nor U53281 ( n52273,n51414,n52241 );
   nor U53282 ( n52271,n52275,n52276 );
   nor U53283 ( n52276,n51409,n52244 );
   nor U53284 ( n52275,n51410,n52245 );
   not U53285 ( n51313,n50606 );
   nor U53286 ( n50606,n51315,n51314 );
   nand U53287 ( n51314,n51189,n52277 );
   nand U53288 ( n52277,n52278,n52279 );
   nor U53289 ( n52279,n52280,n52281 );
   nand U53290 ( n52281,n52282,n52283 );
   nor U53291 ( n52283,n52284,n52285 );
   nor U53292 ( n52285,n51475,n52208 );
   nor U53293 ( n52284,n51476,n52209 );
   nor U53294 ( n52282,n52286,n52287 );
   nor U53295 ( n52287,n51471,n52212 );
   nor U53296 ( n52286,n51472,n52213 );
   nand U53297 ( n52280,n52288,n52289 );
   nor U53298 ( n52289,n52290,n52291 );
   nor U53299 ( n52291,n47276,n52218 );
   nor U53300 ( n52290,n51485,n52219 );
   nor U53301 ( n52288,n52292,n52293 );
   nor U53302 ( n52293,n51481,n52222 );
   nor U53303 ( n52292,n51482,n52223 );
   nor U53304 ( n52278,n52294,n52295 );
   nand U53305 ( n52295,n52296,n52297 );
   nor U53306 ( n52297,n52298,n52299 );
   nor U53307 ( n52299,n51453,n52230 );
   nor U53308 ( n52298,n51454,n52231 );
   nor U53309 ( n52296,n52300,n52301 );
   nor U53310 ( n52301,n51449,n52234 );
   nor U53311 ( n52300,n51450,n52235 );
   nand U53312 ( n52294,n52302,n52303 );
   nor U53313 ( n52303,n52304,n52305 );
   nor U53314 ( n52305,n51463,n52240 );
   nor U53315 ( n52304,n51464,n52241 );
   nor U53316 ( n52302,n52306,n52307 );
   nor U53317 ( n52307,n51459,n52244 );
   nor U53318 ( n52306,n51460,n52245 );
   or U53319 ( n51315,n51253,n51252 );
   nand U53320 ( n51252,n52308,n51189 );
   nand U53321 ( n52308,n52309,n52310 );
   nor U53322 ( n52310,n52311,n52312 );
   nand U53323 ( n52312,n52313,n52314 );
   nor U53324 ( n52314,n52315,n52316 );
   nor U53325 ( n52316,n51991,n52240 );
   nor U53326 ( n52315,n51970,n52241 );
   nor U53327 ( n52313,n52317,n52318 );
   nor U53328 ( n52318,n51971,n52244 );
   nor U53329 ( n52317,n51978,n52245 );
   nand U53330 ( n52311,n52319,n52320 );
   nor U53331 ( n52320,n52321,n52322 );
   nor U53332 ( n52322,n51992,n52230 );
   nor U53333 ( n52321,n51979,n52231 );
   nor U53334 ( n52319,n52323,n52324 );
   nor U53335 ( n52324,n51982,n52234 );
   nor U53336 ( n52323,n51983,n52235 );
   nor U53337 ( n52309,n52325,n52326 );
   nand U53338 ( n52326,n52327,n52328 );
   nor U53339 ( n52328,n52329,n52330 );
   nor U53340 ( n52330,n47292,n52218 );
   nor U53341 ( n52329,n51956,n52219 );
   nor U53342 ( n52327,n52331,n52332 );
   nor U53343 ( n52332,n51957,n52222 );
   nor U53344 ( n52331,n51960,n52223 );
   nand U53345 ( n52325,n52333,n52334 );
   nor U53346 ( n52334,n52335,n52336 );
   nor U53347 ( n52336,n51988,n52208 );
   nor U53348 ( n52335,n51961,n52209 );
   nor U53349 ( n52333,n52337,n52338 );
   nor U53350 ( n52338,n51966,n52212 );
   nor U53351 ( n52337,n51967,n52213 );
   or U53352 ( n51253,n51266,n51265 );
   nand U53353 ( n51265,n52339,n51189 );
   nand U53354 ( n52339,n52340,n52341 );
   nor U53355 ( n52341,n52342,n52343 );
   nand U53356 ( n52343,n52344,n52345 );
   nor U53357 ( n52345,n52346,n52347 );
   nor U53358 ( n52347,n51943,n52240 );
   nor U53359 ( n52346,n51922,n52241 );
   nor U53360 ( n52344,n52348,n52349 );
   nor U53361 ( n52349,n51923,n52244 );
   nor U53362 ( n52348,n51930,n52245 );
   nand U53363 ( n52342,n52350,n52351 );
   nor U53364 ( n52351,n52352,n52353 );
   nor U53365 ( n52353,n51944,n52230 );
   nor U53366 ( n52352,n51931,n52231 );
   nor U53367 ( n52350,n52354,n52355 );
   nor U53368 ( n52355,n51934,n52234 );
   nor U53369 ( n52354,n51935,n52235 );
   nor U53370 ( n52340,n52356,n52357 );
   nand U53371 ( n52357,n52358,n52359 );
   nor U53372 ( n52359,n52360,n52361 );
   nor U53373 ( n52361,n47308,n52218 );
   nor U53374 ( n52360,n51908,n52219 );
   nor U53375 ( n52358,n52362,n52363 );
   nor U53376 ( n52363,n51909,n52222 );
   nor U53377 ( n52362,n51912,n52223 );
   nand U53378 ( n52356,n52364,n52365 );
   nor U53379 ( n52365,n52366,n52367 );
   nor U53380 ( n52367,n51940,n52208 );
   nor U53381 ( n52366,n51913,n52209 );
   nor U53382 ( n52364,n52368,n52369 );
   nor U53383 ( n52369,n51918,n52212 );
   nor U53384 ( n52368,n51919,n52213 );
   or U53385 ( n51266,n51291,n51290 );
   nand U53386 ( n51290,n52370,n51189 );
   nand U53387 ( n52370,n52371,n52372 );
   nor U53388 ( n52372,n52373,n52374 );
   nand U53389 ( n52374,n52375,n52376 );
   nor U53390 ( n52376,n52377,n52378 );
   nor U53391 ( n52378,n51514,n52240 );
   nor U53392 ( n52377,n51515,n52241 );
   nor U53393 ( n52375,n52379,n52380 );
   nor U53394 ( n52380,n51510,n52244 );
   nor U53395 ( n52379,n51511,n52245 );
   nand U53396 ( n52373,n52381,n52382 );
   nor U53397 ( n52382,n52383,n52384 );
   nor U53398 ( n52384,n51504,n52230 );
   nor U53399 ( n52383,n51505,n52231 );
   nor U53400 ( n52381,n52385,n52386 );
   nor U53401 ( n52386,n51500,n52234 );
   nor U53402 ( n52385,n51501,n52235 );
   nor U53403 ( n52371,n52387,n52388 );
   nand U53404 ( n52388,n52389,n52390 );
   nor U53405 ( n52390,n52391,n52392 );
   nor U53406 ( n52392,n47323,n52218 );
   nor U53407 ( n52391,n51536,n52219 );
   nor U53408 ( n52389,n52393,n52394 );
   nor U53409 ( n52394,n51532,n52222 );
   nor U53410 ( n52393,n51533,n52223 );
   nand U53411 ( n52387,n52395,n52396 );
   nor U53412 ( n52396,n52397,n52398 );
   nor U53413 ( n52398,n51526,n52208 );
   nor U53414 ( n52397,n51527,n52209 );
   nor U53415 ( n52395,n52399,n52400 );
   nor U53416 ( n52400,n51522,n52212 );
   nor U53417 ( n52399,n51523,n52213 );
   or U53418 ( n51291,n51302,n51301 );
   nand U53419 ( n51301,n52401,n51189 );
   nand U53420 ( n52401,n52402,n52403 );
   nor U53421 ( n52403,n52404,n52405 );
   nand U53422 ( n52405,n52406,n52407 );
   nor U53423 ( n52407,n52408,n52409 );
   nor U53424 ( n52409,n51564,n52240 );
   nor U53425 ( n52408,n51565,n52241 );
   nor U53426 ( n52406,n52410,n52411 );
   nor U53427 ( n52411,n51560,n52244 );
   nor U53428 ( n52410,n51561,n52245 );
   nand U53429 ( n52404,n52412,n52413 );
   nor U53430 ( n52413,n52414,n52415 );
   nor U53431 ( n52415,n51554,n52230 );
   nor U53432 ( n52414,n51555,n52231 );
   nor U53433 ( n52412,n52416,n52417 );
   nor U53434 ( n52417,n51550,n52234 );
   nor U53435 ( n52416,n51551,n52235 );
   nor U53436 ( n52402,n52418,n52419 );
   nand U53437 ( n52419,n52420,n52421 );
   nor U53438 ( n52421,n52422,n52423 );
   nor U53439 ( n52423,n47339,n52218 );
   nor U53440 ( n52422,n51586,n52219 );
   nor U53441 ( n52420,n52424,n52425 );
   nor U53442 ( n52425,n51582,n52222 );
   nor U53443 ( n52424,n51583,n52223 );
   nand U53444 ( n52418,n52426,n52427 );
   nor U53445 ( n52427,n52428,n52429 );
   nor U53446 ( n52429,n51576,n52208 );
   nor U53447 ( n52428,n51577,n52209 );
   nor U53448 ( n52426,n52430,n52431 );
   nor U53449 ( n52431,n51572,n52212 );
   nor U53450 ( n52430,n51573,n52213 );
   or U53451 ( n51302,n51278,n51279 );
   nand U53452 ( n51279,n51189,n52432 );
   nand U53453 ( n52432,n52433,n52434 );
   nor U53454 ( n52434,n52435,n52436 );
   nand U53455 ( n52436,n52437,n52438 );
   nor U53456 ( n52438,n52439,n52440 );
   nor U53457 ( n52440,n51626,n52208 );
   nand U53458 ( n52208,n52441,n52442 );
   nor U53459 ( n52439,n51627,n52209 );
   nand U53460 ( n52209,n52443,n52441 );
   nor U53461 ( n52443,p1_instqueuerd_addr_reg_2_,n52444 );
   nor U53462 ( n52437,n52445,n52446 );
   nor U53463 ( n52446,n51622,n52212 );
   nand U53464 ( n52212,n52447,n52441 );
   nor U53465 ( n52447,p1_instqueuerd_addr_reg_2_,n52448 );
   nor U53466 ( n52445,n51623,n52213 );
   nand U53467 ( n52213,n52441,n52183 );
   nand U53468 ( n52435,n52449,n52450 );
   nor U53469 ( n52450,n52451,n52452 );
   nor U53470 ( n52452,n47364,n52218 );
   nand U53471 ( n52218,n52441,n52453 );
   nor U53472 ( n52451,n51636,n52219 );
   nand U53473 ( n52219,n52441,n52454 );
   nor U53474 ( n52449,n52455,n52456 );
   nor U53475 ( n52456,n51632,n52222 );
   nand U53476 ( n52222,n52441,n52457 );
   nor U53477 ( n52455,n51633,n52223 );
   nand U53478 ( n52223,n52441,n52181 );
   nor U53479 ( n52433,n52458,n52459 );
   nand U53480 ( n52459,n52460,n52461 );
   nor U53481 ( n52461,n52462,n52463 );
   nor U53482 ( n52463,n51604,n52230 );
   nand U53483 ( n52230,n52442,n52464 );
   nor U53484 ( n52462,n51605,n52231 );
   nand U53485 ( n52231,n52465,n52107 );
   nor U53486 ( n52460,n52466,n52467 );
   nor U53487 ( n52467,n51600,n52234 );
   nand U53488 ( n52234,n52465,n52110 );
   nor U53489 ( n52465,p1_instqueuerd_addr_reg_2_,n52441 );
   nor U53490 ( n52466,n51601,n52235 );
   nand U53491 ( n52235,n52183,n52464 );
   nand U53492 ( n52458,n52468,n52469 );
   nor U53493 ( n52469,n52470,n52471 );
   nor U53494 ( n52471,n51614,n52240 );
   nand U53495 ( n52240,n52453,n52464 );
   nor U53496 ( n52470,n51615,n52241 );
   nand U53497 ( n52241,n52454,n52464 );
   nor U53498 ( n52468,n52472,n52473 );
   nor U53499 ( n52473,n51610,n52244 );
   nand U53500 ( n52244,n52457,n52464 );
   nor U53501 ( n52472,n51611,n52245 );
   nand U53502 ( n52245,n52181,n52464 );
   not U53503 ( n52464,n52441 );
   nor U53504 ( n52441,n52474,n52139 );
   nand U53505 ( n51278,n51189,n52475 );
   nand U53506 ( n52475,n52476,n52477 );
   nor U53507 ( n52477,n52478,n52479 );
   nand U53508 ( n52479,n52480,n52481 );
   nor U53509 ( n52481,n52482,n52483 );
   nor U53510 ( n52483,n51371,n51203 );
   nand U53511 ( n51203,n52484,n52151 );
   nor U53512 ( n52482,n51373,n51202 );
   nand U53513 ( n51202,n52484,n52154 );
   nor U53514 ( n52480,n52485,n52486 );
   nor U53515 ( n52486,n51365,n51199 );
   nand U53516 ( n51199,n52484,n52176 );
   nor U53517 ( n52485,n51367,n51198 );
   nand U53518 ( n51198,n52484,n52150 );
   nor U53519 ( n52484,n52487,n52488 );
   nand U53520 ( n52478,n52489,n52490 );
   nor U53521 ( n52490,n52491,n52492 );
   nor U53522 ( n52492,n47243,n51213 );
   nand U53523 ( n51213,n52493,n52151 );
   nor U53524 ( n52491,n51386,n51212 );
   nand U53525 ( n51212,n52493,n52154 );
   nor U53526 ( n52489,n52494,n52495 );
   nor U53527 ( n52495,n51379,n51209 );
   nand U53528 ( n51209,n52493,n52176 );
   nor U53529 ( n52494,n51381,n51208 );
   nand U53530 ( n51208,n52493,n52150 );
   nor U53531 ( n52493,n52487,n52496 );
   nor U53532 ( n52476,n52497,n52498 );
   nand U53533 ( n52498,n52499,n52500 );
   nor U53534 ( n52500,n52501,n52502 );
   nor U53535 ( n52502,n51341,n51225 );
   nand U53536 ( n51225,n52503,n52151 );
   nor U53537 ( n52501,n51343,n51224 );
   nand U53538 ( n51224,n52503,n52154 );
   nor U53539 ( n52499,n52504,n52505 );
   nor U53540 ( n52505,n51335,n51221 );
   nand U53541 ( n51221,n52503,n52176 );
   nor U53542 ( n52504,n51337,n51220 );
   nand U53543 ( n51220,n52503,n52150 );
   nor U53544 ( n52503,n52488,n52506 );
   not U53545 ( n52488,n52496 );
   nand U53546 ( n52497,n52507,n52508 );
   nor U53547 ( n52508,n52509,n52510 );
   nor U53548 ( n52510,n51355,n51235 );
   nand U53549 ( n51235,n52511,n52151 );
   nor U53550 ( n52151,n52512,n45451 );
   nor U53551 ( n52509,n51357,n51234 );
   nand U53552 ( n51234,n52511,n52154 );
   nor U53553 ( n52154,n52512,p1_instqueuerd_addr_reg_0_ );
   not U53554 ( n52512,n45460 );
   nor U53555 ( n52507,n52513,n52514 );
   nor U53556 ( n52514,n51349,n51231 );
   nand U53557 ( n51231,n52511,n52176 );
   nor U53558 ( n52176,n45451,n45460 );
   nor U53559 ( n52513,n51351,n51230 );
   nand U53560 ( n51230,n52511,n52150 );
   nor U53561 ( n52150,n45460,p1_instqueuerd_addr_reg_0_ );
   nor U53562 ( n45460,n47399,n52106 );
   nor U53563 ( n52511,n52506,n52496 );
   nor U53564 ( n52496,n52515,n52442 );
   not U53565 ( n52506,n52487 );
   nand U53566 ( n52487,n52516,n52517 );
   or U53567 ( n52517,n50913,n52515 );
   nor U53568 ( n52515,n47402,n52106 );
   nand U53569 ( n52516,n52139,n47407 );
   nand U53570 ( n51189,n52518,n52519 );
   nand U53571 ( n52519,n47416,p1_state2_reg_0_ );
   not U53572 ( n47416,n45851 );
   nand U53573 ( n45851,n52520,n45329 );
   and U53574 ( n52520,n47351,n45853 );
   nand U53575 ( n52518,n49622,n45853 );
   nor U53576 ( n45853,n47420,n45878 );
   nand U53577 ( n47420,n52521,n49431 );
   nor U53578 ( n49431,n47255,n49602 );
   nor U53579 ( n52521,n48247,n47426 );
   nand U53580 ( n50604,p1_state2_reg_2_,n52522 );
   nand U53581 ( n52522,n48289,n47255 );
   nor U53582 ( n52185,n52523,n52524 );
   nor U53583 ( n52524,n50609,n49327 );
   not U53584 ( n49327,p1_eax_reg_30_ );
   not U53585 ( n50609,n50593 );
   nor U53586 ( n50593,n47236,n28375 );
   nor U53587 ( n52523,n50610,n48828 );
   not U53588 ( n48828,p1_phyaddrpointer_reg_30_ );
   not U53589 ( n50610,n49013 );
   nor U53590 ( n49013,n47377,p1_state2_reg_2_ );
   not U53591 ( n50010,n49979 );
   nand U53592 ( n49979,n52525,p1_state2_reg_1_ );
   nor U53593 ( n52525,n50566,n49010 );
   xor U53594 ( n49010,p1_phyaddrpointer_reg_31_,n52189 );
   nand U53595 ( n52189,p1_phyaddrpointer_reg_30_,n52191 );
   nor U53596 ( n52191,n48802,n50602 );
   or U53597 ( n50602,n48787,n51310 );
   nand U53598 ( n51310,n52526,p1_phyaddrpointer_reg_27_ );
   not U53599 ( n52526,n51254 );
   nand U53600 ( n51254,n52527,p1_phyaddrpointer_reg_26_ );
   nor U53601 ( n52527,n48727,n51298 );
   not U53602 ( n51298,n51262 );
   nor U53603 ( n51262,n48708,n51275 );
   or U53604 ( n51275,n48694,n51066 );
   nand U53605 ( n51066,n52528,p1_phyaddrpointer_reg_22_ );
   nor U53606 ( n52528,n48655,n51187 );
   not U53607 ( n51187,n51068 );
   nor U53608 ( n51068,n48635,n51108 );
   or U53609 ( n51108,n48620,n50638 );
   nand U53610 ( n50638,n52529,p1_phyaddrpointer_reg_18_ );
   nor U53611 ( n52529,n48587,n51024 );
   not U53612 ( n51024,n50640 );
   nor U53613 ( n50640,n48572,n50742 );
   or U53614 ( n50742,n48551,n50744 );
   nand U53615 ( n50744,n52530,p1_phyaddrpointer_reg_14_ );
   nor U53616 ( n52530,n48511,n50761 );
   nand U53617 ( n50761,n52531,p1_phyaddrpointer_reg_12_ );
   nor U53618 ( n52531,n48481,n50792 );
   nand U53619 ( n50792,n52532,p1_phyaddrpointer_reg_10_ );
   nor U53620 ( n52532,n48445,n50809 );
   nand U53621 ( n50809,n52533,p1_phyaddrpointer_reg_8_ );
   nor U53622 ( n52533,n48411,n50825 );
   nand U53623 ( n50825,n52534,p1_phyaddrpointer_reg_6_ );
   nor U53624 ( n52534,n48377,n50932 );
   nand U53625 ( n50932,n52535,p1_phyaddrpointer_reg_4_ );
   nor U53626 ( n52535,n48349,n50890 );
   nand U53627 ( n50890,p1_phyaddrpointer_reg_2_,p1_phyaddrpointer_reg_1_ );
   not U53628 ( n48349,p1_phyaddrpointer_reg_3_ );
   not U53629 ( n48377,p1_phyaddrpointer_reg_5_ );
   not U53630 ( n48411,p1_phyaddrpointer_reg_7_ );
   not U53631 ( n48445,p1_phyaddrpointer_reg_9_ );
   not U53632 ( n48481,p1_phyaddrpointer_reg_11_ );
   not U53633 ( n48511,p1_phyaddrpointer_reg_13_ );
   not U53634 ( n48551,p1_phyaddrpointer_reg_15_ );
   not U53635 ( n48572,p1_phyaddrpointer_reg_16_ );
   not U53636 ( n48587,p1_phyaddrpointer_reg_17_ );
   not U53637 ( n48620,p1_phyaddrpointer_reg_19_ );
   not U53638 ( n48635,p1_phyaddrpointer_reg_20_ );
   not U53639 ( n48655,p1_phyaddrpointer_reg_21_ );
   not U53640 ( n48694,p1_phyaddrpointer_reg_23_ );
   not U53641 ( n48708,p1_phyaddrpointer_reg_24_ );
   not U53642 ( n48727,p1_phyaddrpointer_reg_25_ );
   not U53643 ( n48787,p1_phyaddrpointer_reg_28_ );
   not U53644 ( n48802,p1_phyaddrpointer_reg_29_ );
   nand U53645 ( n50579,n28286,n49823 );
   not U53646 ( n49823,n48244 );
   xor U53647 ( n48244,n52536,n52537 );
   nand U53648 ( n52537,n50563,n50564 );
   xor U53649 ( n50564,n45329,n52538 );
   nand U53650 ( n52538,n52539,n52540 );
   nand U53651 ( n52540,p1_ebx_reg_30_,n28342 );
   nand U53652 ( n52539,p1_instaddrpointer_reg_30_,n28276 );
   nor U53653 ( n50563,n50526,n50546 );
   xor U53654 ( n50546,n28404,n52541 );
   nand U53655 ( n52541,n52542,n52543 );
   nand U53656 ( n52543,p1_ebx_reg_29_,n49852 );
   nand U53657 ( n52542,p1_instaddrpointer_reg_29_,n49870 );
   or U53658 ( n50526,n50528,n50527 );
   xor U53659 ( n50527,n28403,n52544 );
   nand U53660 ( n52544,n52545,n52546 );
   nand U53661 ( n52546,p1_ebx_reg_28_,n28342 );
   nand U53662 ( n52545,p1_instaddrpointer_reg_28_,n28276 );
   or U53663 ( n50528,n50482,n50503 );
   xor U53664 ( n50503,n28406,n52547 );
   nand U53665 ( n52547,n52548,n52549 );
   nand U53666 ( n52549,p1_ebx_reg_27_,n49852 );
   nand U53667 ( n52548,p1_instaddrpointer_reg_27_,n28276 );
   or U53668 ( n50482,n50484,n50483 );
   xor U53669 ( n50483,n28403,n52550 );
   nand U53670 ( n52550,n52551,n52552 );
   nand U53671 ( n52552,p1_ebx_reg_26_,n49852 );
   nand U53672 ( n52551,p1_instaddrpointer_reg_26_,n49870 );
   or U53673 ( n50484,n50435,n50455 );
   xor U53674 ( n50455,n28404,n52553 );
   nand U53675 ( n52553,n52554,n52555 );
   nand U53676 ( n52555,p1_ebx_reg_25_,n49852 );
   nand U53677 ( n52554,p1_instaddrpointer_reg_25_,n28276 );
   or U53678 ( n50435,n50437,n50436 );
   xor U53679 ( n50436,n28404,n52556 );
   nand U53680 ( n52556,n52557,n52558 );
   nand U53681 ( n52558,p1_ebx_reg_24_,n49852 );
   nand U53682 ( n52557,p1_instaddrpointer_reg_24_,n28276 );
   or U53683 ( n50437,n50392,n50412 );
   xor U53684 ( n50412,n28405,n52559 );
   nand U53685 ( n52559,n52560,n52561 );
   nand U53686 ( n52561,p1_ebx_reg_23_,n49852 );
   nand U53687 ( n52560,p1_instaddrpointer_reg_23_,n28276 );
   or U53688 ( n50392,n50394,n50393 );
   xor U53689 ( n50393,n28405,n52562 );
   nand U53690 ( n52562,n52563,n52564 );
   nand U53691 ( n52564,p1_ebx_reg_22_,n49852 );
   nand U53692 ( n52563,p1_instaddrpointer_reg_22_,n49870 );
   or U53693 ( n50394,n50343,n50363 );
   xor U53694 ( n50363,n28403,n52565 );
   nand U53695 ( n52565,n52566,n52567 );
   nand U53696 ( n52567,p1_ebx_reg_21_,n49852 );
   nand U53697 ( n52566,p1_instaddrpointer_reg_21_,n49870 );
   or U53698 ( n50343,n50345,n50344 );
   xor U53699 ( n50344,n28405,n52568 );
   nand U53700 ( n52568,n52569,n52570 );
   nand U53701 ( n52570,p1_ebx_reg_20_,n49852 );
   nand U53702 ( n52569,p1_instaddrpointer_reg_20_,n49870 );
   or U53703 ( n50345,n50296,n50317 );
   xor U53704 ( n50317,n28403,n52571 );
   nand U53705 ( n52571,n52572,n52573 );
   nand U53706 ( n52573,p1_ebx_reg_19_,n49852 );
   nand U53707 ( n52572,p1_instaddrpointer_reg_19_,n49870 );
   or U53708 ( n50296,n50298,n50297 );
   xor U53709 ( n50297,n28406,n52574 );
   nand U53710 ( n52574,n52575,n52576 );
   nand U53711 ( n52576,p1_ebx_reg_18_,n49852 );
   nand U53712 ( n52575,p1_instaddrpointer_reg_18_,n49870 );
   or U53713 ( n50298,n50248,n50271 );
   xor U53714 ( n50271,n28405,n52577 );
   nand U53715 ( n52577,n52578,n52579 );
   nand U53716 ( n52579,p1_ebx_reg_17_,n49852 );
   nand U53717 ( n52578,p1_instaddrpointer_reg_17_,n49870 );
   or U53718 ( n50248,n50250,n50249 );
   xor U53719 ( n50249,n28405,n52580 );
   nand U53720 ( n52580,n52581,n52582 );
   nand U53721 ( n52582,p1_ebx_reg_16_,n49852 );
   nand U53722 ( n52581,p1_instaddrpointer_reg_16_,n28276 );
   or U53723 ( n50250,n50200,n50225 );
   xor U53724 ( n50225,n28404,n52583 );
   nand U53725 ( n52583,n52584,n52585 );
   nand U53726 ( n52585,p1_ebx_reg_15_,n49852 );
   nand U53727 ( n52584,p1_instaddrpointer_reg_15_,n49870 );
   or U53728 ( n50200,n50202,n50201 );
   xor U53729 ( n50201,n28404,n52586 );
   nand U53730 ( n52586,n52587,n52588 );
   nand U53731 ( n52588,p1_ebx_reg_14_,n49852 );
   nand U53732 ( n52587,p1_instaddrpointer_reg_14_,n49870 );
   or U53733 ( n50202,n50153,n50175 );
   xor U53734 ( n50175,n28406,n52589 );
   nand U53735 ( n52589,n52590,n52591 );
   nand U53736 ( n52591,p1_ebx_reg_13_,n49852 );
   nand U53737 ( n52590,p1_instaddrpointer_reg_13_,n49870 );
   or U53738 ( n50153,n50155,n50154 );
   xor U53739 ( n50154,n28404,n52592 );
   nand U53740 ( n52592,n52593,n52594 );
   nand U53741 ( n52594,p1_ebx_reg_12_,n49852 );
   nand U53742 ( n52593,p1_instaddrpointer_reg_12_,n49870 );
   or U53743 ( n50155,n50101,n50125 );
   xor U53744 ( n50125,n28406,n52595 );
   nand U53745 ( n52595,n52596,n52597 );
   nand U53746 ( n52597,p1_ebx_reg_11_,n28342 );
   nand U53747 ( n52596,p1_instaddrpointer_reg_11_,n28276 );
   or U53748 ( n50101,n50103,n50102 );
   xor U53749 ( n50102,n28403,n52598 );
   nand U53750 ( n52598,n52599,n52600 );
   nand U53751 ( n52600,p1_ebx_reg_10_,n28342 );
   nand U53752 ( n52599,p1_instaddrpointer_reg_10_,n49870 );
   or U53753 ( n50103,n50054,n50076 );
   xor U53754 ( n50076,n28404,n52601 );
   nand U53755 ( n52601,n52602,n52603 );
   nand U53756 ( n52603,p1_ebx_reg_9_,n28342 );
   nand U53757 ( n52602,p1_instaddrpointer_reg_9_,n49870 );
   or U53758 ( n50054,n50056,n50055 );
   xor U53759 ( n50055,n28405,n52604 );
   nand U53760 ( n52604,n52605,n52606 );
   nand U53761 ( n52606,p1_ebx_reg_8_,n28342 );
   nand U53762 ( n52605,p1_instaddrpointer_reg_8_,n49870 );
   or U53763 ( n50056,n50005,n50031 );
   xor U53764 ( n50031,n28405,n52607 );
   nand U53765 ( n52607,n52608,n52609 );
   nand U53766 ( n52609,p1_ebx_reg_7_,n28342 );
   nand U53767 ( n52608,p1_instaddrpointer_reg_7_,n49870 );
   or U53768 ( n50005,n50007,n50006 );
   xor U53769 ( n50006,n28403,n52610 );
   nand U53770 ( n52610,n52611,n52612 );
   nand U53771 ( n52612,p1_ebx_reg_6_,n28342 );
   nand U53772 ( n52611,p1_instaddrpointer_reg_6_,n49870 );
   or U53773 ( n50007,n49948,n49977 );
   xor U53774 ( n49977,n28403,n52613 );
   nand U53775 ( n52613,n52614,n52615 );
   nand U53776 ( n52615,p1_ebx_reg_5_,n28342 );
   nand U53777 ( n52614,p1_instaddrpointer_reg_5_,n49870 );
   or U53778 ( n49948,n49950,n49949 );
   xor U53779 ( n49949,n28406,n52616 );
   nand U53780 ( n52616,n52617,n52618 );
   nand U53781 ( n52618,p1_ebx_reg_4_,n28342 );
   nand U53782 ( n52617,p1_instaddrpointer_reg_4_,n49870 );
   nand U53783 ( n49950,n49926,n49927 );
   xor U53784 ( n49927,n45329,n52619 );
   nand U53785 ( n52619,n52620,n52621 );
   nand U53786 ( n52621,p1_ebx_reg_3_,n28342 );
   nand U53787 ( n52620,p1_instaddrpointer_reg_3_,n49870 );
   nor U53788 ( n49926,n49902,n49901 );
   xor U53789 ( n49901,n28406,n52622 );
   nand U53790 ( n52622,n52623,n52624 );
   nand U53791 ( n52624,p1_ebx_reg_2_,n28342 );
   nand U53792 ( n52623,p1_instaddrpointer_reg_2_,n28276 );
   not U53793 ( n49870,n52625 );
   nand U53794 ( n49902,n52626,n52627 );
   nand U53795 ( n52627,n52628,n52625 );
   or U53796 ( n52628,n49868,n49871 );
   nand U53797 ( n52626,n49868,n49871 );
   nand U53798 ( n49871,n49853,n28342 );
   xor U53799 ( n49853,n52629,n28406 );
   nor U53800 ( n52629,n52630,n52631 );
   nor U53801 ( n52631,n45448,n52625 );
   not U53802 ( n45448,p1_instaddrpointer_reg_0_ );
   nor U53803 ( n52630,n52632,n49855 );
   not U53804 ( n49855,p1_ebx_reg_0_ );
   xor U53805 ( n49868,n52633,n45329 );
   nor U53806 ( n52633,n52634,n52635 );
   nor U53807 ( n52635,n45479,n52625 );
   not U53808 ( n45479,p1_instaddrpointer_reg_1_ );
   and U53809 ( n52634,n49852,p1_ebx_reg_1_ );
   not U53810 ( n49852,n52632 );
   nor U53811 ( n52536,n45329,n52636 );
   nor U53812 ( n52636,n52637,n52638 );
   nor U53813 ( n52638,n45480,n52625 );
   nand U53814 ( n52625,n49620,n52639 );
   nand U53815 ( n52639,n51880,n47351 );
   not U53816 ( n45480,p1_instaddrpointer_reg_31_ );
   nor U53817 ( n52637,n52632,n52640 );
   nor U53818 ( n52632,n45329,n48210 );
   nor U53819 ( n48210,n47303,n45876 );
   nor U53820 ( n45329,n45877,n48289 );
   and U53821 ( n49851,n52641,n52642 );
   nor U53822 ( n52642,n52643,n49620 );
   and U53823 ( n52641,p1_ebx_reg_31_,n49952 );
   nor U53824 ( n50577,n49016,n49837 );
   not U53825 ( n49837,n49883 );
   nor U53826 ( n49883,n45501,n50566 );
   not U53827 ( n49016,p1_phyaddrpointer_reg_31_ );
   nor U53828 ( n50575,n52644,n52645 );
   nand U53829 ( n52645,n52646,n52647 );
   nand U53830 ( n52647,p1_reip_reg_31_,n52648 );
   nand U53831 ( n52648,n52649,n52650 );
   nand U53832 ( n52650,n28140,n45529 );
   not U53833 ( n45529,p1_reip_reg_30_ );
   not U53834 ( n52649,n50573 );
   nand U53835 ( n50573,n50554,n52651 );
   nand U53836 ( n52651,n28140,n45534 );
   not U53837 ( n45534,p1_reip_reg_29_ );
   nor U53838 ( n50554,n50535,n52652 );
   nor U53839 ( n52652,n49841,p1_reip_reg_28_ );
   nand U53840 ( n50535,n49840,n52653 );
   nand U53841 ( n52653,n28141,n50537 );
   not U53842 ( n50537,n52654 );
   nand U53843 ( n52646,n52655,n45527 );
   not U53844 ( n45527,p1_reip_reg_31_ );
   nor U53845 ( n52655,n50553,n52656 );
   nand U53846 ( n52656,p1_reip_reg_29_,p1_reip_reg_30_ );
   nand U53847 ( n50553,n52657,n52654 );
   nor U53848 ( n52654,n52658,n50493 );
   nand U53849 ( n50493,n52659,n50468 );
   nor U53850 ( n50468,n52660,n50403 );
   nand U53851 ( n50403,n52661,n50376 );
   nor U53852 ( n50376,n52662,n50310 );
   nand U53853 ( n50310,n52663,n50287 );
   nor U53854 ( n50287,n52664,n50218 );
   nand U53855 ( n50218,n52665,n50191 );
   nor U53856 ( n50191,n52666,n50118 );
   nand U53857 ( n50118,n52667,n50092 );
   nor U53858 ( n50092,n52668,n50024 );
   nand U53859 ( n50024,n52669,n49966 );
   not U53860 ( n49966,n49994 );
   nand U53861 ( n49994,n52670,p1_reip_reg_2_ );
   nor U53862 ( n52670,n45674,n45664 );
   not U53863 ( n45664,p1_reip_reg_3_ );
   nor U53864 ( n52669,n45654,n45659 );
   not U53865 ( n45659,p1_reip_reg_4_ );
   not U53866 ( n45654,p1_reip_reg_5_ );
   nand U53867 ( n52668,p1_reip_reg_7_,p1_reip_reg_6_ );
   nor U53868 ( n52667,n45634,n45639 );
   not U53869 ( n45639,p1_reip_reg_8_ );
   not U53870 ( n45634,p1_reip_reg_9_ );
   nand U53871 ( n52666,p1_reip_reg_11_,p1_reip_reg_10_ );
   nor U53872 ( n52665,n45614,n45619 );
   not U53873 ( n45619,p1_reip_reg_12_ );
   not U53874 ( n45614,p1_reip_reg_13_ );
   nand U53875 ( n52664,p1_reip_reg_15_,p1_reip_reg_14_ );
   nor U53876 ( n52663,n45594,n45599 );
   not U53877 ( n45599,p1_reip_reg_16_ );
   not U53878 ( n45594,p1_reip_reg_17_ );
   nand U53879 ( n52662,p1_reip_reg_19_,p1_reip_reg_18_ );
   nor U53880 ( n52661,n45574,n45579 );
   not U53881 ( n45579,p1_reip_reg_20_ );
   not U53882 ( n45574,p1_reip_reg_21_ );
   nand U53883 ( n52660,p1_reip_reg_23_,p1_reip_reg_22_ );
   nor U53884 ( n52659,n45554,n45559 );
   not U53885 ( n45559,p1_reip_reg_24_ );
   not U53886 ( n45554,p1_reip_reg_25_ );
   nand U53887 ( n52658,p1_reip_reg_27_,p1_reip_reg_26_ );
   nor U53888 ( n52657,n45539,n28250 );
   nand U53889 ( n49841,n52671,n49952 );
   nor U53890 ( n52671,n52672,n52673 );
   not U53891 ( n52673,n52643 );
   nor U53892 ( n52672,n52674,n51878 );
   nor U53893 ( n52674,n45351,n48912 );
   not U53894 ( n48912,n45358 );
   not U53895 ( n45539,p1_reip_reg_28_ );
   nor U53896 ( n52644,n52640,n49856 );
   nand U53897 ( n49856,n49952,n52675 );
   nand U53898 ( n52675,n52676,n52677 );
   nand U53899 ( n52677,n52678,n51878 );
   nor U53900 ( n52678,p1_ebx_reg_31_,n52643 );
   nand U53901 ( n52676,n45358,n45795 );
   nand U53902 ( n45795,n52643,n45360 );
   nor U53903 ( n52643,p1_statebs16_reg,n45701 );
   not U53904 ( n45701,n45346 );
   nor U53905 ( n49952,n28374,n50566 );
   not U53906 ( n50566,n49840 );
   nand U53907 ( n49840,n52679,n52680 );
   nor U53908 ( n52680,n52681,n45767 );
   and U53909 ( n45767,n52682,n28407 );
   nor U53910 ( n49843,p1_state2_reg_2_,p1_statebs16_reg );
   nor U53911 ( n52682,p1_state2_reg_0_,n45432 );
   not U53912 ( n52681,n45777 );
   nand U53913 ( n45777,n52683,n45352 );
   nor U53914 ( n45352,p1_state2_reg_1_,p1_state2_reg_2_ );
   nor U53915 ( n52683,n45347,n45501 );
   not U53916 ( n45501,p1_state2_reg_3_ );
   nor U53917 ( n52679,n45325,n48272 );
   nor U53918 ( n48272,p1_state2_reg_2_,n49019 );
   not U53919 ( n49019,n45342 );
   nor U53920 ( n45342,n45464,p1_state2_reg_0_ );
   not U53921 ( n45464,n45443 );
   nor U53922 ( n45443,p1_state2_reg_1_,p1_state2_reg_3_ );
   and U53923 ( n45325,n45759,n52684 );
   nand U53924 ( n52684,n52685,n52686 );
   nand U53925 ( n52686,n51860,n48279 );
   nor U53926 ( n51860,n47429,n28095 );
   nand U53927 ( n47429,n45328,n49630 );
   nor U53928 ( n52685,n52687,n52688 );
   nor U53929 ( n52688,n45836,n52689 );
   nand U53930 ( n52689,p1_state2_reg_0_,n45869 );
   nand U53931 ( n45836,n49951,n49630 );
   nor U53932 ( n49951,n48289,n47351 );
   not U53933 ( n52640,p1_ebx_reg_31_ );
   nor U53934 ( n52690,n52692,n52693 );
   nor U53935 ( n52693,n45372,n52694 );
   or U53936 ( n52694,p1_datawidth_reg_1_,p1_reip_reg_1_ );
   and U53937 ( n52692,n45372,p1_byteenable_reg_3_ );
   nand U53938 ( n52696,p1_byteenable_reg_1_,n45372 );
   and U53939 ( n52695,n52691,n45369 );
   not U53940 ( n45369,n45376 );
   nor U53941 ( n45376,n45674,n45372 );
   not U53942 ( n45674,p1_reip_reg_1_ );
   nand U53943 ( n52691,n52697,n52698 );
   nor U53944 ( n52698,p1_reip_reg_0_,p1_datawidth_reg_1_ );
   nor U53945 ( n52697,p1_datawidth_reg_0_,n45372 );
   nand U53946 ( n45372,n52699,n52700 );
   nor U53947 ( n52700,n52701,n52702 );
   nand U53948 ( n52702,n52703,n52704 );
   nor U53949 ( n52704,n52705,n52706 );
   nand U53950 ( n52706,n45748,n45749 );
   not U53951 ( n45749,p1_datawidth_reg_29_ );
   not U53952 ( n45748,p1_datawidth_reg_28_ );
   nand U53953 ( n52705,n45722,n45750 );
   not U53954 ( n45750,p1_datawidth_reg_30_ );
   not U53955 ( n45722,p1_datawidth_reg_2_ );
   nor U53956 ( n52703,n52707,n52708 );
   nand U53957 ( n52708,n45744,n45745 );
   not U53958 ( n45745,p1_datawidth_reg_25_ );
   not U53959 ( n45744,p1_datawidth_reg_24_ );
   nand U53960 ( n52707,n45746,n45747 );
   not U53961 ( n45747,p1_datawidth_reg_27_ );
   not U53962 ( n45746,p1_datawidth_reg_26_ );
   nand U53963 ( n52701,n52709,n52710 );
   nor U53964 ( n52710,n52711,n52712 );
   nand U53965 ( n52712,n45726,n45727 );
   not U53966 ( n45727,p1_datawidth_reg_7_ );
   not U53967 ( n45726,p1_datawidth_reg_6_ );
   nand U53968 ( n52711,n45728,n45729 );
   not U53969 ( n45729,p1_datawidth_reg_9_ );
   not U53970 ( n45728,p1_datawidth_reg_8_ );
   nor U53971 ( n52709,n52713,n52714 );
   nand U53972 ( n52714,n45751,n45723 );
   not U53973 ( n45723,p1_datawidth_reg_3_ );
   not U53974 ( n45751,p1_datawidth_reg_31_ );
   nand U53975 ( n52713,n45724,n45725 );
   not U53976 ( n45725,p1_datawidth_reg_5_ );
   not U53977 ( n45724,p1_datawidth_reg_4_ );
   nor U53978 ( n52699,n52715,n52716 );
   nand U53979 ( n52716,n52717,n52718 );
   nor U53980 ( n52718,n52719,n52720 );
   nand U53981 ( n52720,n45732,n45733 );
   not U53982 ( n45733,p1_datawidth_reg_13_ );
   not U53983 ( n45732,p1_datawidth_reg_12_ );
   nand U53984 ( n52719,n45734,n45735 );
   not U53985 ( n45735,p1_datawidth_reg_15_ );
   not U53986 ( n45734,p1_datawidth_reg_14_ );
   nor U53987 ( n52717,n52721,n52722 );
   nand U53988 ( n52722,n45730,n45731 );
   not U53989 ( n45731,p1_datawidth_reg_11_ );
   not U53990 ( n45730,p1_datawidth_reg_10_ );
   and U53991 ( n52721,p1_datawidth_reg_0_,p1_datawidth_reg_1_ );
   nand U53992 ( n52715,n52723,n52724 );
   nor U53993 ( n52724,n52725,n52726 );
   nand U53994 ( n52726,n45740,n45741 );
   not U53995 ( n45741,p1_datawidth_reg_21_ );
   not U53996 ( n45740,p1_datawidth_reg_20_ );
   nand U53997 ( n52725,n45742,n45743 );
   not U53998 ( n45743,p1_datawidth_reg_23_ );
   not U53999 ( n45742,p1_datawidth_reg_22_ );
   nor U54000 ( n52723,n52727,n52728 );
   nand U54001 ( n52728,n45736,n45737 );
   not U54002 ( n45737,p1_datawidth_reg_17_ );
   not U54003 ( n45736,p1_datawidth_reg_16_ );
   nand U54004 ( n52727,n45738,n45739 );
   not U54005 ( n45739,p1_datawidth_reg_19_ );
   not U54006 ( n45738,p1_datawidth_reg_18_ );
   nand U54007 ( n52729,p1_flush_reg,n45365 );
   nand U54008 ( n45365,n45771,n45856 );
   nand U54009 ( n45856,n52730,n52731 );
   nand U54010 ( n52731,n45346,n52732 );
   nand U54011 ( n52732,n52733,n45351 );
   not U54012 ( n45351,n45360 );
   nor U54013 ( n45360,n51880,p1_state_reg_0_ );
   nand U54014 ( n51880,n45509,n52734 );
   nand U54015 ( n52734,p1_state_reg_2_,p1_state_reg_1_ );
   not U54016 ( n45509,n45513 );
   nor U54017 ( n52733,n51878,n45328 );
   nand U54018 ( n45346,ready11_reg,ready1 );
   nand U54019 ( n49020,n52735,n52736 );
   nor U54020 ( n52736,n45877,n52737 );
   nand U54021 ( n52737,n45869,n45432 );
   not U54022 ( n45877,n47303 );
   nor U54023 ( n52735,n52738,n52739 );
   nand U54024 ( n52739,n48249,n47446 );
   nor U54025 ( n48249,n48286,n45355 );
   not U54026 ( n48286,n49614 );
   nor U54027 ( n52740,n52742,n52743 );
   nor U54028 ( n52743,n47377,n28155 );
   not U54029 ( n45508,n45506 );
   not U54030 ( n47377,p1_statebs16_reg );
   nor U54031 ( n52742,n45506,n28898 );
   not U54032 ( n28898,bs16 );
   nand U54033 ( n52741,n45513,n45685 );
   not U54034 ( n45685,p1_state_reg_0_ );
   nor U54035 ( n45513,p1_state_reg_1_,p1_state_reg_2_ );
   nor U54036 ( n52744,n52745,n52746 );
   and U54037 ( n52746,n45332,p1_d_c_n_reg );
   nor U54038 ( n52745,p1_codefetch_reg,n45332 );
   not U54039 ( n45332,n45333 );
   nor U54040 ( n45333,n45686,p1_state_reg_0_ );
   nand U54041 ( n52748,p1_codefetch_reg,n52749 );
   nand U54042 ( n52749,n52730,n45771 );
   and U54043 ( n52730,n52750,n52751 );
   nand U54044 ( n52751,n52752,n52753 );
   or U54045 ( n52753,n45873,n45880 );
   not U54046 ( n45880,n45869 );
   nand U54047 ( n52752,n49630,n45876 );
   nor U54048 ( n52750,n48269,n52754 );
   nor U54049 ( n52754,n48279,n48169 );
   not U54050 ( n48169,n45328 );
   nor U54051 ( n45328,n47334,n47351 );
   not U54052 ( n48279,n45865 );
   nor U54053 ( n48269,n45869,n48289 );
   nand U54054 ( n52747,n45326,p1_state2_reg_0_ );
   nand U54055 ( n52755,p1_ads_n_reg,p1_state_reg_0_ );
   nor U54056 ( n45506,n52756,n45710 );
   nor U54057 ( n45710,p1_state_reg_0_,p1_state_reg_1_ );
   and U54058 ( n52756,n52757,p1_state_reg_0_ );
   nor U54059 ( n52757,p1_state_reg_2_,n45686 );
   not U54060 ( n45686,p1_state_reg_1_ );
   nand U54061 ( n52759,p1_memoryfetch_reg,n52760 );
   nand U54062 ( n52760,n52761,n52762 );
   nor U54063 ( n52762,n45865,n49624 );
   nand U54064 ( n45865,n52763,n52764 );
   nand U54065 ( n52764,n52765,n52766 );
   nor U54066 ( n52766,n52767,n52768 );
   nor U54067 ( n52765,n52769,n52770 );
   and U54068 ( n52761,n51664,n49630 );
   nor U54069 ( n49630,n48264,n47446 );
   not U54070 ( n47446,n45878 );
   or U54071 ( n48264,n45879,n47303 );
   nand U54072 ( n45879,n52771,n49614 );
   nor U54073 ( n49614,n48218,n47426 );
   not U54074 ( n47426,n47236 );
   not U54075 ( n48218,n47255 );
   nor U54076 ( n52771,n49602,n47287 );
   nor U54077 ( n52758,n52687,n45326 );
   and U54078 ( n45326,n45341,n45432 );
   not U54079 ( n45432,p1_state2_reg_1_ );
   nor U54080 ( n45341,p1_state2_reg_2_,p1_state2_reg_3_ );
   nor U54081 ( n52687,n48283,n45873 );
   nand U54082 ( n45873,n51876,n27892 );
   not U54083 ( n51876,n47433 );
   nand U54084 ( n47433,n52772,n52773 );
   nor U54085 ( n52773,n45878,n52774 );
   nand U54086 ( n52774,n47236,n47303 );
   nand U54087 ( n47303,n52775,n52776 );
   nor U54088 ( n52776,n52777,n52778 );
   nand U54089 ( n52778,n52779,n52780 );
   nor U54090 ( n52780,n52781,n52782 );
   nor U54091 ( n52782,n52783,n51923 );
   not U54092 ( n51923,p1_instqueue_reg_10__3_ );
   nor U54093 ( n52781,n52784,n51943 );
   not U54094 ( n51943,p1_instqueue_reg_8__3_ );
   nor U54095 ( n52779,n52785,n52786 );
   nor U54096 ( n52786,n52787,n51935 );
   not U54097 ( n51935,p1_instqueue_reg_15__3_ );
   nor U54098 ( n52785,n52788,n51934 );
   not U54099 ( n51934,p1_instqueue_reg_14__3_ );
   nand U54100 ( n52777,n52789,n52790 );
   nor U54101 ( n52790,n52791,n52792 );
   nor U54102 ( n52792,n52793,n47308 );
   not U54103 ( n47308,p1_instqueue_reg_0__3_ );
   nor U54104 ( n52791,n52794,n51912 );
   not U54105 ( n51912,p1_instqueue_reg_3__3_ );
   nor U54106 ( n52789,n52795,n52796 );
   nor U54107 ( n52796,n52797,n51944 );
   not U54108 ( n51944,p1_instqueue_reg_12__3_ );
   nor U54109 ( n52795,n52798,n51930 );
   not U54110 ( n51930,p1_instqueue_reg_11__3_ );
   nor U54111 ( n52775,n52799,n52800 );
   nand U54112 ( n52800,n52801,n52802 );
   nor U54113 ( n52802,n52803,n52804 );
   nor U54114 ( n52804,n52805,n51918 );
   not U54115 ( n51918,p1_instqueue_reg_6__3_ );
   nor U54116 ( n52803,n52806,n51913 );
   not U54117 ( n51913,p1_instqueue_reg_5__3_ );
   nor U54118 ( n52801,n52807,n52808 );
   nor U54119 ( n52808,n52809,n51940 );
   not U54120 ( n51940,p1_instqueue_reg_4__3_ );
   nor U54121 ( n52807,n52810,n51909 );
   not U54122 ( n51909,p1_instqueue_reg_2__3_ );
   nand U54123 ( n52799,n52811,n52812 );
   nor U54124 ( n52812,n52813,n52814 );
   nor U54125 ( n52814,n52815,n51922 );
   not U54126 ( n51922,p1_instqueue_reg_9__3_ );
   nor U54127 ( n52813,n52816,n51931 );
   not U54128 ( n51931,p1_instqueue_reg_13__3_ );
   nor U54129 ( n52811,n52817,n52818 );
   nor U54130 ( n52818,n52819,n51908 );
   not U54131 ( n51908,p1_instqueue_reg_1__3_ );
   nor U54132 ( n52817,n52179,n51919 );
   not U54133 ( n51919,p1_instqueue_reg_7__3_ );
   nand U54134 ( n47236,n52820,n52821 );
   nor U54135 ( n52821,n52822,n52823 );
   nand U54136 ( n52823,n52824,n52825 );
   nor U54137 ( n52825,n52826,n52827 );
   nor U54138 ( n52827,n52783,n51349 );
   not U54139 ( n51349,p1_instqueue_reg_10__7_ );
   nor U54140 ( n52826,n52784,n51355 );
   not U54141 ( n51355,p1_instqueue_reg_8__7_ );
   nor U54142 ( n52824,n52828,n52829 );
   nor U54143 ( n52829,n52787,n51337 );
   not U54144 ( n51337,p1_instqueue_reg_15__7_ );
   nor U54145 ( n52828,n52788,n51335 );
   not U54146 ( n51335,p1_instqueue_reg_14__7_ );
   nand U54147 ( n52822,n52830,n52831 );
   nor U54148 ( n52831,n52832,n52833 );
   nor U54149 ( n52833,n52793,n47243 );
   not U54150 ( n47243,p1_instqueue_reg_0__7_ );
   nor U54151 ( n52832,n52794,n51381 );
   not U54152 ( n51381,p1_instqueue_reg_3__7_ );
   nor U54153 ( n52830,n52834,n52835 );
   nor U54154 ( n52835,n52797,n51341 );
   not U54155 ( n51341,p1_instqueue_reg_12__7_ );
   nor U54156 ( n52834,n52798,n51351 );
   not U54157 ( n51351,p1_instqueue_reg_11__7_ );
   nor U54158 ( n52820,n52836,n52837 );
   nand U54159 ( n52837,n52838,n52839 );
   nor U54160 ( n52839,n52840,n52841 );
   nor U54161 ( n52841,n52805,n51365 );
   not U54162 ( n51365,p1_instqueue_reg_6__7_ );
   nor U54163 ( n52840,n52806,n51373 );
   not U54164 ( n51373,p1_instqueue_reg_5__7_ );
   nor U54165 ( n52838,n52842,n52843 );
   nor U54166 ( n52843,n52809,n51371 );
   not U54167 ( n51371,p1_instqueue_reg_4__7_ );
   nor U54168 ( n52842,n52810,n51379 );
   not U54169 ( n51379,p1_instqueue_reg_2__7_ );
   nand U54170 ( n52836,n52844,n52845 );
   nor U54171 ( n52845,n52846,n52847 );
   nor U54172 ( n52847,n52815,n51357 );
   not U54173 ( n51357,p1_instqueue_reg_9__7_ );
   nor U54174 ( n52846,n52816,n51343 );
   not U54175 ( n51343,p1_instqueue_reg_13__7_ );
   nor U54176 ( n52844,n52848,n52849 );
   nor U54177 ( n52849,n52819,n51386 );
   not U54178 ( n51386,p1_instqueue_reg_1__7_ );
   nor U54179 ( n52848,n52179,n51367 );
   not U54180 ( n51367,p1_instqueue_reg_7__7_ );
   nand U54181 ( n45878,n52850,n52851 );
   nor U54182 ( n52851,n52852,n52853 );
   nand U54183 ( n52853,n52854,n52855 );
   nor U54184 ( n52855,n52856,n52857 );
   nor U54185 ( n52857,n52783,n51510 );
   not U54186 ( n51510,p1_instqueue_reg_10__2_ );
   nor U54187 ( n52856,n52784,n51514 );
   not U54188 ( n51514,p1_instqueue_reg_8__2_ );
   nor U54189 ( n52854,n52858,n52859 );
   nor U54190 ( n52859,n52787,n51501 );
   not U54191 ( n51501,p1_instqueue_reg_15__2_ );
   nor U54192 ( n52858,n52788,n51500 );
   not U54193 ( n51500,p1_instqueue_reg_14__2_ );
   nand U54194 ( n52852,n52860,n52861 );
   nor U54195 ( n52861,n52862,n52863 );
   nor U54196 ( n52863,n52793,n47323 );
   not U54197 ( n47323,p1_instqueue_reg_0__2_ );
   nor U54198 ( n52862,n52794,n51533 );
   not U54199 ( n51533,p1_instqueue_reg_3__2_ );
   nor U54200 ( n52860,n52864,n52865 );
   nor U54201 ( n52865,n52797,n51504 );
   not U54202 ( n51504,p1_instqueue_reg_12__2_ );
   nor U54203 ( n52864,n52798,n51511 );
   not U54204 ( n51511,p1_instqueue_reg_11__2_ );
   nor U54205 ( n52850,n52866,n52867 );
   nand U54206 ( n52867,n52868,n52869 );
   nor U54207 ( n52869,n52870,n52871 );
   nor U54208 ( n52871,n52805,n51522 );
   not U54209 ( n51522,p1_instqueue_reg_6__2_ );
   nor U54210 ( n52870,n52806,n51527 );
   not U54211 ( n51527,p1_instqueue_reg_5__2_ );
   nor U54212 ( n52868,n52872,n52873 );
   nor U54213 ( n52873,n52809,n51526 );
   not U54214 ( n51526,p1_instqueue_reg_4__2_ );
   nor U54215 ( n52872,n52810,n51532 );
   not U54216 ( n51532,p1_instqueue_reg_2__2_ );
   nand U54217 ( n52866,n52874,n52875 );
   nor U54218 ( n52875,n52876,n52877 );
   nor U54219 ( n52877,n52815,n51515 );
   not U54220 ( n51515,p1_instqueue_reg_9__2_ );
   nor U54221 ( n52876,n52816,n51505 );
   not U54222 ( n51505,p1_instqueue_reg_13__2_ );
   nor U54223 ( n52874,n52878,n52879 );
   nor U54224 ( n52879,n52819,n51536 );
   not U54225 ( n51536,p1_instqueue_reg_1__2_ );
   nor U54226 ( n52878,n52179,n51523 );
   not U54227 ( n51523,p1_instqueue_reg_7__2_ );
   nor U54228 ( n52772,n47255,n52880 );
   nand U54229 ( n52880,n49602,n48247 );
   nand U54230 ( n47255,n52881,n52882 );
   nor U54231 ( n52882,n52883,n52884 );
   nand U54232 ( n52884,n52885,n52886 );
   nor U54233 ( n52886,n52887,n52888 );
   nor U54234 ( n52888,n52783,n51409 );
   not U54235 ( n51409,p1_instqueue_reg_10__6_ );
   nor U54236 ( n52887,n52784,n51413 );
   not U54237 ( n51413,p1_instqueue_reg_8__6_ );
   nor U54238 ( n52885,n52889,n52890 );
   nor U54239 ( n52890,n52787,n51400 );
   not U54240 ( n51400,p1_instqueue_reg_15__6_ );
   nor U54241 ( n52889,n52788,n51399 );
   not U54242 ( n51399,p1_instqueue_reg_14__6_ );
   nand U54243 ( n52883,n52891,n52892 );
   nor U54244 ( n52892,n52893,n52894 );
   nor U54245 ( n52894,n52793,n47260 );
   not U54246 ( n47260,p1_instqueue_reg_0__6_ );
   nor U54247 ( n52893,n52895,n51432 );
   not U54248 ( n51432,p1_instqueue_reg_3__6_ );
   nor U54249 ( n52891,n52896,n52897 );
   nor U54250 ( n52897,n52797,n51403 );
   not U54251 ( n51403,p1_instqueue_reg_12__6_ );
   nor U54252 ( n52896,n52798,n51410 );
   not U54253 ( n51410,p1_instqueue_reg_11__6_ );
   nor U54254 ( n52881,n52898,n52899 );
   nand U54255 ( n52899,n52900,n52901 );
   nor U54256 ( n52901,n52902,n52903 );
   nor U54257 ( n52903,n52805,n51421 );
   not U54258 ( n51421,p1_instqueue_reg_6__6_ );
   nor U54259 ( n52902,n52806,n51426 );
   not U54260 ( n51426,p1_instqueue_reg_5__6_ );
   nor U54261 ( n52900,n52904,n52905 );
   nor U54262 ( n52905,n52809,n51425 );
   not U54263 ( n51425,p1_instqueue_reg_4__6_ );
   nor U54264 ( n52904,n52810,n51431 );
   not U54265 ( n51431,p1_instqueue_reg_2__6_ );
   nand U54266 ( n52898,n52906,n52907 );
   nor U54267 ( n52907,n52908,n52909 );
   nor U54268 ( n52909,n52815,n51414 );
   not U54269 ( n51414,p1_instqueue_reg_9__6_ );
   nor U54270 ( n52908,n52816,n51404 );
   not U54271 ( n51404,p1_instqueue_reg_13__6_ );
   nor U54272 ( n52906,n52910,n52911 );
   nor U54273 ( n52911,n52819,n51435 );
   not U54274 ( n51435,p1_instqueue_reg_1__6_ );
   nor U54275 ( n52910,n52179,n51422 );
   not U54276 ( n51422,p1_instqueue_reg_7__6_ );
   nand U54277 ( n48283,n45771,n45869 );
   nand U54278 ( n45869,n52912,n52913 );
   nand U54279 ( n52913,n52914,n52915 );
   nand U54280 ( n52915,n52916,n52917 );
   nand U54281 ( n52917,n52918,n52919 );
   nand U54282 ( n52918,n52920,n52921 );
   nand U54283 ( n52921,n52768,n48270 );
   nand U54284 ( n52920,n52922,n52767 );
   nand U54285 ( n52916,n52923,n52924 );
   nand U54286 ( n52924,n52925,n52926 );
   nor U54287 ( n52923,n52927,n52928 );
   nor U54288 ( n52928,n52929,n52930 );
   nor U54289 ( n52930,n52931,n52932 );
   and U54290 ( n52932,n52933,n52934 );
   nor U54291 ( n52931,n52935,n52936 );
   nor U54292 ( n52936,n52934,n52933 );
   nand U54293 ( n52933,n52937,n52938 );
   nand U54294 ( n52938,n52939,n48870 );
   nor U54295 ( n48870,n48289,n49602 );
   nor U54296 ( n52939,n52940,n48270 );
   nand U54297 ( n52937,n52941,n52942 );
   nor U54298 ( n52941,n52940,n52943 );
   nor U54299 ( n52943,n52944,n52945 );
   and U54300 ( n52940,n52946,n52738 );
   nand U54301 ( n52738,n52947,n52948 );
   nor U54302 ( n52947,n49602,n45876 );
   and U54303 ( n52946,n52945,n52949 );
   and U54304 ( n52945,n52950,n52951 );
   nand U54305 ( n52951,p1_instqueuewr_addr_reg_0_,n45451 );
   nand U54306 ( n52934,n52952,n52953 );
   nor U54307 ( n52953,n49602,n45350 );
   nor U54308 ( n52952,n52954,n52955 );
   nor U54309 ( n52955,n48289,n52057 );
   nor U54310 ( n52954,n52956,n48270 );
   nor U54311 ( n52935,n52944,n52956 );
   not U54312 ( n52956,n52770 );
   xor U54313 ( n52770,n52957,n52958 );
   xor U54314 ( n52957,n45842,n45825 );
   nor U54315 ( n52929,n52925,n52926 );
   nand U54316 ( n52926,n52949,n52959 );
   nand U54317 ( n52959,n52769,n51730 );
   nand U54318 ( n52949,n48289,n52960 );
   or U54319 ( n52960,n47271,n49622 );
   not U54320 ( n47271,n49602 );
   and U54321 ( n52925,n52942,n52961 );
   nand U54322 ( n52961,n52769,n52919 );
   xor U54323 ( n52769,n52962,n52963 );
   xor U54324 ( n52962,n45840,n47402 );
   nand U54325 ( n52942,n51733,n52057 );
   nor U54326 ( n52927,n48270,n52964 );
   nand U54327 ( n52964,n52768,n52944 );
   xor U54328 ( n52768,n52965,n52966 );
   xor U54329 ( n52965,n46275,n50913 );
   nor U54330 ( n52914,n52967,n52968 );
   nor U54331 ( n52968,n52944,n52969 );
   nand U54332 ( n52969,n52970,n48270 );
   not U54333 ( n52944,n52919 );
   nor U54334 ( n52967,n52922,n52919 );
   and U54335 ( n52922,n52971,n52972 );
   nand U54336 ( n52972,n51730,n52767 );
   xor U54337 ( n52767,n52973,n52974 );
   xor U54338 ( n52973,p1_instqueuewr_addr_reg_4_,p1_instqueuerd_addr_reg_4_ );
   not U54339 ( n51730,n48270 );
   nand U54340 ( n52971,p1_instqueuerd_addr_reg_4_,n28095 );
   nand U54341 ( n52912,n52975,n52970 );
   not U54342 ( n52970,n52763 );
   nand U54343 ( n52763,n52976,n52977 );
   nand U54344 ( n52977,p1_instqueuewr_addr_reg_4_,n52978 );
   nand U54345 ( n52978,p1_instqueuerd_addr_reg_4_,n52974 );
   or U54346 ( n52976,n52974,p1_instqueuerd_addr_reg_4_ );
   nand U54347 ( n52974,n52979,n52980 );
   nand U54348 ( n52980,n52981,n46275 );
   not U54349 ( n46275,p1_instqueuewr_addr_reg_3_ );
   or U54350 ( n52981,n52966,p1_instqueuerd_addr_reg_3_ );
   nand U54351 ( n52979,p1_instqueuerd_addr_reg_3_,n52966 );
   nand U54352 ( n52966,n52982,n52983 );
   nand U54353 ( n52983,n52984,n45840 );
   not U54354 ( n45840,p1_instqueuewr_addr_reg_2_ );
   or U54355 ( n52984,n52963,p1_instqueuerd_addr_reg_2_ );
   nand U54356 ( n52982,p1_instqueuerd_addr_reg_2_,n52963 );
   nand U54357 ( n52963,n52985,n52986 );
   nand U54358 ( n52986,n52987,n45842 );
   not U54359 ( n45842,p1_instqueuewr_addr_reg_1_ );
   nand U54360 ( n52987,n45825,n52950 );
   not U54361 ( n52950,n52958 );
   nand U54362 ( n52985,n52958,p1_instqueuerd_addr_reg_1_ );
   nor U54363 ( n52958,n45451,p1_instqueuewr_addr_reg_0_ );
   nor U54364 ( n52975,n52919,n48270 );
   nand U54365 ( n48270,n52988,p1_state2_reg_0_ );
   nor U54366 ( n52988,n48247,n45876 );
   not U54367 ( n48247,n47287 );
   nand U54368 ( n52919,n52989,n52990 );
   nor U54369 ( n52990,n45350,n49622 );
   nor U54370 ( n49622,n47334,n51733 );
   nor U54371 ( n45350,n51733,n48289 );
   not U54372 ( n51733,n51664 );
   nor U54373 ( n51664,n47351,n45347 );
   nor U54374 ( n52989,n52991,n52992 );
   nor U54375 ( n52992,n49620,n52057 );
   not U54376 ( n52057,n52948 );
   nor U54377 ( n52948,n47287,n28095 );
   nand U54378 ( n47287,n52993,n52994 );
   nor U54379 ( n52994,n52995,n52996 );
   nand U54380 ( n52996,n52997,n52998 );
   nor U54381 ( n52998,n52999,n53000 );
   nor U54382 ( n53000,n52783,n51971 );
   not U54383 ( n51971,p1_instqueue_reg_10__4_ );
   nor U54384 ( n52999,n52784,n51991 );
   not U54385 ( n51991,p1_instqueue_reg_8__4_ );
   nor U54386 ( n52997,n53001,n53002 );
   nor U54387 ( n53002,n52787,n51983 );
   not U54388 ( n51983,p1_instqueue_reg_15__4_ );
   nor U54389 ( n53001,n52788,n51982 );
   not U54390 ( n51982,p1_instqueue_reg_14__4_ );
   nand U54391 ( n52995,n53003,n53004 );
   nor U54392 ( n53004,n53005,n53006 );
   nor U54393 ( n53006,n52793,n47292 );
   not U54394 ( n47292,p1_instqueue_reg_0__4_ );
   nor U54395 ( n53005,n52895,n51960 );
   not U54396 ( n51960,p1_instqueue_reg_3__4_ );
   nor U54397 ( n53003,n53007,n53008 );
   nor U54398 ( n53008,n52797,n51992 );
   not U54399 ( n51992,p1_instqueue_reg_12__4_ );
   nor U54400 ( n53007,n52798,n51978 );
   not U54401 ( n51978,p1_instqueue_reg_11__4_ );
   nor U54402 ( n52993,n53009,n53010 );
   nand U54403 ( n53010,n53011,n53012 );
   nor U54404 ( n53012,n53013,n53014 );
   nor U54405 ( n53014,n52805,n51966 );
   not U54406 ( n51966,p1_instqueue_reg_6__4_ );
   nor U54407 ( n53013,n52806,n51961 );
   not U54408 ( n51961,p1_instqueue_reg_5__4_ );
   nor U54409 ( n53011,n53015,n53016 );
   nor U54410 ( n53016,n52809,n51988 );
   not U54411 ( n51988,p1_instqueue_reg_4__4_ );
   nor U54412 ( n53015,n52810,n51957 );
   not U54413 ( n51957,p1_instqueue_reg_2__4_ );
   nand U54414 ( n53009,n53017,n53018 );
   nor U54415 ( n53018,n53019,n53020 );
   nor U54416 ( n53020,n52815,n51970 );
   not U54417 ( n51970,p1_instqueue_reg_9__4_ );
   nor U54418 ( n53019,n52816,n51979 );
   not U54419 ( n51979,p1_instqueue_reg_13__4_ );
   nor U54420 ( n53017,n53021,n53022 );
   nor U54421 ( n53022,n52819,n51956 );
   not U54422 ( n51956,p1_instqueue_reg_1__4_ );
   nor U54423 ( n53021,n52179,n51967 );
   not U54424 ( n51967,p1_instqueue_reg_7__4_ );
   not U54425 ( n49620,n51878 );
   nor U54426 ( n51878,n48289,n45876 );
   not U54427 ( n48289,n47334 );
   nor U54428 ( n52991,n53023,n45347 );
   nor U54429 ( n53023,n49602,n45358 );
   nor U54430 ( n45358,n47334,n45876 );
   not U54431 ( n45876,n47351 );
   nand U54432 ( n47351,n53024,n53025 );
   nor U54433 ( n53025,n53026,n53027 );
   nand U54434 ( n53027,n53028,n53029 );
   nor U54435 ( n53029,n53030,n53031 );
   nor U54436 ( n53031,n52783,n51610 );
   not U54437 ( n51610,p1_instqueue_reg_10__0_ );
   nor U54438 ( n53030,n52784,n51614 );
   not U54439 ( n51614,p1_instqueue_reg_8__0_ );
   nor U54440 ( n53028,n53032,n53033 );
   nor U54441 ( n53033,n52787,n51601 );
   not U54442 ( n51601,p1_instqueue_reg_15__0_ );
   nor U54443 ( n53032,n52788,n51600 );
   not U54444 ( n51600,p1_instqueue_reg_14__0_ );
   nand U54445 ( n53026,n53034,n53035 );
   nor U54446 ( n53035,n53036,n53037 );
   nor U54447 ( n53037,n52793,n47364 );
   not U54448 ( n47364,p1_instqueue_reg_0__0_ );
   nor U54449 ( n53036,n52794,n51633 );
   not U54450 ( n51633,p1_instqueue_reg_3__0_ );
   nor U54451 ( n53034,n53038,n53039 );
   nor U54452 ( n53039,n52797,n51604 );
   not U54453 ( n51604,p1_instqueue_reg_12__0_ );
   nor U54454 ( n53038,n52798,n51611 );
   not U54455 ( n51611,p1_instqueue_reg_11__0_ );
   nor U54456 ( n53024,n53040,n53041 );
   nand U54457 ( n53041,n53042,n53043 );
   nor U54458 ( n53043,n53044,n53045 );
   nor U54459 ( n53045,n52805,n51622 );
   not U54460 ( n51622,p1_instqueue_reg_6__0_ );
   nor U54461 ( n53044,n52806,n51627 );
   not U54462 ( n51627,p1_instqueue_reg_5__0_ );
   nor U54463 ( n53042,n53046,n53047 );
   nor U54464 ( n53047,n52809,n51626 );
   not U54465 ( n51626,p1_instqueue_reg_4__0_ );
   nor U54466 ( n53046,n52810,n51632 );
   not U54467 ( n51632,p1_instqueue_reg_2__0_ );
   nand U54468 ( n53040,n53048,n53049 );
   nor U54469 ( n53049,n53050,n53051 );
   nor U54470 ( n53051,n52815,n51615 );
   not U54471 ( n51615,p1_instqueue_reg_9__0_ );
   nor U54472 ( n53050,n52816,n51605 );
   not U54473 ( n51605,p1_instqueue_reg_13__0_ );
   nor U54474 ( n53048,n53052,n53053 );
   nor U54475 ( n53053,n52819,n51636 );
   not U54476 ( n51636,p1_instqueue_reg_1__0_ );
   nor U54477 ( n53052,n52179,n51623 );
   not U54478 ( n51623,p1_instqueue_reg_7__0_ );
   nand U54479 ( n47334,n53054,n53055 );
   nor U54480 ( n53055,n53056,n53057 );
   nand U54481 ( n53057,n53058,n53059 );
   nor U54482 ( n53059,n53060,n53061 );
   nor U54483 ( n53061,n52783,n51560 );
   not U54484 ( n51560,p1_instqueue_reg_10__1_ );
   nor U54485 ( n53060,n52784,n51564 );
   not U54486 ( n51564,p1_instqueue_reg_8__1_ );
   nor U54487 ( n53058,n53062,n53063 );
   nor U54488 ( n53063,n52787,n51551 );
   not U54489 ( n51551,p1_instqueue_reg_15__1_ );
   nor U54490 ( n53062,n52788,n51550 );
   not U54491 ( n51550,p1_instqueue_reg_14__1_ );
   nand U54492 ( n53056,n53064,n53065 );
   nor U54493 ( n53065,n53066,n53067 );
   nor U54494 ( n53067,n52793,n47339 );
   not U54495 ( n47339,p1_instqueue_reg_0__1_ );
   nor U54496 ( n53066,n52794,n51583 );
   not U54497 ( n51583,p1_instqueue_reg_3__1_ );
   nand U54498 ( n52794,n47403,n47399 );
   nor U54499 ( n53064,n53068,n53069 );
   nor U54500 ( n53069,n52797,n51554 );
   not U54501 ( n51554,p1_instqueue_reg_12__1_ );
   nor U54502 ( n53068,n52798,n51561 );
   not U54503 ( n51561,p1_instqueue_reg_11__1_ );
   nor U54504 ( n53054,n53070,n53071 );
   nand U54505 ( n53071,n53072,n53073 );
   nor U54506 ( n53073,n53074,n53075 );
   nor U54507 ( n53075,n52805,n51572 );
   not U54508 ( n51572,p1_instqueue_reg_6__1_ );
   nor U54509 ( n53074,n52806,n51577 );
   not U54510 ( n51577,p1_instqueue_reg_5__1_ );
   nor U54511 ( n53072,n53076,n53077 );
   nor U54512 ( n53077,n52809,n51576 );
   not U54513 ( n51576,p1_instqueue_reg_4__1_ );
   nor U54514 ( n53076,n52810,n51582 );
   not U54515 ( n51582,p1_instqueue_reg_2__1_ );
   nand U54516 ( n53070,n53078,n53079 );
   nor U54517 ( n53079,n53080,n53081 );
   nor U54518 ( n53081,n52815,n51565 );
   not U54519 ( n51565,p1_instqueue_reg_9__1_ );
   nor U54520 ( n53080,n52816,n51555 );
   not U54521 ( n51555,p1_instqueue_reg_13__1_ );
   nor U54522 ( n53078,n53082,n53083 );
   nor U54523 ( n53083,n52819,n51586 );
   not U54524 ( n51586,p1_instqueue_reg_1__1_ );
   nor U54525 ( n53082,n52179,n51573 );
   not U54526 ( n51573,p1_instqueue_reg_7__1_ );
   nor U54527 ( n49602,n51895,n53084 );
   nor U54528 ( n53084,n47276,n52793 );
   nand U54529 ( n52793,n52442,n50913 );
   not U54530 ( n47276,p1_instqueue_reg_0__5_ );
   nand U54531 ( n51895,n53085,n53086 );
   nor U54532 ( n53086,n53087,n53088 );
   nand U54533 ( n53088,n53089,n53090 );
   nor U54534 ( n53090,n53091,n53092 );
   nor U54535 ( n53092,n52788,n51449 );
   not U54536 ( n51449,p1_instqueue_reg_14__5_ );
   nand U54537 ( n52788,n52457,p1_instqueuerd_addr_reg_3_ );
   nor U54538 ( n52457,n52448,n47402 );
   not U54539 ( n52448,n52110 );
   nor U54540 ( n53091,n52783,n51459 );
   not U54541 ( n51459,p1_instqueue_reg_10__5_ );
   nand U54542 ( n52783,n52110,n52474 );
   nor U54543 ( n53089,n53093,n53094 );
   nor U54544 ( n53094,n52816,n51454 );
   not U54545 ( n51454,p1_instqueue_reg_13__5_ );
   nand U54546 ( n52816,n52454,p1_instqueuerd_addr_reg_3_ );
   nor U54547 ( n52454,n52444,n47402 );
   not U54548 ( n52444,n52107 );
   nor U54549 ( n53093,n52787,n51450 );
   not U54550 ( n51450,p1_instqueue_reg_15__5_ );
   nand U54551 ( n52787,n52181,p1_instqueuerd_addr_reg_3_ );
   nor U54552 ( n52181,n47402,n53095 );
   nand U54553 ( n53087,n53096,n53097 );
   nor U54554 ( n53097,n53098,n53099 );
   nor U54555 ( n53099,n52798,n51460 );
   not U54556 ( n51460,p1_instqueue_reg_11__5_ );
   nand U54557 ( n52798,p1_instqueuerd_addr_reg_3_,n52183 );
   nor U54558 ( n53098,n52895,n51482 );
   not U54559 ( n51482,p1_instqueue_reg_3__5_ );
   nand U54560 ( n52895,n52183,n50913 );
   nor U54561 ( n52183,n53095,p1_instqueuerd_addr_reg_2_ );
   not U54562 ( n53095,n47399 );
   nor U54563 ( n53096,n53100,n53101 );
   nor U54564 ( n53101,n52784,n51463 );
   not U54565 ( n51463,p1_instqueue_reg_8__5_ );
   nand U54566 ( n52784,p1_instqueuerd_addr_reg_3_,n52442 );
   nor U54567 ( n52442,n47407,p1_instqueuerd_addr_reg_2_ );
   nor U54568 ( n53100,n52797,n51453 );
   not U54569 ( n51453,p1_instqueue_reg_12__5_ );
   nand U54570 ( n52797,n52453,p1_instqueuerd_addr_reg_3_ );
   nor U54571 ( n52453,n47402,n47407 );
   not U54572 ( n47407,n52106 );
   nor U54573 ( n53085,n53102,n53103 );
   nand U54574 ( n53103,n53104,n53105 );
   or U54575 ( n53105,n51475,n52809 );
   nand U54576 ( n52809,n52139,n52106 );
   nor U54577 ( n52106,p1_instqueuerd_addr_reg_0_,p1_instqueuerd_addr_reg_1_ );
   not U54578 ( n51475,p1_instqueue_reg_4__5_ );
   nor U54579 ( n53104,n53106,n53107 );
   nor U54580 ( n53107,n52810,n51481 );
   not U54581 ( n51481,p1_instqueue_reg_2__5_ );
   nand U54582 ( n52810,n52110,n47403 );
   nor U54583 ( n53106,n52805,n51471 );
   not U54584 ( n51471,p1_instqueue_reg_6__5_ );
   nand U54585 ( n52805,n52139,n52110 );
   nor U54586 ( n52110,n45825,p1_instqueuerd_addr_reg_0_ );
   nand U54587 ( n53102,n53108,n53109 );
   nor U54588 ( n53109,n53110,n53111 );
   nor U54589 ( n53111,n52179,n51472 );
   not U54590 ( n51472,p1_instqueue_reg_7__5_ );
   nand U54591 ( n52179,n52139,n47399 );
   nor U54592 ( n47399,n45825,n45451 );
   not U54593 ( n45825,p1_instqueuerd_addr_reg_1_ );
   nor U54594 ( n53110,n52815,n51464 );
   not U54595 ( n51464,p1_instqueue_reg_9__5_ );
   nand U54596 ( n52815,n52107,n52474 );
   nor U54597 ( n52474,n50913,p1_instqueuerd_addr_reg_2_ );
   not U54598 ( n50913,p1_instqueuerd_addr_reg_3_ );
   nor U54599 ( n53108,n53112,n53113 );
   nor U54600 ( n53113,n52806,n51476 );
   not U54601 ( n51476,p1_instqueue_reg_5__5_ );
   nand U54602 ( n52806,n52139,n52107 );
   nor U54603 ( n52139,n47402,p1_instqueuerd_addr_reg_3_ );
   not U54604 ( n47402,p1_instqueuerd_addr_reg_2_ );
   nor U54605 ( n53112,n52819,n51485 );
   not U54606 ( n51485,p1_instqueue_reg_1__5_ );
   nand U54607 ( n52819,n52107,n47403 );
   nor U54608 ( n47403,p1_instqueuerd_addr_reg_2_,p1_instqueuerd_addr_reg_3_ );
   nor U54609 ( n52107,n45451,p1_instqueuerd_addr_reg_1_ );
   not U54610 ( n45451,p1_instqueuerd_addr_reg_0_ );
   nor U54611 ( n45771,n28094,n49624 );
   not U54612 ( n49624,n45759 );
   nor U54613 ( n45759,n28374,p1_state2_reg_1_ );
   not U54614 ( n45355,p1_state2_reg_2_ );
   not U54615 ( n45347,p1_state2_reg_0_ );
endmodule
