
module b12 ( start, k_3_, k_2_, k_1_, k_0_, count_reg_0_, memory_reg_31__1_,
memory_reg_31__0_, memory_reg_30__1_, memory_reg_30__0_,
memory_reg_29__1_, memory_reg_29__0_, memory_reg_28__1_,
memory_reg_28__0_, memory_reg_27__1_, memory_reg_27__0_,
memory_reg_26__1_, memory_reg_26__0_, memory_reg_25__1_,
memory_reg_25__0_, memory_reg_24__1_, memory_reg_24__0_,
memory_reg_23__1_, memory_reg_23__0_, memory_reg_22__1_,
memory_reg_22__0_, memory_reg_21__1_, memory_reg_21__0_,
memory_reg_20__1_, memory_reg_20__0_, memory_reg_19__1_,
memory_reg_19__0_, memory_reg_18__1_, memory_reg_18__0_,
memory_reg_17__1_, memory_reg_17__0_, memory_reg_16__1_,
memory_reg_16__0_, memory_reg_15__1_, memory_reg_15__0_,
memory_reg_14__1_, memory_reg_14__0_, memory_reg_13__1_,
memory_reg_13__0_, memory_reg_12__1_, memory_reg_12__0_,
memory_reg_11__1_, memory_reg_11__0_, memory_reg_10__1_,
memory_reg_10__0_, memory_reg_9__1_, memory_reg_9__0_,
memory_reg_8__1_, memory_reg_8__0_, memory_reg_7__1_, memory_reg_7__0_,
memory_reg_6__1_, memory_reg_6__0_, memory_reg_5__1_, memory_reg_5__0_,
memory_reg_4__1_, memory_reg_4__0_, memory_reg_3__1_, memory_reg_3__0_,
memory_reg_2__1_, memory_reg_2__0_, memory_reg_1__1_, memory_reg_1__0_,
memory_reg_0__1_, memory_reg_0__0_, nl_reg_3_, nl_reg_2_, nl_reg_1_,
nl_reg_0_, scan_reg_4_, scan_reg_3_, scan_reg_2_, scan_reg_1_,
scan_reg_0_, max_reg_4_, max_reg_3_, max_reg_2_, max_reg_1_,
max_reg_0_, ind_reg_1_, ind_reg_0_, timebase_reg_5_, timebase_reg_4_,
timebase_reg_3_, timebase_reg_2_, timebase_reg_1_, timebase_reg_0_,
count_reg2_5_, count_reg2_4_, count_reg2_3_, count_reg2_2_,
count_reg2_1_, count_reg2_0_, sound_reg_2_, sound_reg_1_, sound_reg_0_,
address_reg_4_, address_reg_3_, address_reg_2_, address_reg_1_,
address_reg_0_, data_in_reg_1_, data_in_reg_0_, s_reg, play_reg,
nloss_reg, speaker_reg, wr_reg, counter_reg_2_, counter_reg_1_,
counter_reg_0_, count_reg_1_, num_reg_1_, num_reg_0_, data_out_reg_1_,
data_out_reg_0_, gamma_reg_4_, gamma_reg_3_, gamma_reg_2_,
gamma_reg_1_, gamma_reg_0_, u1391, u1486, u1485, u1484, u1483, u1482,
u1481, u1480, u1479, u1478, u1477, u1476, u1475, u1474, u1473, u1472,
u1471, u1470, u1469, u1468, u1467, u1466, u1465, u1464, u1463, u1462,
u1461, u1460, u1459, u1458, u1457, u1456, u1455, u1454, u1453, u1452,
u1451, u1450, u1449, u1448, u1447, u1446, u1445, u1444, u1443, u1442,
u1441, u1440, u1439, u1438, u1437, u1436, u1435, u1434, u1433, u1432,
u1431, u1430, u1429, u1428, u1427, u1426, u1425, u1424, u1423, u1422,
u1421, u1420, u1419, u1418, u1417, u1416, u1415, u1414, u1413, u1412,
u1411, u1410, u1409, u1564, u1565, u1566, u1408, u1407, u1406, u1405,
u1567, u1404, u1403, u1568, u1402, u1401, u1400, u1569, u1570, u1571,
u1399, u1398, u1397, u1396, u1395, u1572, u1573, u1394, u1574, u1575,
u1393, u1392, u1381, u1382, u1383, u1563, u1390, u1389, u1384, u1385,
u1386, u1387, u1388 );
input start, k_3_, k_2_, k_1_, k_0_, count_reg_0_, memory_reg_31__1_,
memory_reg_31__0_, memory_reg_30__1_, memory_reg_30__0_,
memory_reg_29__1_, memory_reg_29__0_, memory_reg_28__1_,
memory_reg_28__0_, memory_reg_27__1_, memory_reg_27__0_,
memory_reg_26__1_, memory_reg_26__0_, memory_reg_25__1_,
memory_reg_25__0_, memory_reg_24__1_, memory_reg_24__0_,
memory_reg_23__1_, memory_reg_23__0_, memory_reg_22__1_,
memory_reg_22__0_, memory_reg_21__1_, memory_reg_21__0_,
memory_reg_20__1_, memory_reg_20__0_, memory_reg_19__1_,
memory_reg_19__0_, memory_reg_18__1_, memory_reg_18__0_,
memory_reg_17__1_, memory_reg_17__0_, memory_reg_16__1_,
memory_reg_16__0_, memory_reg_15__1_, memory_reg_15__0_,
memory_reg_14__1_, memory_reg_14__0_, memory_reg_13__1_,
memory_reg_13__0_, memory_reg_12__1_, memory_reg_12__0_,
memory_reg_11__1_, memory_reg_11__0_, memory_reg_10__1_,
memory_reg_10__0_, memory_reg_9__1_, memory_reg_9__0_,
memory_reg_8__1_, memory_reg_8__0_, memory_reg_7__1_,
memory_reg_7__0_, memory_reg_6__1_, memory_reg_6__0_,
memory_reg_5__1_, memory_reg_5__0_, memory_reg_4__1_,
memory_reg_4__0_, memory_reg_3__1_, memory_reg_3__0_,
memory_reg_2__1_, memory_reg_2__0_, memory_reg_1__1_,
memory_reg_1__0_, memory_reg_0__1_, memory_reg_0__0_, nl_reg_3_,
nl_reg_2_, nl_reg_1_, nl_reg_0_, scan_reg_4_, scan_reg_3_,
scan_reg_2_, scan_reg_1_, scan_reg_0_, max_reg_4_, max_reg_3_,
max_reg_2_, max_reg_1_, max_reg_0_, ind_reg_1_, ind_reg_0_,
timebase_reg_5_, timebase_reg_4_, timebase_reg_3_, timebase_reg_2_,
timebase_reg_1_, timebase_reg_0_, count_reg2_5_, count_reg2_4_,
count_reg2_3_, count_reg2_2_, count_reg2_1_, count_reg2_0_,
sound_reg_2_, sound_reg_1_, sound_reg_0_, address_reg_4_,
address_reg_3_, address_reg_2_, address_reg_1_, address_reg_0_,
data_in_reg_1_, data_in_reg_0_, s_reg, play_reg, nloss_reg,
speaker_reg, wr_reg, counter_reg_2_, counter_reg_1_, counter_reg_0_,
count_reg_1_, num_reg_1_, num_reg_0_, data_out_reg_1_,
data_out_reg_0_, gamma_reg_4_, gamma_reg_3_, gamma_reg_2_,
gamma_reg_1_, gamma_reg_0_;
output u1391, u1486, u1485, u1484, u1483, u1482, u1481, u1480, u1479, u1478,
u1477, u1476, u1475, u1474, u1473, u1472, u1471, u1470, u1469, u1468,
u1467, u1466, u1465, u1464, u1463, u1462, u1461, u1460, u1459, u1458,
u1457, u1456, u1455, u1454, u1453, u1452, u1451, u1450, u1449, u1448,
u1447, u1446, u1445, u1444, u1443, u1442, u1441, u1440, u1439, u1438,
u1437, u1436, u1435, u1434, u1433, u1432, u1431, u1430, u1429, u1428,
u1427, u1426, u1425, u1424, u1423, u1422, u1421, u1420, u1419, u1418,
u1417, u1416, u1415, u1414, u1413, u1412, u1411, u1410, u1409, u1564,
u1565, u1566, u1408, u1407, u1406, u1405, u1567, u1404, u1403, u1568,
u1402, u1401, u1400, u1569, u1570, u1571, u1399, u1398, u1397, u1396,
u1395, u1572, u1573, u1394, u1574, u1575, u1393, u1392, u1381, u1382,
u1383, u1563, u1390, u1389, u1384, u1385, u1386, u1387, u1388;
wire   n2947, n2948, n2949, n1460, n1462, n1465, n1466, n1467, n1468, n1469,
n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
n2940, n2941, n2942, n2943, n2944, n2945, n2946;

   not U1579 ( n1460,n2947 );
   not U1580 ( u1381,n1460 );
   not U1581 ( n1462,n2949 );
   not U1582 ( u1563,n1462 );
   not U1583 ( u1383,n2919 );
   not U1584 ( n1465,n1973 );
   not U1585 ( n1468,n1973 );
   not U1586 ( n1466,n1973 );
   not U1587 ( n1467,n1973 );
   not U1588 ( n1469,n1979 );
   not U1589 ( n1472,n1979 );
   not U1590 ( n1470,n1979 );
   not U1591 ( n1471,n1979 );
   not U1592 ( n1473,wr_reg );
   not U1593 ( n1476,wr_reg );
   not U1594 ( n1474,wr_reg );
   not U1595 ( n1475,wr_reg );
   buf U1596 ( n1477,n1513 );
   not U1597 ( n1478,n2294 );
   not U1598 ( u1575,n1479 );
   nor U1599 ( n1479,n1480,n1481 );
   nor U1600 ( n1481,n1482,n1483 );
   not U1601 ( n1483,nloss_reg );
   not U1602 ( n1482,n1484 );
   nor U1603 ( n1480,n1484,n1485 );
   nor U1604 ( n1484,n1486,n1487 );
   not U1605 ( n1487,n1488 );
   nor U1606 ( n1488,n1489,n1490 );
   not U1607 ( u1574,n1491 );
   nor U1608 ( n1491,n1492,n1493 );
   nor U1609 ( n1493,n1494,n1495 );
   nor U1610 ( n1495,n1496,n1497 );
   not U1611 ( n1497,n1498 );
   nor U1612 ( n1498,n1499,n1500 );
   nor U1613 ( n1500,n1501,n1502 );
   not U1614 ( n1502,n1503 );
   nor U1615 ( n1503,n1504,n1505 );
   nor U1616 ( n1505,n1506,n1507 );
   nor U1617 ( n1499,n1508,n1509 );
   nor U1618 ( n1509,n1510,n1511 );
   nor U1619 ( n1510,n1512,n1477 );
   nor U1620 ( n1496,n1514,n1515 );
   nor U1621 ( n1492,n1516,n1517 );
   not U1622 ( n1517,n1494 );
   nor U1623 ( n1494,n1518,n1519 );
   not U1624 ( n1519,n1520 );
   nor U1625 ( n1520,n1521,n1522 );
   nor U1626 ( n1521,n1523,n1478 );
   nor U1627 ( n1523,n1525,n1526 );
   not U1628 ( n1526,n1527 );
   nor U1629 ( n1527,n1528,n1529 );
   nor U1630 ( n1525,n1513,n1530 );
   not U1631 ( n1530,n1531 );
   nor U1632 ( n1531,n1508,n1532 );
   not U1633 ( n1518,n1533 );
   nor U1634 ( n1533,n1534,n1535 );
   not U1635 ( n1535,n1536 );
   nor U1636 ( n1536,n1537,n1538 );
   not U1637 ( u1573,n1539 );
   nor U1638 ( n1539,n1540,n1541 );
   nor U1639 ( n1541,n1542,n1543 );
   not U1640 ( n1543,num_reg_0_ );
   nor U1641 ( n1540,n1544,n1545 );
   not U1642 ( u1572,n1546 );
   nor U1643 ( n1546,n1547,n1548 );
   nor U1644 ( n1548,n1542,n1549 );
   not U1645 ( n1549,num_reg_1_ );
   not U1646 ( n1542,n1544 );
   nor U1647 ( n1547,n1544,n1550 );
   not U1648 ( u1571,n1551 );
   nor U1649 ( n1551,n1552,n1553 );
   nor U1650 ( n1553,n1554,n1555 );
   nor U1651 ( n1555,n1556,n1557 );
   not U1652 ( n1557,n1558 );
   nor U1653 ( n1558,n1559,n1504 );
   nor U1654 ( n1559,n1560,n1561 );
   nor U1655 ( n1556,n1508,n1562 );
   nor U1656 ( n1552,n1563,n1564 );
   not U1657 ( u1570,n1565 );
   nor U1658 ( n1565,n1566,n1567 );
   nor U1659 ( n1567,n1554,n1568 );
   nor U1660 ( n1568,n1569,n1570 );
   nor U1661 ( n1570,n1571,n1560 );
   nor U1662 ( n1569,n1572,n1573 );
   nor U1663 ( n1566,n1574,n1563 );
   not U1664 ( u1569,n1575 );
   nor U1665 ( n1575,n1576,n1577 );
   nor U1666 ( n1577,n1554,n1578 );
   nor U1667 ( n1578,n1579,n1580 );
   nor U1668 ( n1579,n1581,n1582 );
   nor U1669 ( n1576,n1583,n1563 );
   not U1670 ( n1563,n1554 );
   nor U1671 ( n1554,n1584,n1585 );
   not U1672 ( n1585,n1586 );
   nor U1673 ( n1586,n1587,n1522 );
   not U1674 ( n1522,n1588 );
   nor U1675 ( n1588,n1589,n1590 );
   not U1676 ( n1590,n1591 );
   nor U1677 ( n1591,n1592,n1593 );
   nor U1678 ( n1587,n1594,n1478 );
   nor U1679 ( n1594,n1595,n1596 );
   nor U1680 ( n1596,n1582,n1597 );
   not U1681 ( n1584,n1598 );
   nor U1682 ( n1598,n1599,n1538 );
   nor U1683 ( n1538,n1600,n1601 );
   not U1684 ( n1601,n1602 );
   nor U1685 ( n1602,n1603,n1477 );
   not U1686 ( n1600,n1604 );
   nor U1687 ( n1604,n1501,n1605 );
   not U1688 ( u1568,n1606 );
   nor U1689 ( n1606,n1607,n1608 );
   not U1690 ( n1608,n1609 );
   nor U1691 ( n1609,n1610,n1611 );
   nor U1692 ( n1611,n1612,n1613 );
   nor U1693 ( n1613,n1614,n1615 );
   nor U1694 ( n1615,n1616,n1617 );
   nor U1695 ( n1614,n1618,n1478 );
   nor U1696 ( n1618,n1619,n1620 );
   not U1697 ( n1620,n1621 );
   nor U1698 ( n1621,n1622,n1623 );
   nor U1699 ( n1623,n1513,n1617 );
   nor U1700 ( n1622,n1582,n1624 );
   not U1701 ( n1624,n1625 );
   nor U1702 ( n1610,n1626,n1627 );
   not U1703 ( n1627,count_reg2_3_ );
   nor U1704 ( n1607,n1628,n1629 );
   not U1705 ( u1567,n1630 );
   nor U1706 ( n1630,n1631,n1632 );
   nor U1707 ( n1632,n1633,n1634 );
   nor U1708 ( n1634,n1635,n1485 );
   nor U1709 ( n1631,n1636,n1637 );
   not U1710 ( u1566,n1638 );
   nor U1711 ( n1638,n1639,n1640 );
   nor U1712 ( n1640,n1633,n1641 );
   nor U1713 ( n1641,n1642,n1485 );
   not U1714 ( n1642,n1643 );
   nor U1715 ( n1639,n1637,n1644 );
   not U1716 ( u1565,n1645 );
   nor U1717 ( n1645,n1646,n1647 );
   nor U1718 ( n1647,n1648,n1561 );
   not U1719 ( n1561,n1649 );
   nor U1720 ( n1649,k_0_,n1650 );
   nor U1721 ( n1650,k_1_,n1651 );
   nor U1722 ( n1646,n1589,n1652 );
   not U1723 ( u1564,n1653 );
   nor U1724 ( n1653,n1654,n1655 );
   nor U1725 ( n1655,n1571,n1648 );
   not U1726 ( n1648,n1589 );
   nor U1727 ( n1654,n1589,n1656 );
   nor U1728 ( n1589,n1657,n1658 );
   xor U1729 ( n2949,count_reg_1_,count_reg_0_ );
   not U1730 ( u1486,n1659 );
   nor U1731 ( n1659,n1660,n1661 );
   nor U1732 ( n1661,n1662,n1468 );
   nor U1733 ( n1660,n1663,n1664 );
   not U1734 ( u1485,n1665 );
   nor U1735 ( n1665,n1666,n1667 );
   nor U1736 ( n1667,n1662,n1472 );
   nor U1737 ( n1666,n1663,n1668 );
   nor U1738 ( n1663,n1662,n1476 );
   not U1739 ( u1484,n1669 );
   nor U1740 ( n1669,n1670,n1671 );
   nor U1741 ( n1671,n1465,n1672 );
   nor U1742 ( n1670,n1673,n1674 );
   not U1743 ( u1483,n1675 );
   nor U1744 ( n1675,n1676,n1677 );
   nor U1745 ( n1677,n1469,n1672 );
   nor U1746 ( n1676,n1673,n1678 );
   nor U1747 ( n1673,n1475,n1672 );
   not U1748 ( u1482,n1679 );
   nor U1749 ( n1679,n1680,n1681 );
   nor U1750 ( n1681,n1467,n1682 );
   nor U1751 ( n1680,n1683,n1684 );
   not U1752 ( u1481,n1685 );
   nor U1753 ( n1685,n1686,n1687 );
   nor U1754 ( n1687,n1471,n1682 );
   nor U1755 ( n1686,n1683,n1688 );
   nor U1756 ( n1683,n1475,n1682 );
   not U1757 ( u1480,n1689 );
   nor U1758 ( n1689,n1690,n1691 );
   nor U1759 ( n1691,n1467,n1692 );
   nor U1760 ( n1690,n1693,n1694 );
   not U1761 ( u1479,n1695 );
   nor U1762 ( n1695,n1696,n1697 );
   nor U1763 ( n1697,n1471,n1692 );
   nor U1764 ( n1696,n1693,n1698 );
   nor U1765 ( n1693,n1474,n1692 );
   not U1766 ( u1478,n1699 );
   nor U1767 ( n1699,n1700,n1701 );
   nor U1768 ( n1701,n1465,n1702 );
   nor U1769 ( n1700,n1703,n1704 );
   not U1770 ( u1477,n1705 );
   nor U1771 ( n1705,n1706,n1707 );
   nor U1772 ( n1707,n1469,n1702 );
   nor U1773 ( n1706,n1703,n1708 );
   nor U1774 ( n1703,n1474,n1702 );
   not U1775 ( u1476,n1709 );
   nor U1776 ( n1709,n1710,n1711 );
   nor U1777 ( n1711,n1465,n1712 );
   nor U1778 ( n1710,n1713,n1714 );
   not U1779 ( u1475,n1715 );
   nor U1780 ( n1715,n1716,n1717 );
   nor U1781 ( n1717,n1469,n1712 );
   nor U1782 ( n1716,n1713,n1718 );
   nor U1783 ( n1713,n1476,n1712 );
   not U1784 ( u1474,n1719 );
   nor U1785 ( n1719,n1720,n1721 );
   nor U1786 ( n1721,n1468,n1722 );
   nor U1787 ( n1720,n1723,n1724 );
   not U1788 ( u1473,n1725 );
   nor U1789 ( n1725,n1726,n1727 );
   nor U1790 ( n1727,n1472,n1722 );
   nor U1791 ( n1726,n1723,n1728 );
   nor U1792 ( n1723,n1473,n1722 );
   not U1793 ( u1472,n1729 );
   nor U1794 ( n1729,n1730,n1731 );
   nor U1795 ( n1731,n1468,n1732 );
   nor U1796 ( n1730,n1733,n1734 );
   not U1797 ( u1471,n1735 );
   nor U1798 ( n1735,n1736,n1737 );
   nor U1799 ( n1737,n1472,n1732 );
   nor U1800 ( n1736,n1733,n1738 );
   nor U1801 ( n1733,n1474,n1732 );
   not U1802 ( u1470,n1739 );
   nor U1803 ( n1739,n1740,n1741 );
   nor U1804 ( n1741,n1466,n1742 );
   nor U1805 ( n1740,n1743,n1744 );
   not U1806 ( u1469,n1745 );
   nor U1807 ( n1745,n1746,n1747 );
   nor U1808 ( n1747,n1470,n1742 );
   nor U1809 ( n1746,n1743,n1748 );
   nor U1810 ( n1743,n1475,n1742 );
   not U1811 ( u1468,n1749 );
   nor U1812 ( n1749,n1750,n1751 );
   nor U1813 ( n1751,n1466,n1752 );
   nor U1814 ( n1750,n1753,n1754 );
   not U1815 ( u1467,n1755 );
   nor U1816 ( n1755,n1756,n1757 );
   nor U1817 ( n1757,n1470,n1752 );
   nor U1818 ( n1756,n1753,n1758 );
   nor U1819 ( n1753,n1476,n1752 );
   not U1820 ( u1466,n1759 );
   nor U1821 ( n1759,n1760,n1761 );
   nor U1822 ( n1761,n1467,n1762 );
   nor U1823 ( n1760,n1763,n1764 );
   not U1824 ( u1465,n1765 );
   nor U1825 ( n1765,n1766,n1767 );
   nor U1826 ( n1767,n1471,n1762 );
   nor U1827 ( n1766,n1763,n1768 );
   nor U1828 ( n1763,n1473,n1762 );
   not U1829 ( u1464,n1769 );
   nor U1830 ( n1769,n1770,n1771 );
   nor U1831 ( n1771,n1467,n1772 );
   nor U1832 ( n1770,n1773,n1774 );
   not U1833 ( u1463,n1775 );
   nor U1834 ( n1775,n1776,n1777 );
   nor U1835 ( n1777,n1471,n1772 );
   nor U1836 ( n1776,n1773,n1778 );
   nor U1837 ( n1773,n1474,n1772 );
   not U1838 ( u1462,n1779 );
   nor U1839 ( n1779,n1780,n1781 );
   nor U1840 ( n1781,n1466,n1782 );
   nor U1841 ( n1780,n1783,n1784 );
   not U1842 ( u1461,n1785 );
   nor U1843 ( n1785,n1786,n1787 );
   nor U1844 ( n1787,n1470,n1782 );
   nor U1845 ( n1786,n1783,n1788 );
   nor U1846 ( n1783,n1476,n1782 );
   not U1847 ( u1460,n1789 );
   nor U1848 ( n1789,n1790,n1791 );
   nor U1849 ( n1791,n1466,n1792 );
   nor U1850 ( n1790,n1793,n1794 );
   not U1851 ( u1459,n1795 );
   nor U1852 ( n1795,n1796,n1797 );
   nor U1853 ( n1797,n1470,n1792 );
   nor U1854 ( n1796,n1793,n1798 );
   nor U1855 ( n1793,n1475,n1792 );
   not U1856 ( u1458,n1799 );
   nor U1857 ( n1799,n1800,n1801 );
   nor U1858 ( n1801,n1468,n1802 );
   nor U1859 ( n1800,n1803,n1804 );
   not U1860 ( u1457,n1805 );
   nor U1861 ( n1805,n1806,n1807 );
   nor U1862 ( n1807,n1472,n1802 );
   nor U1863 ( n1806,n1803,n1808 );
   nor U1864 ( n1803,n1474,n1802 );
   not U1865 ( u1456,n1809 );
   nor U1866 ( n1809,n1810,n1811 );
   nor U1867 ( n1811,n1468,n1812 );
   nor U1868 ( n1810,n1813,n1814 );
   not U1869 ( u1455,n1815 );
   nor U1870 ( n1815,n1816,n1817 );
   nor U1871 ( n1817,n1472,n1812 );
   nor U1872 ( n1816,n1813,n1818 );
   nor U1873 ( n1813,n1475,n1812 );
   not U1874 ( u1454,n1819 );
   nor U1875 ( n1819,n1820,n1821 );
   nor U1876 ( n1821,n1465,n1822 );
   nor U1877 ( n1820,n1823,n1824 );
   not U1878 ( u1453,n1825 );
   nor U1879 ( n1825,n1826,n1827 );
   nor U1880 ( n1827,n1469,n1822 );
   nor U1881 ( n1826,n1823,n1828 );
   nor U1882 ( n1823,n1473,n1822 );
   not U1883 ( u1452,n1829 );
   nor U1884 ( n1829,n1830,n1831 );
   nor U1885 ( n1831,n1465,n1832 );
   nor U1886 ( n1830,n1833,n1834 );
   not U1887 ( u1451,n1835 );
   nor U1888 ( n1835,n1836,n1837 );
   nor U1889 ( n1837,n1469,n1832 );
   nor U1890 ( n1836,n1833,n1838 );
   nor U1891 ( n1833,n1476,n1832 );
   not U1892 ( u1450,n1839 );
   nor U1893 ( n1839,n1840,n1841 );
   nor U1894 ( n1841,n1467,n1842 );
   nor U1895 ( n1840,n1843,n1844 );
   not U1896 ( u1449,n1845 );
   nor U1897 ( n1845,n1846,n1847 );
   nor U1898 ( n1847,n1471,n1842 );
   nor U1899 ( n1846,n1843,n1848 );
   nor U1900 ( n1843,n1474,n1842 );
   not U1901 ( u1448,n1849 );
   nor U1902 ( n1849,n1850,n1851 );
   nor U1903 ( n1851,n1467,n1852 );
   nor U1904 ( n1850,n1853,n1854 );
   not U1905 ( u1447,n1855 );
   nor U1906 ( n1855,n1856,n1857 );
   nor U1907 ( n1857,n1471,n1852 );
   nor U1908 ( n1856,n1853,n1858 );
   nor U1909 ( n1853,n1473,n1852 );
   not U1910 ( u1446,n1859 );
   nor U1911 ( n1859,n1860,n1861 );
   nor U1912 ( n1861,n1466,n1862 );
   nor U1913 ( n1860,n1863,n1864 );
   not U1914 ( u1445,n1865 );
   nor U1915 ( n1865,n1866,n1867 );
   nor U1916 ( n1867,n1470,n1862 );
   nor U1917 ( n1866,n1863,n1868 );
   nor U1918 ( n1863,n1476,n1862 );
   not U1919 ( u1444,n1869 );
   nor U1920 ( n1869,n1870,n1871 );
   nor U1921 ( n1871,n1468,n1872 );
   nor U1922 ( n1870,n1873,n1874 );
   not U1923 ( u1443,n1875 );
   nor U1924 ( n1875,n1876,n1877 );
   nor U1925 ( n1877,n1472,n1872 );
   nor U1926 ( n1876,n1873,n1878 );
   nor U1927 ( n1873,n1473,n1872 );
   not U1928 ( u1442,n1879 );
   nor U1929 ( n1879,n1880,n1881 );
   nor U1930 ( n1881,n1466,n1882 );
   nor U1931 ( n1880,n1883,n1884 );
   not U1932 ( u1441,n1885 );
   nor U1933 ( n1885,n1886,n1887 );
   nor U1934 ( n1887,n1470,n1882 );
   nor U1935 ( n1886,n1883,n1888 );
   nor U1936 ( n1883,n1473,n1882 );
   not U1937 ( u1440,n1889 );
   nor U1938 ( n1889,n1890,n1891 );
   nor U1939 ( n1891,n1466,n1892 );
   nor U1940 ( n1890,n1893,n1894 );
   not U1941 ( u1439,n1895 );
   nor U1942 ( n1895,n1896,n1897 );
   nor U1943 ( n1897,n1470,n1892 );
   nor U1944 ( n1896,n1893,n1898 );
   nor U1945 ( n1893,n1475,n1892 );
   not U1946 ( u1438,n1899 );
   nor U1947 ( n1899,n1900,n1901 );
   nor U1948 ( n1901,n1465,n1902 );
   nor U1949 ( n1900,n1903,n1904 );
   not U1950 ( u1437,n1905 );
   nor U1951 ( n1905,n1906,n1907 );
   nor U1952 ( n1907,n1469,n1902 );
   nor U1953 ( n1906,n1903,n1908 );
   nor U1954 ( n1903,n1476,n1902 );
   not U1955 ( u1436,n1909 );
   nor U1956 ( n1909,n1910,n1911 );
   nor U1957 ( n1911,n1467,n1912 );
   nor U1958 ( n1910,n1913,n1914 );
   not U1959 ( u1435,n1915 );
   nor U1960 ( n1915,n1916,n1917 );
   nor U1961 ( n1917,n1471,n1912 );
   nor U1962 ( n1916,n1913,n1918 );
   nor U1963 ( n1913,n1473,n1912 );
   not U1964 ( u1434,n1919 );
   nor U1965 ( n1919,n1920,n1921 );
   nor U1966 ( n1921,n1467,n1922 );
   nor U1967 ( n1920,n1923,n1924 );
   not U1968 ( u1433,n1925 );
   nor U1969 ( n1925,n1926,n1927 );
   nor U1970 ( n1927,n1471,n1922 );
   nor U1971 ( n1926,n1923,n1928 );
   nor U1972 ( n1923,n1474,n1922 );
   not U1973 ( u1432,n1929 );
   nor U1974 ( n1929,n1930,n1931 );
   nor U1975 ( n1931,n1465,n1932 );
   nor U1976 ( n1930,n1933,n1934 );
   not U1977 ( u1431,n1935 );
   nor U1978 ( n1935,n1936,n1937 );
   nor U1979 ( n1937,n1469,n1932 );
   nor U1980 ( n1936,n1933,n1938 );
   nor U1981 ( n1933,n1476,n1932 );
   not U1982 ( u1430,n1939 );
   nor U1983 ( n1939,n1940,n1941 );
   nor U1984 ( n1941,n1465,n1942 );
   nor U1985 ( n1940,n1943,n1944 );
   not U1986 ( u1429,n1945 );
   nor U1987 ( n1945,n1946,n1947 );
   nor U1988 ( n1947,n1469,n1942 );
   nor U1989 ( n1946,n1943,n1948 );
   nor U1990 ( n1943,n1475,n1942 );
   not U1991 ( u1428,n1949 );
   nor U1992 ( n1949,n1950,n1951 );
   nor U1993 ( n1951,n1468,n1952 );
   nor U1994 ( n1950,n1953,n1954 );
   not U1995 ( u1427,n1955 );
   nor U1996 ( n1955,n1956,n1957 );
   nor U1997 ( n1957,n1472,n1952 );
   nor U1998 ( n1956,n1953,n1958 );
   nor U1999 ( n1953,n1474,n1952 );
   not U2000 ( u1426,n1959 );
   nor U2001 ( n1959,n1960,n1961 );
   nor U2002 ( n1961,n1468,n1962 );
   nor U2003 ( n1960,n1963,n1964 );
   not U2004 ( u1425,n1965 );
   nor U2005 ( n1965,n1966,n1967 );
   nor U2006 ( n1967,n1472,n1962 );
   nor U2007 ( n1966,n1963,n1968 );
   nor U2008 ( n1963,n1473,n1962 );
   not U2009 ( u1424,n1969 );
   nor U2010 ( n1969,n1970,n1971 );
   nor U2011 ( n1971,n1466,n1972 );
   nor U2012 ( n1973,n1550,n1475 );
   not U2013 ( n1550,data_in_reg_1_ );
   nor U2014 ( n1970,n1974,n1975 );
   not U2015 ( u1423,n1976 );
   nor U2016 ( n1976,n1977,n1978 );
   nor U2017 ( n1978,n1470,n1972 );
   nor U2018 ( n1979,n1545,n1473 );
   not U2019 ( n1545,data_in_reg_0_ );
   nor U2020 ( n1977,n1974,n1980 );
   nor U2021 ( n1974,n1475,n1972 );
   not U2022 ( u1422,n1981 );
   nor U2023 ( n1981,n1982,n1983 );
   not U2024 ( n1983,n1984 );
   nor U2025 ( n1984,n1985,n1986 );
   nor U2026 ( n1986,n1987,n1988 );
   not U2027 ( n1988,nl_reg_3_ );
   nor U2028 ( n1985,n1989,n1990 );
   not U2029 ( n1990,n1991 );
   nor U2030 ( n1991,n1652,n1656 );
   not U2031 ( n1982,n1992 );
   nor U2032 ( n1992,n1993,n1994 );
   nor U2033 ( n1994,n1995,n1996 );
   not U2034 ( n1996,n1997 );
   not U2035 ( u1421,n1998 );
   nor U2036 ( n1998,n1999,n2000 );
   not U2037 ( n2000,n2001 );
   nor U2038 ( n2001,n2002,n2003 );
   nor U2039 ( n2003,n1987,n2004 );
   not U2040 ( n2004,nl_reg_2_ );
   nor U2041 ( n2002,n1989,n2005 );
   not U2042 ( n2005,n2006 );
   nor U2043 ( n2006,ind_reg_0_,n1656 );
   not U2044 ( n1656,ind_reg_1_ );
   not U2045 ( n1999,n2007 );
   nor U2046 ( n2007,n1993,n2008 );
   nor U2047 ( n2008,n1995,n2009 );
   not U2048 ( n2009,n2010 );
   not U2049 ( u1420,n2011 );
   nor U2050 ( n2011,n2012,n2013 );
   not U2051 ( n2013,n2014 );
   nor U2052 ( n2014,n2015,n2016 );
   nor U2053 ( n2016,n1987,n2017 );
   not U2054 ( n2017,nl_reg_1_ );
   nor U2055 ( n2015,n1989,n2018 );
   not U2056 ( n2018,n2019 );
   nor U2057 ( n2019,ind_reg_1_,n1652 );
   not U2058 ( n1652,ind_reg_0_ );
   not U2059 ( n2012,n2020 );
   nor U2060 ( n2020,n1993,n2021 );
   nor U2061 ( n2021,n1995,n2022 );
   not U2062 ( n2022,n2023 );
   nor U2063 ( n2023,data_out_reg_1_,n1562 );
   not U2064 ( u1419,n2024 );
   nor U2065 ( n2024,n2025,n2026 );
   not U2066 ( n2026,n2027 );
   nor U2067 ( n2027,n2028,n2029 );
   nor U2068 ( n2029,n1987,n2030 );
   not U2069 ( n2030,nl_reg_0_ );
   nor U2070 ( n1987,n2031,n2032 );
   not U2071 ( n2032,n2033 );
   nor U2072 ( n2033,n2034,n2035 );
   not U2073 ( n2031,n2036 );
   nor U2074 ( n2028,n1989,n2037 );
   not U2075 ( n2037,n2038 );
   nor U2076 ( n2038,ind_reg_1_,ind_reg_0_ );
   not U2077 ( n1989,n2039 );
   nor U2078 ( n2039,n2034,n2040 );
   not U2079 ( n2040,n2035 );
   nor U2080 ( n2035,n2041,n1485 );
   nor U2081 ( n2041,n2042,n2043 );
   not U2082 ( n2025,n2044 );
   nor U2083 ( n2044,n1993,n2045 );
   nor U2084 ( n2045,n1995,n2046 );
   not U2085 ( n2046,n2047 );
   nor U2086 ( n2047,data_out_reg_1_,data_out_reg_0_ );
   not U2087 ( n1995,n2048 );
   nor U2088 ( n2048,n2034,n2036 );
   nor U2089 ( n2036,n2049,n2050 );
   not U2090 ( n2050,n2051 );
   nor U2091 ( n2051,n2052,n2053 );
   nor U2092 ( n2049,n2054,n1582 );
   nor U2093 ( n1993,n2055,n2056 );
   not U2094 ( n2056,n2057 );
   nor U2095 ( n2057,n2034,n2058 );
   nor U2096 ( n2034,n2059,n2060 );
   not U2097 ( n2060,n2061 );
   nor U2098 ( n2061,n2062,n2063 );
   not U2099 ( n2063,n2064 );
   nor U2100 ( n2064,n2065,n2066 );
   nor U2101 ( n2066,n1513,n2067 );
   not U2102 ( n2067,n2068 );
   nor U2103 ( n2068,n2069,n1603 );
   nor U2104 ( n2065,n1597,n2070 );
   nor U2105 ( n2062,n1514,n2071 );
   not U2106 ( n2071,n2072 );
   not U2107 ( n2059,n2073 );
   nor U2108 ( n2073,n2074,n2075 );
   not U2109 ( n2075,n2076 );
   nor U2110 ( n2076,n2077,n1534 );
   nor U2111 ( n2077,n2078,n1478 );
   nor U2112 ( n2078,n2079,n2080 );
   nor U2113 ( n2080,n2081,n2082 );
   not U2114 ( n2074,n2083 );
   nor U2115 ( n2083,n1593,n1537 );
   nor U2116 ( n1537,n2084,n2085 );
   not U2117 ( n2085,n2086 );
   nor U2118 ( n2086,n1524,n1582 );
   not U2119 ( n2084,n2054 );
   nor U2120 ( n2054,n2087,n1581 );
   not U2121 ( u1418,n2088 );
   nor U2122 ( n2088,n2089,n2090 );
   nor U2123 ( n2090,scan_reg_4_,n2091 );
   not U2124 ( n2091,n2092 );
   nor U2125 ( n2092,n2093,n2094 );
   not U2126 ( n2094,n2095 );
   nor U2127 ( n2095,n2096,n2097 );
   nor U2128 ( n2089,n2098,n2099 );
   nor U2129 ( n2098,n2100,n2101 );
   not U2130 ( n2101,n2102 );
   nor U2131 ( n2100,scan_reg_3_,n2093 );
   not U2132 ( u1417,n2103 );
   nor U2133 ( n2103,n2104,n2105 );
   nor U2134 ( n2105,scan_reg_3_,n2106 );
   not U2135 ( n2106,n2107 );
   nor U2136 ( n2107,n2097,n2093 );
   not U2137 ( n2097,n2108 );
   nor U2138 ( n2104,n2102,n2096 );
   nor U2139 ( n2102,n2109,n2110 );
   nor U2140 ( n2109,n2108,n2093 );
   nor U2141 ( n2108,n2111,n2112 );
   not U2142 ( u1416,n2113 );
   nor U2143 ( n2113,n2114,n2115 );
   nor U2144 ( n2115,scan_reg_2_,n2116 );
   not U2145 ( n2116,n2117 );
   nor U2146 ( n2117,n2093,n2112 );
   not U2147 ( n2112,n2118 );
   nor U2148 ( n2118,n2119,n2120 );
   nor U2149 ( n2114,n2121,n2111 );
   nor U2150 ( n2121,n2122,n2123 );
   not U2151 ( n2123,n2124 );
   nor U2152 ( n2122,scan_reg_1_,n2093 );
   not U2153 ( u1415,n2125 );
   nor U2154 ( n2125,n2126,n2127 );
   nor U2155 ( n2127,scan_reg_1_,n2128 );
   not U2156 ( n2128,n2129 );
   nor U2157 ( n2129,n2120,n2093 );
   nor U2158 ( n2126,n2124,n2119 );
   nor U2159 ( n2124,n2130,n2110 );
   not U2160 ( u1414,n2131 );
   nor U2161 ( n2131,n2130,n2132 );
   nor U2162 ( n2132,n2120,n2133 );
   not U2163 ( n2133,n2110 );
   nor U2164 ( n2130,scan_reg_0_,n2093 );
   not U2165 ( n2093,n2134 );
   nor U2166 ( n2134,n1513,n2135 );
   not U2167 ( n2135,n2136 );
   nor U2168 ( n2136,n2137,n2110 );
   nor U2169 ( n2110,n2138,n2139 );
   not U2170 ( n2139,n2140 );
   nor U2171 ( n2140,n2141,n1544 );
   nor U2172 ( n2138,n1524,n2142 );
   not U2173 ( u1413,n2143 );
   nor U2174 ( n2143,n2144,n2145 );
   nor U2175 ( n2145,max_reg_4_,n2146 );
   not U2176 ( n2146,n2147 );
   nor U2177 ( n2147,n2148,n2149 );
   not U2178 ( n2149,n2150 );
   nor U2179 ( n2150,n2151,n2152 );
   nor U2180 ( n2144,n2153,n2154 );
   nor U2181 ( n2153,n2155,n2156 );
   not U2182 ( n2156,n2157 );
   nor U2183 ( n2155,max_reg_3_,n2148 );
   not U2184 ( u1412,n2158 );
   nor U2185 ( n2158,n2159,n2160 );
   nor U2186 ( n2160,max_reg_3_,n2161 );
   not U2187 ( n2161,n2162 );
   nor U2188 ( n2162,n2152,n2148 );
   nor U2189 ( n2159,n2157,n2151 );
   nor U2190 ( n2157,n2163,n2164 );
   nor U2191 ( n2163,n2165,n2148 );
   not U2192 ( u1411,n2166 );
   nor U2193 ( n2166,n2167,n2168 );
   nor U2194 ( n2168,max_reg_2_,n2169 );
   not U2195 ( n2169,n2170 );
   nor U2196 ( n2170,n2148,n2171 );
   nor U2197 ( n2167,n2172,n2173 );
   nor U2198 ( n2172,n2174,n2175 );
   not U2199 ( n2175,n2176 );
   nor U2200 ( n2174,max_reg_1_,n2148 );
   not U2201 ( u1410,n2177 );
   nor U2202 ( n2177,n2178,n2179 );
   nor U2203 ( n2179,max_reg_1_,n2180 );
   not U2204 ( n2180,n2181 );
   nor U2205 ( n2181,n2182,n2148 );
   nor U2206 ( n2178,n2176,n2183 );
   nor U2207 ( n2176,n2184,n2164 );
   not U2208 ( u1409,n2185 );
   nor U2209 ( n2185,n2184,n2186 );
   nor U2210 ( n2186,n2182,n2187 );
   not U2211 ( n2187,n2164 );
   nor U2212 ( n2184,max_reg_0_,n2148 );
   not U2213 ( n2148,n2188 );
   nor U2214 ( n2188,n2164,n1513 );
   nor U2215 ( n2164,n2189,n1637 );
   nor U2216 ( n2189,n2190,n1478 );
   nor U2217 ( n2190,n2191,n2192 );
   nor U2218 ( n2191,n2193,n2194 );
   not U2219 ( u1408,n2195 );
   nor U2220 ( n2195,n2196,n2197 );
   nor U2221 ( n2197,n1637,n2198 );
   nor U2222 ( n2196,n2199,n2200 );
   not U2223 ( u1407,n2201 );
   nor U2224 ( n2201,n2202,n2203 );
   nor U2225 ( n2203,n1617,n1637 );
   nor U2226 ( n2202,n1628,n2200 );
   nor U2227 ( n1628,n2204,n2205 );
   nor U2228 ( n2205,n2206,n2207 );
   not U2229 ( u1406,n2208 );
   nor U2230 ( n2208,n2209,n2210 );
   nor U2231 ( n2210,n2211,n1637 );
   nor U2232 ( n2209,n2212,n2200 );
   not U2233 ( u1405,n2213 );
   nor U2234 ( n2213,n2214,n2215 );
   nor U2235 ( n2215,n2216,n1637 );
   not U2236 ( n1637,n1633 );
   nor U2237 ( n2214,n2217,n2200 );
   not U2238 ( n2200,n2218 );
   nor U2239 ( n2218,n1633,n1485 );
   nor U2240 ( n1633,n2219,n1486 );
   nor U2241 ( n1486,n1560,n2069 );
   not U2242 ( u1404,n2220 );
   nor U2243 ( n2220,n2221,n2222 );
   not U2244 ( n2222,n2223 );
   nor U2245 ( n2223,n2224,n2225 );
   nor U2246 ( n2225,n1612,n2226 );
   nor U2247 ( n2226,n2227,n2228 );
   nor U2248 ( n2228,n2229,n1643 );
   xor U2249 ( n1643,n2230,n2231 );
   nor U2250 ( n2231,count_reg2_5_,n2232 );
   nor U2251 ( n2232,n1524,n1644 );
   nor U2252 ( n2230,n2233,n2234 );
   nor U2253 ( n2227,n2235,n1644 );
   not U2254 ( n1644,timebase_reg_5_ );
   nor U2255 ( n2224,n1626,n2236 );
   not U2256 ( n2236,count_reg2_5_ );
   not U2257 ( u1403,n2237 );
   nor U2258 ( n2237,n2238,n2239 );
   not U2259 ( n2239,n2240 );
   nor U2260 ( n2240,n2241,n2242 );
   nor U2261 ( n2242,n2198,n2243 );
   nor U2262 ( n2241,n1629,n2199 );
   xor U2263 ( n2199,n2234,n2233 );
   not U2264 ( n2233,n2244 );
   nor U2265 ( n2244,count_reg2_4_,n2245 );
   nor U2266 ( n2245,n1524,n2198 );
   not U2267 ( n2198,timebase_reg_4_ );
   not U2268 ( n2234,n2204 );
   nor U2269 ( n2204,n2246,n2247 );
   not U2270 ( n2247,n2206 );
   nor U2271 ( n2206,count_reg2_3_,n2248 );
   nor U2272 ( n2248,n1524,n1617 );
   not U2273 ( n1617,timebase_reg_3_ );
   not U2274 ( n2246,n2207 );
   nor U2275 ( n2238,n1626,n2249 );
   not U2276 ( n2249,count_reg2_4_ );
   not U2277 ( u1402,n2250 );
   nor U2278 ( n2250,n2251,n2252 );
   not U2279 ( n2252,n2253 );
   nor U2280 ( n2253,n2254,n2255 );
   nor U2281 ( n2255,n2211,n2243 );
   nor U2282 ( n2254,n2212,n1629 );
   nor U2283 ( n2212,n2207,n2256 );
   nor U2284 ( n2256,n2257,n2258 );
   nor U2285 ( n2207,n2259,n2260 );
   not U2286 ( n2260,n2257 );
   nor U2287 ( n2257,count_reg2_2_,n2261 );
   nor U2288 ( n2261,n1478,n2211 );
   not U2289 ( n2211,timebase_reg_2_ );
   not U2290 ( n2259,n2258 );
   nor U2291 ( n2251,n1626,n2262 );
   not U2292 ( n2262,count_reg2_2_ );
   not U2293 ( u1401,n2263 );
   nor U2294 ( n2263,n2264,n2265 );
   not U2295 ( n2265,n2266 );
   nor U2296 ( n2266,n2267,n2268 );
   nor U2297 ( n2268,n2216,n2243 );
   not U2298 ( n2243,n2269 );
   nor U2299 ( n2269,n1612,n2270 );
   nor U2300 ( n2270,n2271,n2272 );
   not U2301 ( n2272,n1616 );
   nor U2302 ( n1616,n2273,n2274 );
   not U2303 ( n2274,n2275 );
   nor U2304 ( n2275,n2276,n2277 );
   nor U2305 ( n2277,n1560,n2278 );
   not U2306 ( n2278,n2279 );
   nor U2307 ( n2279,n1657,n2280 );
   not U2308 ( n2273,n1572 );
   nor U2309 ( n1572,n2281,n2053 );
   nor U2310 ( n2267,n2217,n1629 );
   not U2311 ( n1629,n2282 );
   nor U2312 ( n2282,n1612,n2283 );
   nor U2313 ( n2283,n2284,n2285 );
   not U2314 ( n2285,n2286 );
   nor U2315 ( n2286,n2287,n2288 );
   nor U2316 ( n2288,n2289,n2290 );
   not U2317 ( n2290,n2291 );
   nor U2318 ( n2291,n2280,n1560 );
   nor U2319 ( n2284,n1513,n2292 );
   not U2320 ( n2292,n2293 );
   nor U2321 ( n2293,n2081,n2294 );
   nor U2322 ( n2217,n2258,n2295 );
   nor U2323 ( n2295,n2296,n1635 );
   nor U2324 ( n2258,n2297,n2298 );
   not U2325 ( n2298,n2296 );
   nor U2326 ( n2296,count_reg2_1_,n2299 );
   nor U2327 ( n2299,n1524,n2216 );
   not U2328 ( n2216,timebase_reg_1_ );
   nor U2329 ( n2264,n1626,n2300 );
   not U2330 ( n2300,count_reg2_1_ );
   not U2331 ( u1400,n2301 );
   nor U2332 ( n2301,n2221,n2302 );
   not U2333 ( n2302,n2303 );
   nor U2334 ( n2303,n2304,n2305 );
   nor U2335 ( n2305,n1612,n2306 );
   nor U2336 ( n2306,n2307,n2308 );
   nor U2337 ( n2308,n2229,n2297 );
   not U2338 ( n2297,n1635 );
   nor U2339 ( n1635,count_reg2_0_,n2309 );
   nor U2340 ( n2309,n1524,n1636 );
   nor U2341 ( n2229,n2310,n2311 );
   not U2342 ( n2311,n2312 );
   nor U2343 ( n2312,n2287,n2313 );
   nor U2344 ( n2313,n1560,n2289 );
   not U2345 ( n2289,n1657 );
   nor U2346 ( n2287,n2294,n2314 );
   nor U2347 ( n2314,n2315,n1619 );
   not U2348 ( n1619,n2316 );
   nor U2349 ( n2316,n2317,n2318 );
   not U2350 ( n2318,n2319 );
   nor U2351 ( n2319,n1507,n2320 );
   nor U2352 ( n2317,n1485,n1501 );
   nor U2353 ( n2315,n1508,n2058 );
   nor U2354 ( n2310,n2321,n2294 );
   nor U2355 ( n2321,n2322,n1625 );
   nor U2356 ( n1625,n2280,n1477 );
   nor U2357 ( n2307,n2235,n1636 );
   not U2358 ( n1636,timebase_reg_0_ );
   nor U2359 ( n2235,n2323,n2324 );
   not U2360 ( n2324,n2325 );
   nor U2361 ( n2325,n2326,n2327 );
   nor U2362 ( n2327,n1657,n1560 );
   nor U2363 ( n1657,n1571,n2328 );
   not U2364 ( n2328,n2329 );
   nor U2365 ( n2329,k_3_,k_2_ );
   nor U2366 ( n2326,n2330,n2331 );
   not U2367 ( n2323,n2332 );
   nor U2368 ( n2332,n2271,n2333 );
   not U2369 ( n2333,n2334 );
   nor U2370 ( n2334,n2281,n2276 );
   nor U2371 ( n2276,n2335,n1478 );
   nor U2372 ( n2335,n2336,n2337 );
   nor U2373 ( n2336,n2280,n2082 );
   nor U2374 ( n2281,n2280,n2193 );
   nor U2375 ( n2271,n2338,n2339 );
   not U2376 ( n2339,n2340 );
   nor U2377 ( n2340,n1524,n1477 );
   nor U2378 ( n2304,n1626,n2341 );
   not U2379 ( n2341,count_reg2_0_ );
   not U2380 ( n1626,n1612 );
   nor U2381 ( n2221,n1560,n2342 );
   not U2382 ( n2342,n2343 );
   nor U2383 ( n2343,n2330,n1612 );
   nor U2384 ( n1612,n2344,n2345 );
   not U2385 ( n2345,n2346 );
   nor U2386 ( n2346,n2347,n2348 );
   not U2387 ( n2348,n2349 );
   nor U2388 ( n2349,n2350,n2351 );
   not U2389 ( n2351,n2352 );
   nor U2390 ( n2352,n2353,n2354 );
   nor U2391 ( n2354,n2058,n2355 );
   not U2392 ( n2355,n2356 );
   nor U2393 ( n2356,n2294,n2357 );
   nor U2394 ( n2353,n1512,n2358 );
   not U2395 ( n2358,n2053 );
   nor U2396 ( n2053,n2331,n2359 );
   not U2397 ( n2350,n2360 );
   nor U2398 ( n2360,n2361,n2362 );
   nor U2399 ( n2362,n1506,n2363 );
   not U2400 ( n2363,n2364 );
   nor U2401 ( n2364,n2330,n2055 );
   nor U2402 ( n2361,n2365,n1477 );
   nor U2403 ( n2365,n2366,n2367 );
   not U2404 ( n2367,n2368 );
   nor U2405 ( n2368,n2369,n2370 );
   nor U2406 ( n2370,n1582,n2371 );
   not U2407 ( n2371,n2372 );
   nor U2408 ( n2372,n2081,n1508 );
   nor U2409 ( n2369,n1514,n2373 );
   not U2410 ( n2373,n2374 );
   nor U2411 ( n2374,n2294,n1597 );
   nor U2412 ( n2366,n2280,n2375 );
   not U2413 ( n2347,n2376 );
   nor U2414 ( n2376,n2377,n2378 );
   nor U2415 ( n2377,n1506,n2194 );
   not U2416 ( n2344,n2379 );
   nor U2417 ( n2379,n2380,n2381 );
   not U2418 ( n2381,n2382 );
   nor U2419 ( n2382,n2383,n2384 );
   nor U2420 ( n2384,n1514,n2385 );
   nor U2421 ( n2383,n2338,n2386 );
   not U2422 ( n2386,n2387 );
   nor U2423 ( n2387,n1514,n1485 );
   not U2424 ( n2380,n2388 );
   nor U2425 ( n2388,n2389,n1593 );
   nor U2426 ( n1593,n1597,n2390 );
   not U2427 ( n2390,n2391 );
   nor U2428 ( n2391,n2193,n1582 );
   not U2429 ( u1399,n2392 );
   nor U2430 ( n2392,n2393,n2394 );
   not U2431 ( n2394,n2395 );
   nor U2432 ( n2395,n2396,n2397 );
   nor U2433 ( n2397,n2154,n2398 );
   nor U2434 ( n2396,n2099,n2399 );
   nor U2435 ( n2393,n2400,n2401 );
   not U2436 ( u1398,n2402 );
   nor U2437 ( n2402,n2403,n2404 );
   not U2438 ( n2404,n2405 );
   nor U2439 ( n2405,n2406,n2407 );
   nor U2440 ( n2407,n2151,n2398 );
   nor U2441 ( n2406,n2096,n2399 );
   nor U2442 ( n2403,n2408,n2401 );
   not U2443 ( u1397,n2409 );
   nor U2444 ( n2409,n2410,n2411 );
   not U2445 ( n2411,n2412 );
   nor U2446 ( n2412,n2413,n2414 );
   nor U2447 ( n2414,n2173,n2398 );
   nor U2448 ( n2413,n2111,n2399 );
   nor U2449 ( n2410,n2415,n2401 );
   not U2450 ( u1396,n2416 );
   nor U2451 ( n2416,n2417,n2418 );
   not U2452 ( n2418,n2419 );
   nor U2453 ( n2419,n2420,n2421 );
   nor U2454 ( n2421,n2183,n2398 );
   nor U2455 ( n2420,n2119,n2399 );
   nor U2456 ( n2417,n2422,n2401 );
   not U2457 ( u1395,n2423 );
   nor U2458 ( n2423,n2424,n2425 );
   not U2459 ( n2425,n2426 );
   nor U2460 ( n2426,n2427,n2428 );
   nor U2461 ( n2428,n2182,n2398 );
   not U2462 ( n2398,n2429 );
   nor U2463 ( n2429,n2430,n2431 );
   nor U2464 ( n2431,n2320,n2042 );
   nor U2465 ( n2427,n2120,n2399 );
   not U2466 ( n2399,n2432 );
   nor U2467 ( n2432,n2430,n2433 );
   nor U2468 ( n2433,n1511,n1508 );
   nor U2469 ( n2424,n2434,n2401 );
   not U2470 ( n2401,n2430 );
   nor U2471 ( n2430,n2435,n2436 );
   nor U2472 ( n2436,n2437,n2193 );
   nor U2473 ( n2437,n2320,n2438 );
   nor U2474 ( n2438,n1514,n2280 );
   not U2475 ( u1394,n2439 );
   nor U2476 ( n2439,n2440,n2441 );
   nor U2477 ( n2440,n2442,n2443 );
   not U2478 ( n2443,s_reg );
   nor U2479 ( n2442,n1516,n2444 );
   not U2480 ( u1393,n2445 );
   nor U2481 ( n2445,n2446,n2441 );
   nor U2482 ( n2441,n2444,n2447 );
   not U2483 ( n2447,n2448 );
   nor U2484 ( n2448,s_reg,n1516 );
   not U2485 ( n2444,n2449 );
   nor U2486 ( n2446,n2450,n2451 );
   not U2487 ( n2451,n2452 );
   nor U2488 ( n2452,n2449,n1516 );
   nor U2489 ( n2449,n2453,n2454 );
   not U2490 ( n2450,speaker_reg );
   not U2491 ( u1392,n2455 );
   nor U2492 ( n2455,n2456,n1544 );
   nor U2493 ( n1544,n2375,n2457 );
   not U2494 ( n2457,n2458 );
   nor U2495 ( n2458,n1506,n2280 );
   nor U2496 ( n2456,n2459,n1474 );
   nor U2497 ( n2459,n1560,n2460 );
   not U2498 ( n2460,n2461 );
   nor U2499 ( n2461,n1512,n1508 );
   not U2500 ( u1391,count_reg_0_ );
   not U2501 ( u1390,n2462 );
   nor U2502 ( n2462,n2463,n2464 );
   not U2503 ( n2464,n2465 );
   nor U2504 ( n2465,n2466,n2467 );
   not U2505 ( n2467,n2468 );
   nor U2506 ( n2468,n2469,n2470 );
   not U2507 ( n2470,n2471 );
   nor U2508 ( n2471,n2472,n2473 );
   not U2509 ( n2473,n2474 );
   nor U2510 ( n2474,n2475,n2476 );
   nor U2511 ( n2476,n1972,n1975 );
   not U2512 ( n1975,memory_reg_0__1_ );
   nor U2513 ( n2475,n1962,n1964 );
   not U2514 ( n1964,memory_reg_1__1_ );
   not U2515 ( n2472,n2477 );
   nor U2516 ( n2477,n2478,n2479 );
   nor U2517 ( n2479,n1952,n1954 );
   not U2518 ( n1954,memory_reg_2__1_ );
   nor U2519 ( n2478,n1942,n1944 );
   not U2520 ( n1944,memory_reg_3__1_ );
   not U2521 ( n2469,n2480 );
   nor U2522 ( n2480,n2481,n2482 );
   not U2523 ( n2482,n2483 );
   nor U2524 ( n2483,n2484,n2485 );
   nor U2525 ( n2485,n1932,n1934 );
   not U2526 ( n1934,memory_reg_4__1_ );
   nor U2527 ( n2484,n1922,n1924 );
   not U2528 ( n1924,memory_reg_5__1_ );
   not U2529 ( n2481,n2486 );
   nor U2530 ( n2486,n2487,n2488 );
   nor U2531 ( n2488,n1912,n1914 );
   not U2532 ( n1914,memory_reg_6__1_ );
   nor U2533 ( n2487,n1902,n1904 );
   not U2534 ( n1904,memory_reg_7__1_ );
   not U2535 ( n2466,n2489 );
   nor U2536 ( n2489,n2490,n2491 );
   not U2537 ( n2491,n2492 );
   nor U2538 ( n2492,n2493,n2494 );
   not U2539 ( n2494,n2495 );
   nor U2540 ( n2495,n2496,n2497 );
   nor U2541 ( n2497,n1892,n1894 );
   not U2542 ( n1894,memory_reg_8__1_ );
   nor U2543 ( n2496,n1882,n1884 );
   not U2544 ( n1884,memory_reg_9__1_ );
   not U2545 ( n2493,n2498 );
   nor U2546 ( n2498,n2499,n2500 );
   nor U2547 ( n2500,n1872,n1874 );
   not U2548 ( n1874,memory_reg_10__1_ );
   nor U2549 ( n2499,n1862,n1864 );
   not U2550 ( n1864,memory_reg_11__1_ );
   not U2551 ( n2490,n2501 );
   nor U2552 ( n2501,n2502,n2503 );
   not U2553 ( n2503,n2504 );
   nor U2554 ( n2504,n2505,n2506 );
   nor U2555 ( n2506,n1852,n1854 );
   not U2556 ( n1854,memory_reg_12__1_ );
   nor U2557 ( n2505,n1842,n1844 );
   not U2558 ( n1844,memory_reg_13__1_ );
   not U2559 ( n2502,n2507 );
   nor U2560 ( n2507,n2508,n2509 );
   nor U2561 ( n2509,n1832,n1834 );
   not U2562 ( n1834,memory_reg_14__1_ );
   nor U2563 ( n2508,n1822,n1824 );
   not U2564 ( n1824,memory_reg_15__1_ );
   not U2565 ( n2463,n2510 );
   nor U2566 ( n2510,n2511,n2512 );
   not U2567 ( n2512,n2513 );
   nor U2568 ( n2513,n2514,n2515 );
   not U2569 ( n2515,n2516 );
   nor U2570 ( n2516,n2517,n2518 );
   not U2571 ( n2518,n2519 );
   nor U2572 ( n2519,n2520,n2521 );
   nor U2573 ( n2521,n1812,n1814 );
   not U2574 ( n1814,memory_reg_16__1_ );
   nor U2575 ( n2520,n1802,n1804 );
   not U2576 ( n1804,memory_reg_17__1_ );
   not U2577 ( n2517,n2522 );
   nor U2578 ( n2522,n2523,n2524 );
   nor U2579 ( n2524,n1792,n1794 );
   not U2580 ( n1794,memory_reg_18__1_ );
   nor U2581 ( n2523,n1782,n1784 );
   not U2582 ( n1784,memory_reg_19__1_ );
   not U2583 ( n2514,n2525 );
   nor U2584 ( n2525,n2526,n2527 );
   not U2585 ( n2527,n2528 );
   nor U2586 ( n2528,n2529,n2530 );
   nor U2587 ( n2530,n1772,n1774 );
   not U2588 ( n1774,memory_reg_20__1_ );
   nor U2589 ( n2529,n1762,n1764 );
   not U2590 ( n1764,memory_reg_21__1_ );
   not U2591 ( n2526,n2531 );
   nor U2592 ( n2531,n2532,n2533 );
   nor U2593 ( n2533,n1752,n1754 );
   not U2594 ( n1754,memory_reg_22__1_ );
   nor U2595 ( n2532,n1742,n1744 );
   not U2596 ( n1744,memory_reg_23__1_ );
   not U2597 ( n2511,n2534 );
   nor U2598 ( n2534,n2535,n2536 );
   not U2599 ( n2536,n2537 );
   nor U2600 ( n2537,n2538,n2539 );
   not U2601 ( n2539,n2540 );
   nor U2602 ( n2540,n2541,n2542 );
   nor U2603 ( n2542,n1732,n1734 );
   not U2604 ( n1734,memory_reg_24__1_ );
   nor U2605 ( n2541,n1722,n1724 );
   not U2606 ( n1724,memory_reg_25__1_ );
   not U2607 ( n2538,n2543 );
   nor U2608 ( n2543,n2544,n2545 );
   nor U2609 ( n2545,n1712,n1714 );
   not U2610 ( n1714,memory_reg_26__1_ );
   nor U2611 ( n2544,n1702,n1704 );
   not U2612 ( n1704,memory_reg_27__1_ );
   not U2613 ( n2535,n2546 );
   nor U2614 ( n2546,n2547,n2548 );
   not U2615 ( n2548,n2549 );
   nor U2616 ( n2549,n2550,n2551 );
   nor U2617 ( n2551,n1692,n1694 );
   not U2618 ( n1694,memory_reg_28__1_ );
   nor U2619 ( n2550,n1682,n1684 );
   not U2620 ( n1684,memory_reg_29__1_ );
   not U2621 ( n2547,n2552 );
   nor U2622 ( n2552,n2553,n2554 );
   nor U2623 ( n2554,n1672,n1674 );
   not U2624 ( n1674,memory_reg_30__1_ );
   nor U2625 ( n2553,n1662,n1664 );
   not U2626 ( n1664,memory_reg_31__1_ );
   not U2627 ( u1389,n2555 );
   nor U2628 ( n2555,n2556,n2557 );
   not U2629 ( n2557,n2558 );
   nor U2630 ( n2558,n2559,n2560 );
   not U2631 ( n2560,n2561 );
   nor U2632 ( n2561,n2562,n2563 );
   not U2633 ( n2563,n2564 );
   nor U2634 ( n2564,n2565,n2566 );
   not U2635 ( n2566,n2567 );
   nor U2636 ( n2567,n2568,n2569 );
   nor U2637 ( n2569,n1972,n1980 );
   not U2638 ( n1980,memory_reg_0__0_ );
   not U2639 ( n1972,n2570 );
   nor U2640 ( n2570,n2571,n2572 );
   nor U2641 ( n2568,n1962,n1968 );
   not U2642 ( n1968,memory_reg_1__0_ );
   not U2643 ( n1962,n2573 );
   nor U2644 ( n2573,n2574,n2572 );
   not U2645 ( n2565,n2575 );
   nor U2646 ( n2575,n2576,n2577 );
   nor U2647 ( n2577,n1952,n1958 );
   not U2648 ( n1958,memory_reg_2__0_ );
   not U2649 ( n1952,n2578 );
   nor U2650 ( n2578,n2571,n2579 );
   nor U2651 ( n2576,n1942,n1948 );
   not U2652 ( n1948,memory_reg_3__0_ );
   not U2653 ( n1942,n2580 );
   nor U2654 ( n2580,n2574,n2579 );
   not U2655 ( n2562,n2581 );
   nor U2656 ( n2581,n2582,n2583 );
   not U2657 ( n2583,n2584 );
   nor U2658 ( n2584,n2585,n2586 );
   nor U2659 ( n2586,n1932,n1938 );
   not U2660 ( n1938,memory_reg_4__0_ );
   not U2661 ( n1932,n2587 );
   nor U2662 ( n2587,n2588,n2572 );
   nor U2663 ( n2585,n1922,n1928 );
   not U2664 ( n1928,memory_reg_5__0_ );
   not U2665 ( n1922,n2589 );
   nor U2666 ( n2589,n2590,n2572 );
   not U2667 ( n2572,n2591 );
   nor U2668 ( n2591,address_reg_1_,n2592 );
   not U2669 ( n2582,n2593 );
   nor U2670 ( n2593,n2594,n2595 );
   nor U2671 ( n2595,n1912,n1918 );
   not U2672 ( n1918,memory_reg_6__0_ );
   not U2673 ( n1912,n2596 );
   nor U2674 ( n2596,n2588,n2579 );
   nor U2675 ( n2594,n1902,n1908 );
   not U2676 ( n1908,memory_reg_7__0_ );
   not U2677 ( n1902,n2597 );
   nor U2678 ( n2597,n2590,n2579 );
   not U2679 ( n2579,n2598 );
   nor U2680 ( n2598,n2422,n2592 );
   not U2681 ( n2592,n2599 );
   nor U2682 ( n2599,address_reg_4_,address_reg_3_ );
   not U2683 ( n2559,n2600 );
   nor U2684 ( n2600,n2601,n2602 );
   not U2685 ( n2602,n2603 );
   nor U2686 ( n2603,n2604,n2605 );
   not U2687 ( n2605,n2606 );
   nor U2688 ( n2606,n2607,n2608 );
   nor U2689 ( n2608,n1892,n1898 );
   not U2690 ( n1898,memory_reg_8__0_ );
   not U2691 ( n1892,n2609 );
   nor U2692 ( n2609,n2571,n2610 );
   nor U2693 ( n2607,n1882,n1888 );
   not U2694 ( n1888,memory_reg_9__0_ );
   not U2695 ( n1882,n2611 );
   nor U2696 ( n2611,n2574,n2610 );
   not U2697 ( n2604,n2612 );
   nor U2698 ( n2612,n2613,n2614 );
   nor U2699 ( n2614,n1872,n1878 );
   not U2700 ( n1878,memory_reg_10__0_ );
   not U2701 ( n1872,n2615 );
   nor U2702 ( n2615,n2571,n2616 );
   nor U2703 ( n2613,n1862,n1868 );
   not U2704 ( n1868,memory_reg_11__0_ );
   not U2705 ( n1862,n2617 );
   nor U2706 ( n2617,n2574,n2616 );
   not U2707 ( n2601,n2618 );
   nor U2708 ( n2618,n2619,n2620 );
   not U2709 ( n2620,n2621 );
   nor U2710 ( n2621,n2622,n2623 );
   nor U2711 ( n2623,n1852,n1858 );
   not U2712 ( n1858,memory_reg_12__0_ );
   not U2713 ( n1852,n2624 );
   nor U2714 ( n2624,n2588,n2610 );
   nor U2715 ( n2622,n1842,n1848 );
   not U2716 ( n1848,memory_reg_13__0_ );
   not U2717 ( n1842,n2625 );
   nor U2718 ( n2625,n2590,n2610 );
   not U2719 ( n2610,n2626 );
   nor U2720 ( n2626,n2408,n2627 );
   not U2721 ( n2627,n2628 );
   nor U2722 ( n2628,address_reg_4_,address_reg_1_ );
   not U2723 ( n2619,n2629 );
   nor U2724 ( n2629,n2630,n2631 );
   nor U2725 ( n2631,n1832,n1838 );
   not U2726 ( n1838,memory_reg_14__0_ );
   not U2727 ( n1832,n2632 );
   nor U2728 ( n2632,n2588,n2616 );
   nor U2729 ( n2630,n1822,n1828 );
   not U2730 ( n1828,memory_reg_15__0_ );
   not U2731 ( n1822,n2633 );
   nor U2732 ( n2633,n2590,n2616 );
   not U2733 ( n2616,n2634 );
   nor U2734 ( n2634,n2408,n2635 );
   not U2735 ( n2635,n2636 );
   nor U2736 ( n2636,address_reg_4_,n2422 );
   not U2737 ( n2556,n2637 );
   nor U2738 ( n2637,n2638,n2639 );
   not U2739 ( n2639,n2640 );
   nor U2740 ( n2640,n2641,n2642 );
   not U2741 ( n2642,n2643 );
   nor U2742 ( n2643,n2644,n2645 );
   not U2743 ( n2645,n2646 );
   nor U2744 ( n2646,n2647,n2648 );
   nor U2745 ( n2648,n1812,n1818 );
   not U2746 ( n1818,memory_reg_16__0_ );
   not U2747 ( n1812,n2649 );
   nor U2748 ( n2649,n2571,n2650 );
   nor U2749 ( n2647,n1802,n1808 );
   not U2750 ( n1808,memory_reg_17__0_ );
   not U2751 ( n1802,n2651 );
   nor U2752 ( n2651,n2574,n2650 );
   not U2753 ( n2644,n2652 );
   nor U2754 ( n2652,n2653,n2654 );
   nor U2755 ( n2654,n1792,n1798 );
   not U2756 ( n1798,memory_reg_18__0_ );
   not U2757 ( n1792,n2655 );
   nor U2758 ( n2655,n2571,n2656 );
   nor U2759 ( n2653,n1782,n1788 );
   not U2760 ( n1788,memory_reg_19__0_ );
   not U2761 ( n1782,n2657 );
   nor U2762 ( n2657,n2574,n2656 );
   not U2763 ( n2641,n2658 );
   nor U2764 ( n2658,n2659,n2660 );
   not U2765 ( n2660,n2661 );
   nor U2766 ( n2661,n2662,n2663 );
   nor U2767 ( n2663,n1772,n1778 );
   not U2768 ( n1778,memory_reg_20__0_ );
   not U2769 ( n1772,n2664 );
   nor U2770 ( n2664,n2588,n2650 );
   nor U2771 ( n2662,n1762,n1768 );
   not U2772 ( n1768,memory_reg_21__0_ );
   not U2773 ( n1762,n2665 );
   nor U2774 ( n2665,n2590,n2650 );
   not U2775 ( n2650,n2666 );
   nor U2776 ( n2666,n2400,n2667 );
   not U2777 ( n2667,n2668 );
   nor U2778 ( n2668,address_reg_3_,address_reg_1_ );
   not U2779 ( n2659,n2669 );
   nor U2780 ( n2669,n2670,n2671 );
   nor U2781 ( n2671,n1752,n1758 );
   not U2782 ( n1758,memory_reg_22__0_ );
   not U2783 ( n1752,n2672 );
   nor U2784 ( n2672,n2588,n2656 );
   nor U2785 ( n2670,n1742,n1748 );
   not U2786 ( n1748,memory_reg_23__0_ );
   not U2787 ( n1742,n2673 );
   nor U2788 ( n2673,n2590,n2656 );
   not U2789 ( n2656,n2674 );
   nor U2790 ( n2674,n2400,n2675 );
   not U2791 ( n2675,n2676 );
   nor U2792 ( n2676,address_reg_3_,n2422 );
   not U2793 ( n2638,n2677 );
   nor U2794 ( n2677,n2678,n2679 );
   not U2795 ( n2679,n2680 );
   nor U2796 ( n2680,n2681,n2682 );
   not U2797 ( n2682,n2683 );
   nor U2798 ( n2683,n2684,n2685 );
   nor U2799 ( n2685,n1732,n1738 );
   not U2800 ( n1738,memory_reg_24__0_ );
   not U2801 ( n1732,n2686 );
   nor U2802 ( n2686,n2687,n2571 );
   nor U2803 ( n2684,n1722,n1728 );
   not U2804 ( n1728,memory_reg_25__0_ );
   not U2805 ( n1722,n2688 );
   nor U2806 ( n2688,n2687,n2574 );
   not U2807 ( n2681,n2689 );
   nor U2808 ( n2689,n2690,n2691 );
   nor U2809 ( n2691,n1712,n1718 );
   not U2810 ( n1718,memory_reg_26__0_ );
   not U2811 ( n1712,n2692 );
   nor U2812 ( n2692,n2693,n2571 );
   not U2813 ( n2571,n2694 );
   nor U2814 ( n2694,address_reg_2_,address_reg_0_ );
   nor U2815 ( n2690,n1702,n1708 );
   not U2816 ( n1708,memory_reg_27__0_ );
   not U2817 ( n1702,n2695 );
   nor U2818 ( n2695,n2693,n2574 );
   not U2819 ( n2574,n2696 );
   nor U2820 ( n2696,address_reg_2_,n2434 );
   not U2821 ( n2678,n2697 );
   nor U2822 ( n2697,n2698,n2699 );
   not U2823 ( n2699,n2700 );
   nor U2824 ( n2700,n2701,n2702 );
   nor U2825 ( n2702,n1692,n1698 );
   not U2826 ( n1698,memory_reg_28__0_ );
   not U2827 ( n1692,n2703 );
   nor U2828 ( n2703,n2588,n2687 );
   nor U2829 ( n2701,n1682,n1688 );
   not U2830 ( n1688,memory_reg_29__0_ );
   not U2831 ( n1682,n2704 );
   nor U2832 ( n2704,n2590,n2687 );
   not U2833 ( n2687,n2705 );
   nor U2834 ( n2705,n2400,n2706 );
   not U2835 ( n2706,n2707 );
   nor U2836 ( n2707,address_reg_1_,n2408 );
   not U2837 ( n2698,n2708 );
   nor U2838 ( n2708,n2709,n2710 );
   nor U2839 ( n2710,n1672,n1678 );
   not U2840 ( n1678,memory_reg_30__0_ );
   not U2841 ( n1672,n2711 );
   nor U2842 ( n2711,n2693,n2588 );
   not U2843 ( n2588,n2712 );
   nor U2844 ( n2712,address_reg_0_,n2415 );
   nor U2845 ( n2709,n1662,n1668 );
   not U2846 ( n1668,memory_reg_31__0_ );
   not U2847 ( n1662,n2713 );
   nor U2848 ( n2713,n2693,n2590 );
   not U2849 ( n2590,n2714 );
   nor U2850 ( n2714,n2434,n2415 );
   not U2851 ( n2415,address_reg_2_ );
   not U2852 ( n2434,address_reg_0_ );
   not U2853 ( n2693,n2715 );
   nor U2854 ( n2715,n2400,n2716 );
   not U2855 ( n2716,n2717 );
   nor U2856 ( n2717,n2422,n2408 );
   not U2857 ( n2408,address_reg_3_ );
   not U2858 ( n2422,address_reg_1_ );
   not U2859 ( n2400,address_reg_4_ );
   not U2860 ( u1388,n2718 );
   nor U2861 ( n2718,n2719,n2720 );
   not U2862 ( n2720,n2721 );
   nor U2863 ( n2721,n2722,n2723 );
   not U2864 ( n2723,n2724 );
   nor U2865 ( n2724,n2725,n2726 );
   nor U2866 ( n2725,n2727,n1658 );
   nor U2867 ( n2727,n2728,n2729 );
   nor U2868 ( n2729,data_out_reg_1_,n2730 );
   nor U2869 ( n2730,n2731,n2732 );
   not U2870 ( n2732,n2733 );
   nor U2871 ( n2731,data_out_reg_0_,n2734 );
   nor U2872 ( n2728,n1571,n2735 );
   not U2873 ( n2735,n2736 );
   nor U2874 ( n2736,n2737,n2738 );
   nor U2875 ( n2738,data_out_reg_0_,n2739 );
   nor U2876 ( n2739,n2733,n1651 );
   nor U2877 ( n2737,n2740,n1562 );
   nor U2878 ( n2740,n2741,n2742 );
   not U2879 ( n2742,n2743 );
   nor U2880 ( n2743,k_2_,n2733 );
   nor U2881 ( n2733,data_out_reg_1_,n2744 );
   nor U2882 ( n2744,n2745,n2746 );
   not U2883 ( n2746,n2747 );
   nor U2884 ( n2747,k_0_,n1562 );
   not U2885 ( n2722,n2748 );
   nor U2886 ( n2748,n2749,n2750 );
   nor U2887 ( n2750,n2751,n1478 );
   nor U2888 ( n2751,n2752,n2753 );
   not U2889 ( n2753,n2754 );
   nor U2890 ( n2754,n2755,n2192 );
   not U2891 ( n2192,n2756 );
   nor U2892 ( n2756,n2757,n2758 );
   nor U2893 ( n2758,n2137,n2759 );
   nor U2894 ( n2749,n2294,n2760 );
   nor U2895 ( n2760,n2761,n2762 );
   not U2896 ( n2762,n2763 );
   nor U2897 ( n2763,n2764,n1595 );
   nor U2898 ( n1595,n1512,n2055 );
   not U2899 ( n2055,n1507 );
   not U2900 ( n2761,n2765 );
   nor U2901 ( n2765,n2766,n2052 );
   not U2902 ( n2719,n2767 );
   nor U2903 ( n2767,n2768,n2769 );
   not U2904 ( n2769,n2770 );
   nor U2905 ( n2770,n2435,n2771 );
   nor U2906 ( n2435,n2338,n2070 );
   not U2907 ( n2070,n2772 );
   nor U2908 ( n2772,n1485,n1560 );
   nor U2909 ( n2768,n1582,n2773 );
   not U2910 ( n2773,n2774 );
   nor U2911 ( n2774,n1506,n1532 );
   not U2912 ( u1387,n2775 );
   nor U2913 ( n2775,n2776,n2777 );
   not U2914 ( n2777,n2778 );
   nor U2915 ( n2778,n2779,n2780 );
   not U2916 ( n2780,n2781 );
   nor U2917 ( n2781,n2726,n2782 );
   not U2918 ( n2782,n2783 );
   nor U2919 ( n2783,n2784,n2785 );
   nor U2920 ( n2785,n1501,n1560 );
   not U2921 ( n1560,n2043 );
   nor U2922 ( n2784,n2043,n1532 );
   nor U2923 ( n2043,n1506,n1514 );
   not U2924 ( n2726,n2786 );
   nor U2925 ( n2786,n2787,n2788 );
   not U2926 ( n2788,n2789 );
   nor U2927 ( n2789,n2790,n2791 );
   nor U2928 ( n2791,n2137,n2142 );
   nor U2929 ( n2790,n1532,n2193 );
   not U2930 ( n2193,n1581 );
   nor U2931 ( n1581,n1508,n1506 );
   not U2932 ( n2779,n2792 );
   nor U2933 ( n2792,n1534,n2793 );
   nor U2934 ( n2793,n1506,n2069 );
   not U2935 ( n2776,n2794 );
   nor U2936 ( n2794,n2795,n2796 );
   not U2937 ( n2796,n2797 );
   nor U2938 ( n2797,n1592,n2219 );
   nor U2939 ( n2219,n2798,n2799 );
   not U2940 ( n2799,n2800 );
   nor U2941 ( n2800,n2801,n1603 );
   not U2942 ( n2795,n2802 );
   nor U2943 ( n2802,n2803,n2052 );
   not U2944 ( u1386,n2804 );
   nor U2945 ( n2804,n2805,n2806 );
   not U2946 ( n2806,n2807 );
   nor U2947 ( n2807,n2808,n2809 );
   not U2948 ( n2809,n2810 );
   nor U2949 ( n2810,n2752,n2811 );
   not U2950 ( n2811,n2812 );
   nor U2951 ( n2812,n2813,n2814 );
   nor U2952 ( n2814,n1513,n2194 );
   not U2953 ( n2194,n2755 );
   nor U2954 ( n2755,n1582,n2338 );
   nor U2955 ( n2813,n1506,n1597 );
   not U2956 ( n2752,n2815 );
   nor U2957 ( n2815,n2079,n1529 );
   nor U2958 ( n2079,n1532,n1477 );
   not U2959 ( n2808,n2816 );
   nor U2960 ( n2816,n2378,n2787 );
   not U2961 ( n2787,n2817 );
   nor U2962 ( n2817,n2072,n2818 );
   nor U2963 ( n2818,n2819,n2294 );
   nor U2964 ( n2819,n1528,n2820 );
   not U2965 ( n2378,n2821 );
   nor U2966 ( n2821,n1592,n2822 );
   nor U2967 ( n2822,n2823,n2294 );
   nor U2968 ( n2823,n2766,n2764 );
   nor U2969 ( n1592,n1603,n2759 );
   not U2970 ( n2759,n2764 );
   nor U2971 ( n2764,n1513,n2824 );
   not U2972 ( n2824,n2320 );
   nor U2973 ( n2320,n1501,n1582 );
   not U2974 ( n2805,n2825 );
   nor U2975 ( n2825,n2826,n2827 );
   not U2976 ( n2827,n2828 );
   nor U2977 ( n2828,n1599,n2771 );
   nor U2978 ( n2771,n2375,n2359 );
   not U2979 ( n2359,n2829 );
   nor U2980 ( n2829,n2330,n1477 );
   not U2981 ( n2375,n2337 );
   nor U2982 ( n2337,n2058,n2331 );
   nor U2983 ( n1599,n1513,n2830 );
   not U2984 ( n2830,n1534 );
   nor U2985 ( n1534,n1514,n2069 );
   not U2986 ( n2069,n2087 );
   nor U2987 ( n2087,n1508,n1501 );
   not U2988 ( n2826,n2831 );
   nor U2989 ( n2831,n1489,n2052 );
   nor U2990 ( n2052,n1597,n2832 );
   not U2991 ( n2832,n1504 );
   nor U2992 ( n1504,n1582,n1477 );
   nor U2993 ( n1489,n2833,n1658 );
   not U2994 ( n1658,n2803 );
   nor U2995 ( n2833,n2834,n2835 );
   not U2996 ( n2835,n2836 );
   nor U2997 ( n2836,n2837,n2838 );
   nor U2998 ( n2838,n1562,n2734 );
   not U2999 ( n2734,k_0_ );
   nor U3000 ( n2837,k_0_,n2839 );
   not U3001 ( n2839,n2840 );
   nor U3002 ( n2840,data_out_reg_0_,n2745 );
   not U3003 ( n2745,k_1_ );
   not U3004 ( n2834,n2841 );
   nor U3005 ( n2841,n2842,n2843 );
   nor U3006 ( n2843,n1571,n2844 );
   nor U3007 ( n2844,n2845,n2846 );
   nor U3008 ( n2846,k_2_,n2847 );
   not U3009 ( n2847,n2848 );
   nor U3010 ( n2848,n1997,n2741 );
   not U3011 ( n2741,k_3_ );
   nor U3012 ( n1997,n1562,n1573 );
   not U3013 ( n1562,data_out_reg_0_ );
   nor U3014 ( n2845,n2010,n1651 );
   not U3015 ( n1651,k_2_ );
   nor U3016 ( n2010,data_out_reg_0_,n1573 );
   not U3017 ( n1571,n2849 );
   nor U3018 ( n2842,n2849,n1573 );
   not U3019 ( n1573,data_out_reg_1_ );
   nor U3020 ( n2849,k_1_,k_0_ );
   not U3021 ( u1385,n2850 );
   nor U3022 ( n2850,n2851,n2852 );
   not U3023 ( n2852,n2853 );
   nor U3024 ( n2853,n2854,n2855 );
   not U3025 ( n2855,n2856 );
   nor U3026 ( n2856,n2857,n2858 );
   nor U3027 ( n2858,n2294,n2385 );
   nor U3028 ( n2857,n1603,n2142 );
   not U3029 ( n2142,n2820 );
   nor U3030 ( n2820,n2331,n2859 );
   not U3031 ( n2859,n2860 );
   nor U3032 ( n2860,n1513,n1597 );
   not U3033 ( n2331,n2861 );
   nor U3034 ( n2861,n1508,n1514 );
   not U3035 ( n2854,n2862 );
   nor U3036 ( n2862,n2863,n2864 );
   nor U3037 ( n2864,n2865,n2357 );
   nor U3038 ( n2865,n2322,n2866 );
   not U3039 ( n2866,n2867 );
   nor U3040 ( n2867,n2081,n1511 );
   nor U3041 ( n2863,n2868,n2798 );
   nor U3042 ( n2868,n2801,n1478 );
   not U3043 ( n2851,n2869 );
   nor U3044 ( n2869,n2870,n2871 );
   not U3045 ( n2871,n2872 );
   nor U3046 ( n2872,n2803,n2072 );
   nor U3047 ( n2072,n1532,n2082 );
   nor U3048 ( n2803,n2294,n1515 );
   not U3049 ( n2870,n2873 );
   nor U3050 ( n2873,n2141,n2874 );
   not U3051 ( n2874,n2875 );
   nor U3052 ( n2875,n1529,n1507 );
   nor U3053 ( n1507,n1485,n1582 );
   not U3054 ( n1582,n1514 );
   nor U3055 ( n1529,n2082,n2338 );
   not U3056 ( n2338,n2322 );
   nor U3057 ( n2322,n2330,n2058 );
   nor U3058 ( n2141,n2798,n2876 );
   not U3059 ( n2876,n2877 );
   nor U3060 ( n2877,n2137,n1478 );
   not U3061 ( u1384,n2878 );
   nor U3062 ( n2878,n2879,n2880 );
   not U3063 ( n2880,n2881 );
   nor U3064 ( n2881,n1490,n2882 );
   nor U3065 ( n2882,n1524,n2385 );
   not U3066 ( n2385,n1528 );
   nor U3067 ( n1528,n1597,n2082 );
   not U3068 ( n1597,n1511 );
   nor U3069 ( n1511,n1512,n2280 );
   nor U3070 ( n1490,n1515,n1478 );
   not U3071 ( n1515,n2757 );
   nor U3072 ( n2757,n2357,n1532 );
   not U3073 ( n1532,n2042 );
   nor U3074 ( n2042,n2058,n2280 );
   not U3075 ( n2280,n2330 );
   not U3076 ( n2058,n1512 );
   not U3077 ( n2357,n2883 );
   nor U3078 ( n2883,n1506,n1485 );
   not U3079 ( n2879,n2884 );
   nor U3080 ( n2884,n2389,n1514 );
   nor U3081 ( n1514,start,n2885 );
   not U3082 ( n2885,gamma_reg_4_ );
   nor U3083 ( n2389,n2798,n2886 );
   not U3084 ( n2886,n2887 );
   nor U3085 ( n2887,n1605,n1603 );
   not U3086 ( n1603,n2888 );
   nor U3087 ( n2888,n1524,n2889 );
   not U3088 ( n2889,n2137 );
   nor U3089 ( n2137,n2890,n2891 );
   not U3090 ( n2891,n2892 );
   nor U3091 ( n2892,n2893,n2894 );
   xor U3092 ( n2894,n2096,n2151 );
   not U3093 ( n2096,scan_reg_3_ );
   xor U3094 ( n2893,n2111,n2173 );
   not U3095 ( n2111,scan_reg_2_ );
   not U3096 ( n2890,n2895 );
   nor U3097 ( n2895,n2896,n2897 );
   not U3098 ( n2897,n2898 );
   nor U3099 ( n2898,n2899,n2900 );
   xor U3100 ( n2900,n2119,n2183 );
   not U3101 ( n2119,scan_reg_1_ );
   xor U3102 ( n2899,n2099,n2154 );
   not U3103 ( n2099,scan_reg_4_ );
   xor U3104 ( n2896,n2120,n2182 );
   not U3105 ( n2120,scan_reg_0_ );
   not U3106 ( n1524,n2294 );
   nor U3107 ( n2294,n2901,n2902 );
   not U3108 ( n2902,n2903 );
   nor U3109 ( n2903,count_reg2_0_,n2904 );
   not U3110 ( n2904,n2905 );
   nor U3111 ( n2905,count_reg2_2_,count_reg2_1_ );
   not U3112 ( n2901,n2906 );
   nor U3113 ( n2906,count_reg2_3_,n2907 );
   not U3114 ( n2907,n2908 );
   nor U3115 ( n2908,count_reg2_5_,count_reg2_4_ );
   not U3116 ( n1605,n2801 );
   nor U3117 ( n2801,n2152,n2909 );
   not U3118 ( n2909,n2910 );
   nor U3119 ( n2910,n2154,n2151 );
   not U3120 ( n2151,max_reg_3_ );
   not U3121 ( n2154,max_reg_4_ );
   not U3122 ( n2152,n2165 );
   nor U3123 ( n2165,n2173,n2171 );
   not U3124 ( n2171,n2911 );
   nor U3125 ( n2911,n2183,n2182 );
   not U3126 ( n2182,max_reg_0_ );
   not U3127 ( n2183,max_reg_1_ );
   not U3128 ( n2173,max_reg_2_ );
   not U3129 ( n2798,n2766 );
   nor U3130 ( n2766,n1501,n2082 );
   not U3131 ( n2082,n1580 );
   nor U3132 ( n1580,n1485,n1477 );
   not U3133 ( n1513,n1506 );
   nor U3134 ( n1506,start,n2912 );
   not U3135 ( n2912,gamma_reg_2_ );
   not U3136 ( n1485,n1508 );
   nor U3137 ( n1508,start,n2913 );
   not U3138 ( n2913,gamma_reg_3_ );
   not U3139 ( n1501,n2081 );
   nor U3140 ( n2081,n2330,n1512 );
   nor U3141 ( n1512,start,gamma_reg_0_ );
   nor U3142 ( n2330,start,n2914 );
   not U3143 ( n2914,gamma_reg_1_ );
   not U3144 ( u1382,n2915 );
   nor U3145 ( n2915,n2916,n2917 );
   nor U3146 ( n2917,n2918,n2919 );
   not U3147 ( n2919,n2948 );
   nor U3148 ( n2948,counter_reg_0_,n2920 );
   nor U3149 ( n2916,counter_reg_1_,n2921 );
   not U3150 ( n2921,n2922 );
   nor U3151 ( n2922,n2923,n2920 );
   nor U3152 ( n2947,n2924,n2920 );
   not U3153 ( n2920,n2925 );
   nor U3154 ( n2925,n2926,n2927 );
   not U3155 ( n2927,n2928 );
   nor U3156 ( n2928,n2454,n1516 );
   not U3157 ( n1516,play_reg );
   nor U3158 ( n2454,n1574,n1583 );
   not U3159 ( n2926,n2453 );
   nor U3160 ( n2453,n2929,n2930 );
   nor U3161 ( n2930,n2931,n2932 );
   not U3162 ( n2932,n2933 );
   not U3163 ( n2931,counter_reg_2_ );
   nor U3164 ( n2929,n2934,n2935 );
   nor U3165 ( n2935,n2933,counter_reg_2_ );
   nor U3166 ( n2933,sound_reg_1_,n2936 );
   nor U3167 ( n2936,sound_reg_0_,n1583 );
   nor U3168 ( n2934,n2937,n2938 );
   nor U3169 ( n2938,n2939,n2918 );
   nor U3170 ( n2939,sound_reg_1_,n2940 );
   not U3171 ( n2940,n2941 );
   nor U3172 ( n2941,n2942,n2943 );
   nor U3173 ( n2943,n1583,n1564 );
   not U3174 ( n1564,sound_reg_0_ );
   not U3175 ( n1583,sound_reg_2_ );
   nor U3176 ( n2942,sound_reg_0_,n2923 );
   nor U3177 ( n2937,n2923,n2944 );
   not U3178 ( n2944,n2945 );
   nor U3179 ( n2945,sound_reg_0_,n1574 );
   not U3180 ( n1574,sound_reg_1_ );
   nor U3181 ( n2924,n2946,counter_reg_2_ );
   nor U3182 ( n2946,n2923,n2918 );
   not U3183 ( n2918,counter_reg_1_ );
   not U3184 ( n2923,counter_reg_0_ );
endmodule
