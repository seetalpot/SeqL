
module b20 ( si_31_, si_30_, si_29_, si_28_, si_27_, si_26_, si_25_, si_24_,         si_23_, si_22_, si_21_, si_20_, si_19_, si_18_, si_17_, si_16_, si_15_,         si_14_, si_13_, si_12_, si_11_, si_10_, si_9_, si_8_, si_7_, si_6_,         si_5_, si_4_, si_3_, si_2_, si_1_, si_0_, p1_ir_reg_0_, p1_ir_reg_1_,         p1_ir_reg_2_, p1_ir_reg_3_, p1_ir_reg_4_, p1_ir_reg_5_, p1_ir_reg_6_,         p1_ir_reg_7_, p1_ir_reg_8_, p1_ir_reg_9_, p1_ir_reg_10_, p1_ir_reg_11_,         p1_ir_reg_12_, p1_ir_reg_13_, p1_ir_reg_14_, p1_ir_reg_15_,         p1_ir_reg_16_, p1_ir_reg_17_, p1_ir_reg_18_, p1_ir_reg_19_,         p1_ir_reg_20_, p1_ir_reg_21_, p1_ir_reg_22_, p1_ir_reg_23_,         p1_ir_reg_24_, p1_ir_reg_25_, p1_ir_reg_26_, p1_ir_reg_27_,         p1_ir_reg_28_, p1_ir_reg_29_, p1_ir_reg_30_, p1_ir_reg_31_,         p1_d_reg_0_, p1_d_reg_1_, p1_d_reg_2_, p1_d_reg_3_, p1_d_reg_4_,         p1_d_reg_5_, p1_d_reg_6_, p1_d_reg_7_, p1_d_reg_8_, p1_d_reg_9_,         p1_d_reg_10_, p1_d_reg_11_, p1_d_reg_12_, p1_d_reg_13_, p1_d_reg_14_,         p1_d_reg_15_, p1_d_reg_16_, p1_d_reg_17_, p1_d_reg_18_, p1_d_reg_19_,         p1_d_reg_20_, p1_d_reg_21_, p1_d_reg_22_, p1_d_reg_23_, p1_d_reg_24_,         p1_d_reg_25_, p1_d_reg_26_, p1_d_reg_27_, p1_d_reg_28_, p1_d_reg_29_,         p1_d_reg_30_, p1_d_reg_31_, p1_reg0_reg_0_, p1_reg0_reg_1_,         p1_reg0_reg_2_, p1_reg0_reg_3_, p1_reg0_reg_4_, p1_reg0_reg_5_,         p1_reg0_reg_6_, p1_reg0_reg_7_, p1_reg0_reg_8_, p1_reg0_reg_9_,         p1_reg0_reg_10_, p1_reg0_reg_11_, p1_reg0_reg_12_, p1_reg0_reg_13_,         p1_reg0_reg_14_, p1_reg0_reg_15_, p1_reg0_reg_16_, p1_reg0_reg_17_,         p1_reg0_reg_18_, p1_reg0_reg_19_, p1_reg0_reg_20_, p1_reg0_reg_21_,         p1_reg0_reg_22_, p1_reg0_reg_23_, p1_reg0_reg_24_, p1_reg0_reg_25_,         p1_reg0_reg_26_, p1_reg0_reg_27_, p1_reg0_reg_28_, p1_reg0_reg_29_,         p1_reg0_reg_30_, p1_reg0_reg_31_, p1_reg1_reg_0_, p1_reg1_reg_1_,         p1_reg1_reg_2_, p1_reg1_reg_3_, p1_reg1_reg_4_, p1_reg1_reg_5_,         p1_reg1_reg_6_, p1_reg1_reg_7_, p1_reg1_reg_8_, p1_reg1_reg_9_,         p1_reg1_reg_10_, p1_reg1_reg_11_, p1_reg1_reg_12_, p1_reg1_reg_13_,         p1_reg1_reg_14_, p1_reg1_reg_15_, p1_reg1_reg_16_, p1_reg1_reg_17_,         p1_reg1_reg_18_, p1_reg1_reg_19_, p1_reg1_reg_20_, p1_reg1_reg_21_,         p1_reg1_reg_22_, p1_reg1_reg_23_, p1_reg1_reg_24_, p1_reg1_reg_25_,         p1_reg1_reg_26_, p1_reg1_reg_27_, p1_reg1_reg_28_, p1_reg1_reg_29_,         p1_reg1_reg_30_, p1_reg1_reg_31_, p1_reg2_reg_0_, p1_reg2_reg_1_,         p1_reg2_reg_2_, p1_reg2_reg_3_, p1_reg2_reg_4_, p1_reg2_reg_5_,         p1_reg2_reg_6_, p1_reg2_reg_7_, p1_reg2_reg_8_, p1_reg2_reg_9_,         p1_reg2_reg_10_, p1_reg2_reg_11_, p1_reg2_reg_12_, p1_reg2_reg_13_,         p1_reg2_reg_14_, p1_reg2_reg_15_, p1_reg2_reg_16_, p1_reg2_reg_17_,         p1_reg2_reg_18_, p1_reg2_reg_19_, p1_reg2_reg_20_, p1_reg2_reg_21_,         p1_reg2_reg_22_, p1_reg2_reg_23_, p1_reg2_reg_24_, p1_reg2_reg_25_,         p1_reg2_reg_26_, p1_reg2_reg_27_, p1_reg2_reg_28_, p1_reg2_reg_29_,         p1_reg2_reg_30_, p1_reg2_reg_31_, p1_addr_reg_19_, p1_addr_reg_18_,         p1_addr_reg_17_, p1_addr_reg_16_, p1_addr_reg_15_, p1_addr_reg_14_,         p1_addr_reg_13_, p1_addr_reg_12_, p1_addr_reg_11_, p1_addr_reg_10_,         p1_addr_reg_9_, p1_addr_reg_8_, p1_addr_reg_7_, p1_addr_reg_6_,         p1_addr_reg_5_, p1_addr_reg_4_, p1_addr_reg_3_, p1_addr_reg_2_,         p1_addr_reg_1_, p1_addr_reg_0_, p1_datao_reg_0_, p1_datao_reg_1_,         p1_datao_reg_2_, p1_datao_reg_3_, p1_datao_reg_4_, p1_datao_reg_5_,         p1_datao_reg_6_, p1_datao_reg_7_, p1_datao_reg_8_, p1_datao_reg_9_,         p1_datao_reg_10_, p1_datao_reg_11_, p1_datao_reg_12_, p1_datao_reg_13_,         p1_datao_reg_14_, p1_datao_reg_15_, p1_datao_reg_16_, p1_datao_reg_17_,         p1_datao_reg_18_, p1_datao_reg_19_, p1_datao_reg_20_, p1_datao_reg_21_,         p1_datao_reg_22_, p1_datao_reg_23_, p1_datao_reg_24_, p1_datao_reg_25_,         p1_datao_reg_26_, p1_datao_reg_27_, p1_datao_reg_28_, p1_datao_reg_29_,         p1_datao_reg_30_, p1_datao_reg_31_, p1_b_reg, p1_reg3_reg_15_,         p1_reg3_reg_26_, p1_reg3_reg_6_, p1_reg3_reg_18_, p1_reg3_reg_2_,         p1_reg3_reg_11_, p1_reg3_reg_22_, p1_reg3_reg_13_, p1_reg3_reg_20_,         p1_reg3_reg_0_, p1_reg3_reg_9_, p1_reg3_reg_4_, p1_reg3_reg_24_,         p1_reg3_reg_17_, p1_reg3_reg_5_, p1_reg3_reg_16_, p1_reg3_reg_25_,         p1_reg3_reg_12_, p1_reg3_reg_21_, p1_reg3_reg_1_, p1_reg3_reg_8_,         p1_reg3_reg_28_, p1_reg3_reg_19_, p1_reg3_reg_3_, p1_reg3_reg_10_,         p1_reg3_reg_23_, p1_reg3_reg_14_, p1_reg3_reg_27_, p1_reg3_reg_7_,         p1_state_reg, p1_rd_reg, p1_wr_reg, p2_ir_reg_0_, p2_ir_reg_1_,         p2_ir_reg_2_, p2_ir_reg_3_, p2_ir_reg_4_, p2_ir_reg_5_, p2_ir_reg_6_,         p2_ir_reg_7_, p2_ir_reg_8_, p2_ir_reg_9_, p2_ir_reg_10_, p2_ir_reg_11_,         p2_ir_reg_12_, p2_ir_reg_13_, p2_ir_reg_14_, p2_ir_reg_15_,         p2_ir_reg_16_, p2_ir_reg_17_, p2_ir_reg_18_, p2_ir_reg_19_,         p2_ir_reg_20_, p2_ir_reg_21_, p2_ir_reg_22_, p2_ir_reg_23_,         p2_ir_reg_24_, p2_ir_reg_25_, p2_ir_reg_26_, p2_ir_reg_27_,         p2_ir_reg_28_, p2_ir_reg_29_, p2_ir_reg_30_, p2_ir_reg_31_,         p2_d_reg_0_, p2_d_reg_1_, p2_d_reg_2_, p2_d_reg_3_, p2_d_reg_4_,         p2_d_reg_5_, p2_d_reg_6_, p2_d_reg_7_, p2_d_reg_8_, p2_d_reg_9_,         p2_d_reg_10_, p2_d_reg_11_, p2_d_reg_12_, p2_d_reg_13_, p2_d_reg_14_,         p2_d_reg_15_, p2_d_reg_16_, p2_d_reg_17_, p2_d_reg_18_, p2_d_reg_19_,         p2_d_reg_20_, p2_d_reg_21_, p2_d_reg_22_, p2_d_reg_23_, p2_d_reg_24_,         p2_d_reg_25_, p2_d_reg_26_, p2_d_reg_27_, p2_d_reg_28_, p2_d_reg_29_,         p2_d_reg_30_, p2_d_reg_31_, p2_reg0_reg_0_, p2_reg0_reg_1_,         p2_reg0_reg_2_, p2_reg0_reg_3_, p2_reg0_reg_4_, p2_reg0_reg_5_,         p2_reg0_reg_6_, p2_reg0_reg_7_, p2_reg0_reg_8_, p2_reg0_reg_9_,         p2_reg0_reg_10_, p2_reg0_reg_11_, p2_reg0_reg_12_, p2_reg0_reg_13_,         p2_reg0_reg_14_, p2_reg0_reg_15_, p2_reg0_reg_16_, p2_reg0_reg_17_,         p2_reg0_reg_18_, p2_reg0_reg_19_, p2_reg0_reg_20_, p2_reg0_reg_21_,         p2_reg0_reg_22_, p2_reg0_reg_23_, p2_reg0_reg_24_, p2_reg0_reg_25_,         p2_reg0_reg_26_, p2_reg0_reg_27_, p2_reg0_reg_28_, p2_reg0_reg_29_,         p2_reg0_reg_30_, p2_reg0_reg_31_, p2_reg1_reg_0_, p2_reg1_reg_1_,         p2_reg1_reg_2_, p2_reg1_reg_3_, p2_reg1_reg_4_, p2_reg1_reg_5_,         p2_reg1_reg_6_, p2_reg1_reg_7_, p2_reg1_reg_8_, p2_reg1_reg_9_,         p2_reg1_reg_10_, p2_reg1_reg_11_, p2_reg1_reg_12_, p2_reg1_reg_13_,         p2_reg1_reg_14_, p2_reg1_reg_15_, p2_reg1_reg_16_, p2_reg1_reg_17_,         p2_reg1_reg_18_, p2_reg1_reg_19_, p2_reg1_reg_20_, p2_reg1_reg_21_,         p2_reg1_reg_22_, p2_reg1_reg_23_, p2_reg1_reg_24_, p2_reg1_reg_25_,         p2_reg1_reg_26_, p2_reg1_reg_27_, p2_reg1_reg_28_, p2_reg1_reg_29_,         p2_reg1_reg_30_, p2_reg1_reg_31_, p2_reg2_reg_0_, p2_reg2_reg_1_,         p2_reg2_reg_2_, p2_reg2_reg_3_, p2_reg2_reg_4_, p2_reg2_reg_5_,         p2_reg2_reg_6_, p2_reg2_reg_7_, p2_reg2_reg_8_, p2_reg2_reg_9_,         p2_reg2_reg_10_, p2_reg2_reg_11_, p2_reg2_reg_12_, p2_reg2_reg_13_,         p2_reg2_reg_14_, p2_reg2_reg_15_, p2_reg2_reg_16_, p2_reg2_reg_17_,         p2_reg2_reg_18_, p2_reg2_reg_19_, p2_reg2_reg_20_, p2_reg2_reg_21_,         p2_reg2_reg_22_, p2_reg2_reg_23_, p2_reg2_reg_24_, p2_reg2_reg_25_,         p2_reg2_reg_26_, p2_reg2_reg_27_, p2_reg2_reg_28_, p2_reg2_reg_29_,         p2_reg2_reg_30_, p2_reg2_reg_31_, p2_addr_reg_19_, p2_addr_reg_18_,         p2_addr_reg_17_, p2_addr_reg_16_, p2_addr_reg_15_, p2_addr_reg_14_,         p2_addr_reg_13_, p2_addr_reg_12_, p2_addr_reg_11_, p2_addr_reg_10_,         p2_addr_reg_9_, p2_addr_reg_8_, p2_addr_reg_7_, p2_addr_reg_6_,         p2_addr_reg_5_, p2_addr_reg_4_, p2_addr_reg_3_, p2_addr_reg_2_,         p2_addr_reg_1_, p2_addr_reg_0_, p2_datao_reg_0_, p2_datao_reg_1_,         p2_datao_reg_2_, p2_datao_reg_3_, p2_datao_reg_4_, p2_datao_reg_5_,         p2_datao_reg_6_, p2_datao_reg_7_, p2_datao_reg_8_, p2_datao_reg_9_,         p2_datao_reg_10_, p2_datao_reg_11_, p2_datao_reg_12_, p2_datao_reg_13_,         p2_datao_reg_14_, p2_datao_reg_15_, p2_datao_reg_16_, p2_datao_reg_17_,         p2_datao_reg_18_, p2_datao_reg_19_, p2_datao_reg_20_, p2_datao_reg_21_,         p2_datao_reg_22_, p2_datao_reg_23_, p2_datao_reg_24_, p2_datao_reg_25_,         p2_datao_reg_26_, p2_datao_reg_27_, p2_datao_reg_28_, p2_datao_reg_29_,         p2_datao_reg_30_, p2_datao_reg_31_, p2_b_reg, p2_reg3_reg_15_,         p2_reg3_reg_26_, p2_reg3_reg_6_, p2_reg3_reg_18_, p2_reg3_reg_2_,         p2_reg3_reg_11_, p2_reg3_reg_22_, p2_reg3_reg_13_, p2_reg3_reg_20_,         p2_reg3_reg_0_, p2_reg3_reg_9_, p2_reg3_reg_4_, p2_reg3_reg_24_,         p2_reg3_reg_17_, p2_reg3_reg_5_, p2_reg3_reg_16_, p2_reg3_reg_25_,         p2_reg3_reg_12_, p2_reg3_reg_21_, p2_reg3_reg_1_, p2_reg3_reg_8_,         p2_reg3_reg_28_, p2_reg3_reg_19_, p2_reg3_reg_3_, p2_reg3_reg_10_,         p2_reg3_reg_23_, p2_reg3_reg_14_, p2_reg3_reg_27_, p2_reg3_reg_7_,         p2_state_reg, p2_rd_reg, p2_wr_reg, add_1068_u4, add_1068_u55,         add_1068_u56, add_1068_u57, add_1068_u58, add_1068_u59, add_1068_u60,         add_1068_u61, add_1068_u62, add_1068_u63, add_1068_u47, add_1068_u48,         add_1068_u49, add_1068_u50, add_1068_u51, add_1068_u52, add_1068_u53,         add_1068_u54, add_1068_u5, add_1068_u46, u126, u123, p1_u3355,         p1_u3354, p1_u3353, p1_u3352, p1_u3351, p1_u3350, p1_u3349, p1_u3348,         p1_u3347, p1_u3346, p1_u3345, p1_u3344, p1_u3343, p1_u3342, p1_u3341,         p1_u3340, p1_u3339, p1_u3338, p1_u3337, p1_u3336, p1_u3335, p1_u3334,         p1_u3333, p1_u3332, p1_u3331, p1_u3330, p1_u3329, p1_u3328, p1_u3327,         p1_u3326, p1_u3325, p1_u3324, p1_u3439, p1_u3440, p1_u3323, p1_u3322,         p1_u3321, p1_u3320, p1_u3319, p1_u3318, p1_u3317, p1_u3316, p1_u3315,         p1_u3314, p1_u3313, p1_u3312, p1_u3311, p1_u3310, p1_u3309, p1_u3308,         p1_u3307, p1_u3306, p1_u3305, p1_u3304, p1_u3303, p1_u3302, p1_u3301,         p1_u3300, p1_u3299, p1_u3298, p1_u3297, p1_u3296, p1_u3295, p1_u3294,         p1_u3453, p1_u3456, p1_u3459, p1_u3462, p1_u3465, p1_u3468, p1_u3471,         p1_u3474, p1_u3477, p1_u3480, p1_u3483, p1_u3486, p1_u3489, p1_u3492,         p1_u3495, p1_u3498, p1_u3501, p1_u3504, p1_u3507, p1_u3509, p1_u3510,         p1_u3511, p1_u3512, p1_u3513, p1_u3514, p1_u3515, p1_u3516, p1_u3517,         p1_u3518, p1_u3519, p1_u3520, p1_u3521, p1_u3522, p1_u3523, p1_u3524,         p1_u3525, p1_u3526, p1_u3527, p1_u3528, p1_u3529, p1_u3530, p1_u3531,         p1_u3532, p1_u3533, p1_u3534, p1_u3535, p1_u3536, p1_u3537, p1_u3538,         p1_u3539, p1_u3540, p1_u3541, p1_u3542, p1_u3543, p1_u3544, p1_u3545,         p1_u3546, p1_u3547, p1_u3548, p1_u3549, p1_u3550, p1_u3551, p1_u3552,         p1_u3553, p1_u3293, p1_u3292, p1_u3291, p1_u3290, p1_u3289, p1_u3288,         p1_u3287, p1_u3286, p1_u3285, p1_u3284, p1_u3283, p1_u3282, p1_u3281,         p1_u3280, p1_u3279, p1_u3278, p1_u3277, p1_u3276, p1_u3275, p1_u3274,         p1_u3273, p1_u3272, p1_u3271, p1_u3270, p1_u3269, p1_u3268, p1_u3267,         p1_u3266, p1_u3265, p1_u3356, p1_u3264, p1_u3263, p1_u3262, p1_u3261,         p1_u3260, p1_u3259, p1_u3258, p1_u3257, p1_u3256, p1_u3255, p1_u3254,         p1_u3253, p1_u3252, p1_u3251, p1_u3250, p1_u3249, p1_u3248, p1_u3247,         p1_u3246, p1_u3245, p1_u3244, p1_u3243, p1_u3554, p1_u3555, p1_u3556,         p1_u3557, p1_u3558, p1_u3559, p1_u3560, p1_u3561, p1_u3562, p1_u3563,         p1_u3564, p1_u3565, p1_u3566, p1_u3567, p1_u3568, p1_u3569, p1_u3570,         p1_u3571, p1_u3572, p1_u3573, p1_u3574, p1_u3575, p1_u3576, p1_u3577,         p1_u3578, p1_u3579, p1_u3580, p1_u3581, p1_u3582, p1_u3583, p1_u3584,         p1_u3585, p1_u3242, p1_u3241, p1_u3240, p1_u3239, p1_u3238, p1_u3237,         p1_u3236, p1_u3235, p1_u3234, p1_u3233, p1_u3232, p1_u3231, p1_u3230,         p1_u3229, p1_u3228, p1_u3227, p1_u3226, p1_u3225, p1_u3224, p1_u3223,         p1_u3222, p1_u3221, p1_u3220, p1_u3219, p1_u3218, p1_u3217, p1_u3216,         p1_u3215, p1_u3214, p1_u3213, p1_u3086, p1_u3085, p1_u3973, p2_u3295,         p2_u3294, p2_u3293, p2_u3292, p2_u3291, p2_u3290, p2_u3289, p2_u3288,         p2_u3287, p2_u3286, p2_u3285, p2_u3284, p2_u3283, p2_u3282, p2_u3281,         p2_u3280, p2_u3279, p2_u3278, p2_u3277, p2_u3276, p2_u3275, p2_u3274,         p2_u3273, p2_u3272, p2_u3271, p2_u3270, p2_u3269, p2_u3268, p2_u3267,         p2_u3266, p2_u3265, p2_u3264, p2_u3376, p2_u3377, p2_u3263, p2_u3262,         p2_u3261, p2_u3260, p2_u3259, p2_u3258, p2_u3257, p2_u3256, p2_u3255,         p2_u3254, p2_u3253, p2_u3252, p2_u3251, p2_u3250, p2_u3249, p2_u3248,         p2_u3247, p2_u3246, p2_u3245, p2_u3244, p2_u3243, p2_u3242, p2_u3241,         p2_u3240, p2_u3239, p2_u3238, p2_u3237, p2_u3236, p2_u3235, p2_u3234,         p2_u3390, p2_u3393, p2_u3396, p2_u3399, p2_u3402, p2_u3405, p2_u3408,         p2_u3411, p2_u3414, p2_u3417, p2_u3420, p2_u3423, p2_u3426, p2_u3429,         p2_u3432, p2_u3435, p2_u3438, p2_u3441, p2_u3444, p2_u3446, p2_u3447,         p2_u3448, p2_u3449, p2_u3450, p2_u3451, p2_u3452, p2_u3453, p2_u3454,         p2_u3455, p2_u3456, p2_u3457, p2_u3458, p2_u3459, p2_u3460, p2_u3461,         p2_u3462, p2_u3463, p2_u3464, p2_u3465, p2_u3466, p2_u3467, p2_u3468,         p2_u3469, p2_u3470, p2_u3471, p2_u3472, p2_u3473, p2_u3474, p2_u3475,         p2_u3476, p2_u3477, p2_u3478, p2_u3479, p2_u3480, p2_u3481, p2_u3482,         p2_u3483, p2_u3484, p2_u3485, p2_u3486, p2_u3487, p2_u3488, p2_u3489,         p2_u3490, p2_u3233, p2_u3232, p2_u3231, p2_u3230, p2_u3229, p2_u3228,         p2_u3227, p2_u3226, p2_u3225, p2_u3224, p2_u3223, p2_u3222, p2_u3221,         p2_u3220, p2_u3219, p2_u3218, p2_u3217, p2_u3216, p2_u3215, p2_u3214,         p2_u3213, p2_u3212, p2_u3211, p2_u3210, p2_u3209, p2_u3208, p2_u3207,         p2_u3206, p2_u3205, p2_u3204, p2_u3203, p2_u3202, p2_u3201, p2_u3200,         p2_u3199, p2_u3198, p2_u3197, p2_u3196, p2_u3195, p2_u3194, p2_u3193,         p2_u3192, p2_u3191, p2_u3190, p2_u3189, p2_u3188, p2_u3187, p2_u3186,         p2_u3185, p2_u3184, p2_u3183, p2_u3182, p2_u3491, p2_u3492, p2_u3493,         p2_u3494, p2_u3495, p2_u3496, p2_u3497, p2_u3498, p2_u3499, p2_u3500,         p2_u3501, p2_u3502, p2_u3503, p2_u3504, p2_u3505, p2_u3506, p2_u3507,         p2_u3508, p2_u3509, p2_u3510, p2_u3511, p2_u3512, p2_u3513, p2_u3514,         p2_u3515, p2_u3516, p2_u3517, p2_u3518, p2_u3519, p2_u3520, p2_u3521,         p2_u3522, p2_u3296, p2_u3181, p2_u3180, p2_u3179, p2_u3178, p2_u3177,         p2_u3176, p2_u3175, p2_u3174, p2_u3173, p2_u3172, p2_u3171, p2_u3170,         p2_u3169, p2_u3168, p2_u3167, p2_u3166, p2_u3165, p2_u3164, p2_u3163,         p2_u3162, p2_u3161, p2_u3160, p2_u3159, p2_u3158, p2_u3157, p2_u3156,         p2_u3155, p2_u3154, p2_u3153, p2_u3151, p2_u3150, p2_u3893 );
input si_31_, si_30_, si_29_, si_28_, si_27_, si_26_, si_25_, si_24_, si_23_,         si_22_, si_21_, si_20_, si_19_, si_18_, si_17_, si_16_, si_15_,         si_14_, si_13_, si_12_, si_11_, si_10_, si_9_, si_8_, si_7_, si_6_,         si_5_, si_4_, si_3_, si_2_, si_1_, si_0_, p1_ir_reg_0_, p1_ir_reg_1_,         p1_ir_reg_2_, p1_ir_reg_3_, p1_ir_reg_4_, p1_ir_reg_5_, p1_ir_reg_6_,         p1_ir_reg_7_, p1_ir_reg_8_, p1_ir_reg_9_, p1_ir_reg_10_,         p1_ir_reg_11_, p1_ir_reg_12_, p1_ir_reg_13_, p1_ir_reg_14_,         p1_ir_reg_15_, p1_ir_reg_16_, p1_ir_reg_17_, p1_ir_reg_18_,         p1_ir_reg_19_, p1_ir_reg_20_, p1_ir_reg_21_, p1_ir_reg_22_,         p1_ir_reg_23_, p1_ir_reg_24_, p1_ir_reg_25_, p1_ir_reg_26_,         p1_ir_reg_27_, p1_ir_reg_28_, p1_ir_reg_29_, p1_ir_reg_30_,         p1_ir_reg_31_, p1_d_reg_0_, p1_d_reg_1_, p1_d_reg_2_, p1_d_reg_3_,         p1_d_reg_4_, p1_d_reg_5_, p1_d_reg_6_, p1_d_reg_7_, p1_d_reg_8_,         p1_d_reg_9_, p1_d_reg_10_, p1_d_reg_11_, p1_d_reg_12_, p1_d_reg_13_,         p1_d_reg_14_, p1_d_reg_15_, p1_d_reg_16_, p1_d_reg_17_, p1_d_reg_18_,         p1_d_reg_19_, p1_d_reg_20_, p1_d_reg_21_, p1_d_reg_22_, p1_d_reg_23_,         p1_d_reg_24_, p1_d_reg_25_, p1_d_reg_26_, p1_d_reg_27_, p1_d_reg_28_,         p1_d_reg_29_, p1_d_reg_30_, p1_d_reg_31_, p1_reg0_reg_0_,         p1_reg0_reg_1_, p1_reg0_reg_2_, p1_reg0_reg_3_, p1_reg0_reg_4_,         p1_reg0_reg_5_, p1_reg0_reg_6_, p1_reg0_reg_7_, p1_reg0_reg_8_,         p1_reg0_reg_9_, p1_reg0_reg_10_, p1_reg0_reg_11_, p1_reg0_reg_12_,         p1_reg0_reg_13_, p1_reg0_reg_14_, p1_reg0_reg_15_, p1_reg0_reg_16_,         p1_reg0_reg_17_, p1_reg0_reg_18_, p1_reg0_reg_19_, p1_reg0_reg_20_,         p1_reg0_reg_21_, p1_reg0_reg_22_, p1_reg0_reg_23_, p1_reg0_reg_24_,         p1_reg0_reg_25_, p1_reg0_reg_26_, p1_reg0_reg_27_, p1_reg0_reg_28_,         p1_reg0_reg_29_, p1_reg0_reg_30_, p1_reg0_reg_31_, p1_reg1_reg_0_,         p1_reg1_reg_1_, p1_reg1_reg_2_, p1_reg1_reg_3_, p1_reg1_reg_4_,         p1_reg1_reg_5_, p1_reg1_reg_6_, p1_reg1_reg_7_, p1_reg1_reg_8_,         p1_reg1_reg_9_, p1_reg1_reg_10_, p1_reg1_reg_11_, p1_reg1_reg_12_,         p1_reg1_reg_13_, p1_reg1_reg_14_, p1_reg1_reg_15_, p1_reg1_reg_16_,         p1_reg1_reg_17_, p1_reg1_reg_18_, p1_reg1_reg_19_, p1_reg1_reg_20_,         p1_reg1_reg_21_, p1_reg1_reg_22_, p1_reg1_reg_23_, p1_reg1_reg_24_,         p1_reg1_reg_25_, p1_reg1_reg_26_, p1_reg1_reg_27_, p1_reg1_reg_28_,         p1_reg1_reg_29_, p1_reg1_reg_30_, p1_reg1_reg_31_, p1_reg2_reg_0_,         p1_reg2_reg_1_, p1_reg2_reg_2_, p1_reg2_reg_3_, p1_reg2_reg_4_,         p1_reg2_reg_5_, p1_reg2_reg_6_, p1_reg2_reg_7_, p1_reg2_reg_8_,         p1_reg2_reg_9_, p1_reg2_reg_10_, p1_reg2_reg_11_, p1_reg2_reg_12_,         p1_reg2_reg_13_, p1_reg2_reg_14_, p1_reg2_reg_15_, p1_reg2_reg_16_,         p1_reg2_reg_17_, p1_reg2_reg_18_, p1_reg2_reg_19_, p1_reg2_reg_20_,         p1_reg2_reg_21_, p1_reg2_reg_22_, p1_reg2_reg_23_, p1_reg2_reg_24_,         p1_reg2_reg_25_, p1_reg2_reg_26_, p1_reg2_reg_27_, p1_reg2_reg_28_,         p1_reg2_reg_29_, p1_reg2_reg_30_, p1_reg2_reg_31_, p1_addr_reg_19_,         p1_addr_reg_18_, p1_addr_reg_17_, p1_addr_reg_16_, p1_addr_reg_15_,         p1_addr_reg_14_, p1_addr_reg_13_, p1_addr_reg_12_, p1_addr_reg_11_,         p1_addr_reg_10_, p1_addr_reg_9_, p1_addr_reg_8_, p1_addr_reg_7_,         p1_addr_reg_6_, p1_addr_reg_5_, p1_addr_reg_4_, p1_addr_reg_3_,         p1_addr_reg_2_, p1_addr_reg_1_, p1_addr_reg_0_, p1_datao_reg_0_,         p1_datao_reg_1_, p1_datao_reg_2_, p1_datao_reg_3_, p1_datao_reg_4_,         p1_datao_reg_5_, p1_datao_reg_6_, p1_datao_reg_7_, p1_datao_reg_8_,         p1_datao_reg_9_, p1_datao_reg_10_, p1_datao_reg_11_, p1_datao_reg_12_,         p1_datao_reg_13_, p1_datao_reg_14_, p1_datao_reg_15_,         p1_datao_reg_16_, p1_datao_reg_17_, p1_datao_reg_18_,         p1_datao_reg_19_, p1_datao_reg_20_, p1_datao_reg_21_,         p1_datao_reg_22_, p1_datao_reg_23_, p1_datao_reg_24_,         p1_datao_reg_25_, p1_datao_reg_26_, p1_datao_reg_27_,         p1_datao_reg_28_, p1_datao_reg_29_, p1_datao_reg_30_,         p1_datao_reg_31_, p1_b_reg, p1_reg3_reg_15_, p1_reg3_reg_26_,         p1_reg3_reg_6_, p1_reg3_reg_18_, p1_reg3_reg_2_, p1_reg3_reg_11_,         p1_reg3_reg_22_, p1_reg3_reg_13_, p1_reg3_reg_20_, p1_reg3_reg_0_,         p1_reg3_reg_9_, p1_reg3_reg_4_, p1_reg3_reg_24_, p1_reg3_reg_17_,         p1_reg3_reg_5_, p1_reg3_reg_16_, p1_reg3_reg_25_, p1_reg3_reg_12_,         p1_reg3_reg_21_, p1_reg3_reg_1_, p1_reg3_reg_8_, p1_reg3_reg_28_,         p1_reg3_reg_19_, p1_reg3_reg_3_, p1_reg3_reg_10_, p1_reg3_reg_23_,         p1_reg3_reg_14_, p1_reg3_reg_27_, p1_reg3_reg_7_, p1_state_reg,         p1_rd_reg, p1_wr_reg, p2_ir_reg_0_, p2_ir_reg_1_, p2_ir_reg_2_,         p2_ir_reg_3_, p2_ir_reg_4_, p2_ir_reg_5_, p2_ir_reg_6_, p2_ir_reg_7_,         p2_ir_reg_8_, p2_ir_reg_9_, p2_ir_reg_10_, p2_ir_reg_11_,         p2_ir_reg_12_, p2_ir_reg_13_, p2_ir_reg_14_, p2_ir_reg_15_,         p2_ir_reg_16_, p2_ir_reg_17_, p2_ir_reg_18_, p2_ir_reg_19_,         p2_ir_reg_20_, p2_ir_reg_21_, p2_ir_reg_22_, p2_ir_reg_23_,         p2_ir_reg_24_, p2_ir_reg_25_, p2_ir_reg_26_, p2_ir_reg_27_,         p2_ir_reg_28_, p2_ir_reg_29_, p2_ir_reg_30_, p2_ir_reg_31_,         p2_d_reg_0_, p2_d_reg_1_, p2_d_reg_2_, p2_d_reg_3_, p2_d_reg_4_,         p2_d_reg_5_, p2_d_reg_6_, p2_d_reg_7_, p2_d_reg_8_, p2_d_reg_9_,         p2_d_reg_10_, p2_d_reg_11_, p2_d_reg_12_, p2_d_reg_13_, p2_d_reg_14_,         p2_d_reg_15_, p2_d_reg_16_, p2_d_reg_17_, p2_d_reg_18_, p2_d_reg_19_,         p2_d_reg_20_, p2_d_reg_21_, p2_d_reg_22_, p2_d_reg_23_, p2_d_reg_24_,         p2_d_reg_25_, p2_d_reg_26_, p2_d_reg_27_, p2_d_reg_28_, p2_d_reg_29_,         p2_d_reg_30_, p2_d_reg_31_, p2_reg0_reg_0_, p2_reg0_reg_1_,         p2_reg0_reg_2_, p2_reg0_reg_3_, p2_reg0_reg_4_, p2_reg0_reg_5_,         p2_reg0_reg_6_, p2_reg0_reg_7_, p2_reg0_reg_8_, p2_reg0_reg_9_,         p2_reg0_reg_10_, p2_reg0_reg_11_, p2_reg0_reg_12_, p2_reg0_reg_13_,         p2_reg0_reg_14_, p2_reg0_reg_15_, p2_reg0_reg_16_, p2_reg0_reg_17_,         p2_reg0_reg_18_, p2_reg0_reg_19_, p2_reg0_reg_20_, p2_reg0_reg_21_,         p2_reg0_reg_22_, p2_reg0_reg_23_, p2_reg0_reg_24_, p2_reg0_reg_25_,         p2_reg0_reg_26_, p2_reg0_reg_27_, p2_reg0_reg_28_, p2_reg0_reg_29_,         p2_reg0_reg_30_, p2_reg0_reg_31_, p2_reg1_reg_0_, p2_reg1_reg_1_,         p2_reg1_reg_2_, p2_reg1_reg_3_, p2_reg1_reg_4_, p2_reg1_reg_5_,         p2_reg1_reg_6_, p2_reg1_reg_7_, p2_reg1_reg_8_, p2_reg1_reg_9_,         p2_reg1_reg_10_, p2_reg1_reg_11_, p2_reg1_reg_12_, p2_reg1_reg_13_,         p2_reg1_reg_14_, p2_reg1_reg_15_, p2_reg1_reg_16_, p2_reg1_reg_17_,         p2_reg1_reg_18_, p2_reg1_reg_19_, p2_reg1_reg_20_, p2_reg1_reg_21_,         p2_reg1_reg_22_, p2_reg1_reg_23_, p2_reg1_reg_24_, p2_reg1_reg_25_,         p2_reg1_reg_26_, p2_reg1_reg_27_, p2_reg1_reg_28_, p2_reg1_reg_29_,         p2_reg1_reg_30_, p2_reg1_reg_31_, p2_reg2_reg_0_, p2_reg2_reg_1_,         p2_reg2_reg_2_, p2_reg2_reg_3_, p2_reg2_reg_4_, p2_reg2_reg_5_,         p2_reg2_reg_6_, p2_reg2_reg_7_, p2_reg2_reg_8_, p2_reg2_reg_9_,         p2_reg2_reg_10_, p2_reg2_reg_11_, p2_reg2_reg_12_, p2_reg2_reg_13_,         p2_reg2_reg_14_, p2_reg2_reg_15_, p2_reg2_reg_16_, p2_reg2_reg_17_,         p2_reg2_reg_18_, p2_reg2_reg_19_, p2_reg2_reg_20_, p2_reg2_reg_21_,         p2_reg2_reg_22_, p2_reg2_reg_23_, p2_reg2_reg_24_, p2_reg2_reg_25_,         p2_reg2_reg_26_, p2_reg2_reg_27_, p2_reg2_reg_28_, p2_reg2_reg_29_,         p2_reg2_reg_30_, p2_reg2_reg_31_, p2_addr_reg_19_, p2_addr_reg_18_,         p2_addr_reg_17_, p2_addr_reg_16_, p2_addr_reg_15_, p2_addr_reg_14_,         p2_addr_reg_13_, p2_addr_reg_12_, p2_addr_reg_11_, p2_addr_reg_10_,         p2_addr_reg_9_, p2_addr_reg_8_, p2_addr_reg_7_, p2_addr_reg_6_,         p2_addr_reg_5_, p2_addr_reg_4_, p2_addr_reg_3_, p2_addr_reg_2_,         p2_addr_reg_1_, p2_addr_reg_0_, p2_datao_reg_0_, p2_datao_reg_1_,         p2_datao_reg_2_, p2_datao_reg_3_, p2_datao_reg_4_, p2_datao_reg_5_,         p2_datao_reg_6_, p2_datao_reg_7_, p2_datao_reg_8_, p2_datao_reg_9_,         p2_datao_reg_10_, p2_datao_reg_11_, p2_datao_reg_12_,         p2_datao_reg_13_, p2_datao_reg_14_, p2_datao_reg_15_,         p2_datao_reg_16_, p2_datao_reg_17_, p2_datao_reg_18_,         p2_datao_reg_19_, p2_datao_reg_20_, p2_datao_reg_21_,         p2_datao_reg_22_, p2_datao_reg_23_, p2_datao_reg_24_,         p2_datao_reg_25_, p2_datao_reg_26_, p2_datao_reg_27_,         p2_datao_reg_28_, p2_datao_reg_29_, p2_datao_reg_30_,         p2_datao_reg_31_, p2_b_reg, p2_reg3_reg_15_, p2_reg3_reg_26_,         p2_reg3_reg_6_, p2_reg3_reg_18_, p2_reg3_reg_2_, p2_reg3_reg_11_,         p2_reg3_reg_22_, p2_reg3_reg_13_, p2_reg3_reg_20_, p2_reg3_reg_0_,         p2_reg3_reg_9_, p2_reg3_reg_4_, p2_reg3_reg_24_, p2_reg3_reg_17_,         p2_reg3_reg_5_, p2_reg3_reg_16_, p2_reg3_reg_25_, p2_reg3_reg_12_,         p2_reg3_reg_21_, p2_reg3_reg_1_, p2_reg3_reg_8_, p2_reg3_reg_28_,         p2_reg3_reg_19_, p2_reg3_reg_3_, p2_reg3_reg_10_, p2_reg3_reg_23_,         p2_reg3_reg_14_, p2_reg3_reg_27_, p2_reg3_reg_7_, p2_state_reg,         p2_rd_reg, p2_wr_reg;
output add_1068_u4, add_1068_u55, add_1068_u56, add_1068_u57, add_1068_u58,         add_1068_u59, add_1068_u60, add_1068_u61, add_1068_u62, add_1068_u63,         add_1068_u47, add_1068_u48, add_1068_u49, add_1068_u50, add_1068_u51,         add_1068_u52, add_1068_u53, add_1068_u54, add_1068_u5, add_1068_u46,         u126, u123, p1_u3355, p1_u3354, p1_u3353, p1_u3352, p1_u3351,         p1_u3350, p1_u3349, p1_u3348, p1_u3347, p1_u3346, p1_u3345, p1_u3344,         p1_u3343, p1_u3342, p1_u3341, p1_u3340, p1_u3339, p1_u3338, p1_u3337,         p1_u3336, p1_u3335, p1_u3334, p1_u3333, p1_u3332, p1_u3331, p1_u3330,         p1_u3329, p1_u3328, p1_u3327, p1_u3326, p1_u3325, p1_u3324, p1_u3439,         p1_u3440, p1_u3323, p1_u3322, p1_u3321, p1_u3320, p1_u3319, p1_u3318,         p1_u3317, p1_u3316, p1_u3315, p1_u3314, p1_u3313, p1_u3312, p1_u3311,         p1_u3310, p1_u3309, p1_u3308, p1_u3307, p1_u3306, p1_u3305, p1_u3304,         p1_u3303, p1_u3302, p1_u3301, p1_u3300, p1_u3299, p1_u3298, p1_u3297,         p1_u3296, p1_u3295, p1_u3294, p1_u3453, p1_u3456, p1_u3459, p1_u3462,         p1_u3465, p1_u3468, p1_u3471, p1_u3474, p1_u3477, p1_u3480, p1_u3483,         p1_u3486, p1_u3489, p1_u3492, p1_u3495, p1_u3498, p1_u3501, p1_u3504,         p1_u3507, p1_u3509, p1_u3510, p1_u3511, p1_u3512, p1_u3513, p1_u3514,         p1_u3515, p1_u3516, p1_u3517, p1_u3518, p1_u3519, p1_u3520, p1_u3521,         p1_u3522, p1_u3523, p1_u3524, p1_u3525, p1_u3526, p1_u3527, p1_u3528,         p1_u3529, p1_u3530, p1_u3531, p1_u3532, p1_u3533, p1_u3534, p1_u3535,         p1_u3536, p1_u3537, p1_u3538, p1_u3539, p1_u3540, p1_u3541, p1_u3542,         p1_u3543, p1_u3544, p1_u3545, p1_u3546, p1_u3547, p1_u3548, p1_u3549,         p1_u3550, p1_u3551, p1_u3552, p1_u3553, p1_u3293, p1_u3292, p1_u3291,         p1_u3290, p1_u3289, p1_u3288, p1_u3287, p1_u3286, p1_u3285, p1_u3284,         p1_u3283, p1_u3282, p1_u3281, p1_u3280, p1_u3279, p1_u3278, p1_u3277,         p1_u3276, p1_u3275, p1_u3274, p1_u3273, p1_u3272, p1_u3271, p1_u3270,         p1_u3269, p1_u3268, p1_u3267, p1_u3266, p1_u3265, p1_u3356, p1_u3264,         p1_u3263, p1_u3262, p1_u3261, p1_u3260, p1_u3259, p1_u3258, p1_u3257,         p1_u3256, p1_u3255, p1_u3254, p1_u3253, p1_u3252, p1_u3251, p1_u3250,         p1_u3249, p1_u3248, p1_u3247, p1_u3246, p1_u3245, p1_u3244, p1_u3243,         p1_u3554, p1_u3555, p1_u3556, p1_u3557, p1_u3558, p1_u3559, p1_u3560,         p1_u3561, p1_u3562, p1_u3563, p1_u3564, p1_u3565, p1_u3566, p1_u3567,         p1_u3568, p1_u3569, p1_u3570, p1_u3571, p1_u3572, p1_u3573, p1_u3574,         p1_u3575, p1_u3576, p1_u3577, p1_u3578, p1_u3579, p1_u3580, p1_u3581,         p1_u3582, p1_u3583, p1_u3584, p1_u3585, p1_u3242, p1_u3241, p1_u3240,         p1_u3239, p1_u3238, p1_u3237, p1_u3236, p1_u3235, p1_u3234, p1_u3233,         p1_u3232, p1_u3231, p1_u3230, p1_u3229, p1_u3228, p1_u3227, p1_u3226,         p1_u3225, p1_u3224, p1_u3223, p1_u3222, p1_u3221, p1_u3220, p1_u3219,         p1_u3218, p1_u3217, p1_u3216, p1_u3215, p1_u3214, p1_u3213, p1_u3086,         p1_u3085, p1_u3973, p2_u3295, p2_u3294, p2_u3293, p2_u3292, p2_u3291,         p2_u3290, p2_u3289, p2_u3288, p2_u3287, p2_u3286, p2_u3285, p2_u3284,         p2_u3283, p2_u3282, p2_u3281, p2_u3280, p2_u3279, p2_u3278, p2_u3277,         p2_u3276, p2_u3275, p2_u3274, p2_u3273, p2_u3272, p2_u3271, p2_u3270,         p2_u3269, p2_u3268, p2_u3267, p2_u3266, p2_u3265, p2_u3264, p2_u3376,         p2_u3377, p2_u3263, p2_u3262, p2_u3261, p2_u3260, p2_u3259, p2_u3258,         p2_u3257, p2_u3256, p2_u3255, p2_u3254, p2_u3253, p2_u3252, p2_u3251,         p2_u3250, p2_u3249, p2_u3248, p2_u3247, p2_u3246, p2_u3245, p2_u3244,         p2_u3243, p2_u3242, p2_u3241, p2_u3240, p2_u3239, p2_u3238, p2_u3237,         p2_u3236, p2_u3235, p2_u3234, p2_u3390, p2_u3393, p2_u3396, p2_u3399,         p2_u3402, p2_u3405, p2_u3408, p2_u3411, p2_u3414, p2_u3417, p2_u3420,         p2_u3423, p2_u3426, p2_u3429, p2_u3432, p2_u3435, p2_u3438, p2_u3441,         p2_u3444, p2_u3446, p2_u3447, p2_u3448, p2_u3449, p2_u3450, p2_u3451,         p2_u3452, p2_u3453, p2_u3454, p2_u3455, p2_u3456, p2_u3457, p2_u3458,         p2_u3459, p2_u3460, p2_u3461, p2_u3462, p2_u3463, p2_u3464, p2_u3465,         p2_u3466, p2_u3467, p2_u3468, p2_u3469, p2_u3470, p2_u3471, p2_u3472,         p2_u3473, p2_u3474, p2_u3475, p2_u3476, p2_u3477, p2_u3478, p2_u3479,         p2_u3480, p2_u3481, p2_u3482, p2_u3483, p2_u3484, p2_u3485, p2_u3486,         p2_u3487, p2_u3488, p2_u3489, p2_u3490, p2_u3233, p2_u3232, p2_u3231,         p2_u3230, p2_u3229, p2_u3228, p2_u3227, p2_u3226, p2_u3225, p2_u3224,         p2_u3223, p2_u3222, p2_u3221, p2_u3220, p2_u3219, p2_u3218, p2_u3217,         p2_u3216, p2_u3215, p2_u3214, p2_u3213, p2_u3212, p2_u3211, p2_u3210,         p2_u3209, p2_u3208, p2_u3207, p2_u3206, p2_u3205, p2_u3204, p2_u3203,         p2_u3202, p2_u3201, p2_u3200, p2_u3199, p2_u3198, p2_u3197, p2_u3196,         p2_u3195, p2_u3194, p2_u3193, p2_u3192, p2_u3191, p2_u3190, p2_u3189,         p2_u3188, p2_u3187, p2_u3186, p2_u3185, p2_u3184, p2_u3183, p2_u3182,         p2_u3491, p2_u3492, p2_u3493, p2_u3494, p2_u3495, p2_u3496, p2_u3497,         p2_u3498, p2_u3499, p2_u3500, p2_u3501, p2_u3502, p2_u3503, p2_u3504,         p2_u3505, p2_u3506, p2_u3507, p2_u3508, p2_u3509, p2_u3510, p2_u3511,         p2_u3512, p2_u3513, p2_u3514, p2_u3515, p2_u3516, p2_u3517, p2_u3518,         p2_u3519, p2_u3520, p2_u3521, p2_u3522, p2_u3296, p2_u3181, p2_u3180,         p2_u3179, p2_u3178, p2_u3177, p2_u3176, p2_u3175, p2_u3174, p2_u3173,         p2_u3172, p2_u3171, p2_u3170, p2_u3169, p2_u3168, p2_u3167, p2_u3166,         p2_u3165, p2_u3164, p2_u3163, p2_u3162, p2_u3161, p2_u3160, p2_u3159,         p2_u3158, p2_u3157, p2_u3156, p2_u3155, p2_u3154, p2_u3153, p2_u3151,         p2_u3150, p2_u3893;
wire   n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,         n19241, n19242, n19243, n9903, n9904, n9906, n9908, n9910, n9912,         n9914, n9916, n9918, n9920, n9922, n9924, n9926, n9928, n9930, n9932,         n9934, n9936, n9938, n9940, n9942, n10003, n10006, n10009, n10014,         n10017, n10020, n10025, n10028, n10033, n10036, n10047, n10050,         n10053, n10056, n10059, n10062, n10065, n10070, n10075, n10078,         n10281, n10452, n10453, n10454, n10455, n10456, n10457, n10458,         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,         n18771, n18772, n18773, n18774, n18775, n18776;

   nor U9493 ( n17606,n17607,n17608,n17609 );
   nor U9494 ( n17496,n17497,n17498,n17499 );
   nor U9495 ( n17406,n17407,n17408,n17409 );
   nor U9496 ( n11040,n11046,n11047,n11048 );
   or U9497 ( n9903,n14310,n14313 );
   not U9498 ( n15293,n15260 );
   nand U9499 ( n13451,n10650,n14281 );
   nor U9500 ( n11835,n12667,n11836 );
   not U9501 ( n17346,n17417 );
   nand U9502 ( n13450,n11026,n12500,n11031 );
   nand U9503 ( n13467,n11026,n12646,n11031 );
   nand U9504 ( n9904,n10281,p1_d_reg_15_ );
   not U9505 ( p1_u3310,n9904 );
   nand U9506 ( n9906,n14973,p1_d_reg_20_ );
   not U9507 ( p1_u3305,n9906 );
   nand U9508 ( n9908,n14973,p1_d_reg_14_ );
   not U9509 ( p1_u3311,n9908 );
   nand U9510 ( n9910,n10281,p1_d_reg_21_ );
   not U9511 ( p1_u3304,n9910 );
   nand U9512 ( n9912,n10281,p1_d_reg_12_ );
   not U9513 ( p1_u3313,n9912 );
   nand U9514 ( n9914,n14973,p1_d_reg_22_ );
   not U9515 ( p1_u3303,n9914 );
   nand U9516 ( n9916,n14973,p1_d_reg_11_ );
   not U9517 ( p1_u3314,n9916 );
   nand U9518 ( n9918,n14973,p1_d_reg_23_ );
   not U9519 ( p1_u3302,n9918 );
   nand U9520 ( n9920,n10281,p1_d_reg_9_ );
   not U9521 ( p1_u3316,n9920 );
   nand U9522 ( n9922,n14973,p1_d_reg_24_ );
   not U9523 ( p1_u3301,n9922 );
   nand U9524 ( n9924,n14973,p1_d_reg_8_ );
   not U9525 ( p1_u3317,n9924 );
   nand U9526 ( n9926,n10281,p1_d_reg_25_ );
   not U9527 ( p1_u3300,n9926 );
   nand U9528 ( n9928,n10281,p1_d_reg_7_ );
   not U9529 ( p1_u3318,n9928 );
   nand U9530 ( n9930,n14973,p1_d_reg_26_ );
   not U9531 ( p1_u3299,n9930 );
   nand U9532 ( n9932,n10281,p1_d_reg_5_ );
   not U9533 ( p1_u3320,n9932 );
   nand U9534 ( n9934,n10281,p1_d_reg_28_ );
   not U9535 ( p1_u3297,n9934 );
   nand U9536 ( n9936,n14973,p1_d_reg_4_ );
   not U9537 ( p1_u3321,n9936 );
   nand U9538 ( n9938,n14973,p1_d_reg_30_ );
   not U9539 ( p1_u3295,n9938 );
   nand U9540 ( n9940,n14973,p1_d_reg_3_ );
   not U9541 ( p1_u3322,n9940 );
   nand U9542 ( n9942,n10281,p1_d_reg_31_ );
   not U9543 ( p1_u3294,n9942 );
   and U9544 ( n13453,n10650,n14161 );
   buf U9545 ( p2_u3292,n19024 );
   nand U9546 ( n19024,n11569,n11570,n11571,n11572 );
   buf U9547 ( p2_u3293,n19023 );
   nand U9548 ( n19023,n11562,n11563,n11564,n11565 );
   buf U9549 ( p2_u3291,n19025 );
   nand U9550 ( n19025,n11579,n11580,n11581,n11582 );
   buf U9551 ( p2_u3294,n19022 );
   nand U9552 ( n19022,n11552,n11553,n11554,n11555 );
   buf U9553 ( p2_u3290,n19026 );
   nand U9554 ( n19026,n11586,n11587,n11588,n11589 );
   buf U9555 ( p2_u3295,n19021 );
   nand U9556 ( n19021,n11543,n11544,n11545 );
   buf U9557 ( p2_u3289,n19027 );
   nand U9558 ( n19027,n11595,n11596,n11597,n11598 );
   not U9559 ( p1_u3085,n16819 );
   nand U9560 ( n16819,n18638,n14347 );
   buf U9561 ( p2_u3288,n19028 );
   nand U9562 ( n19028,n11602,n11603,n11604,n11605 );
   buf U9563 ( p1_u3218,n19015 );
   nand U9564 ( n19015,n17691,n16730,n17692,n17693 );
   nor U9565 ( n17693,n17694,n17695,n17696 );
   buf U9566 ( p2_u3287,n19029 );
   nand U9567 ( n19029,n11611,n11612,n11613,n11614 );
   buf U9568 ( p1_u3228,n19005 );
   nand U9569 ( n19005,n17519,n17520,n17521,n17522 );
   nand U9570 ( n17520,n17527,n17528,n17366 );
   buf U9571 ( p2_u3286,n19030 );
   nand U9572 ( n19030,n11618,n11619,n11620,n11621 );
   buf U9573 ( p1_u3229,n19004 );
   nand U9574 ( n19004,n17506,n17507,n17508,n17509 );
   buf U9575 ( p2_u3285,n19031 );
   nand U9576 ( n19031,n11627,n11628,n11629,n11630 );
   buf U9577 ( p1_u3230,n19003 );
   nand U9578 ( n19003,n17493,n17494,n17495,n17496 );
   buf U9579 ( p2_u3284,n19032 );
   nand U9580 ( n19032,n11634,n11635,n11636,n11637 );
   buf U9581 ( p1_u3231,n19002 );
   nand U9582 ( n19002,n17481,n17482,n17483,n17484 );
   buf U9583 ( p2_u3283,n19033 );
   nand U9584 ( n19033,n11644,n11645,n11646,n11647 );
   buf U9585 ( p1_u3233,n19000 );
   nand U9586 ( n19000,n17458,n17459,n17460,n17461 );
   buf U9587 ( p2_u3282,n19034 );
   nand U9588 ( n19034,n11651,n11652,n11653,n11654 );
   buf U9589 ( p1_u3234,n18999 );
   nand U9590 ( n18999,n17444,n17445,n17446,n17447 );
   nand U9591 ( n17445,n17451,n17452,n17366 );
   buf U9592 ( p2_u3281,n19035 );
   nand U9593 ( n19035,n11661,n11662,n11663,n11664 );
   buf U9594 ( p1_u3235,n18998 );
   nand U9595 ( n18998,n17431,n17432,n17433,n17434 );
   buf U9596 ( p2_u3280,n19036 );
   nand U9597 ( n19036,n11668,n11669,n11670,n11671 );
   buf U9598 ( p1_u3236,n18997 );
   nand U9599 ( n18997,n17418,n17419,n17420,n17421 );
   nand U9600 ( n17419,n17426,n17366 );
   buf U9601 ( p2_u3279,n19037 );
   nand U9602 ( n19037,n11678,n11679,n11680,n11681 );
   buf U9603 ( p1_u3238,n18995 );
   nand U9604 ( n18995,n17390,n17391,n17392,n17393 );
   buf U9605 ( p2_u3278,n19038 );
   nand U9606 ( n19038,n11685,n11686,n11687,n11688 );
   buf U9607 ( p1_u3239,n18994 );
   nand U9608 ( n18994,n17376,n17377,n17378,n17379 );
   buf U9609 ( p2_u3277,n19039 );
   nand U9610 ( n19039,n11695,n11696,n11697,n11698 );
   buf U9611 ( p1_u3240,n18993 );
   nand U9612 ( n18993,n17357,n17358,n17359,n17360 );
   buf U9613 ( p2_u3276,n19040 );
   nand U9614 ( n19040,n11705,n11706,n11707,n11708 );
   buf U9615 ( p1_u3241,n18992 );
   nand U9616 ( n18992,n17339,n17340,n17341,n17342 );
   or U9617 ( n17340,n17350,n17351 );
   buf U9618 ( p2_u3275,n19041 );
   nand U9619 ( n19041,n11712,n11713,n11714,n11715 );
   buf U9620 ( p1_u3242,n18991 );
   nor U9621 ( n18991,n16822,n16823,n16824 );
   buf U9622 ( p2_u3274,n19042 );
   nand U9623 ( n19042,n11719,n11720,n11721,n11722 );
   buf U9624 ( p1_u3243,n18958 );
   nand U9625 ( n18958,n16798,n16799,n16800,n16801 );
   nand U9626 ( n16801,p1_ir_reg_0_,n16802 );
   buf U9627 ( p2_u3273,n19043 );
   nand U9628 ( n19043,n11728,n11729,n11730,n11731 );
   buf U9629 ( p1_u3244,n18957 );
   nand U9630 ( n18957,n16784,n16785,n16786,n16787 );
   buf U9631 ( p2_u3272,n19044 );
   nand U9632 ( n19044,n11735,n11736,n11737,n11738 );
   buf U9633 ( p1_u3245,n18956 );
   nand U9634 ( n18956,n16751,n16752,n16753,n16754 );
   nor U9635 ( n16754,n16755,n16756,n16757 );
   buf U9636 ( p2_u3271,n19045 );
   nand U9637 ( n19045,n11745,n11746,n11747,n11748 );
   buf U9638 ( p1_u3246,n18955 );
   nand U9639 ( n18955,n16730,n16731,n16732,n16733 );
   buf U9640 ( p2_u3270,n19046 );
   nand U9641 ( n19046,n11752,n11753,n11754,n11755 );
   buf U9642 ( p1_u3248,n18953 );
   nand U9643 ( n18953,n16670,n16671,n16672 );
   nor U9644 ( n16672,n16673,n16674,n16675 );
   buf U9645 ( p2_u3269,n19047 );
   nand U9646 ( n19047,n11762,n11763,n11764,n11765 );
   buf U9647 ( p1_u3249,n18952 );
   nand U9648 ( n18952,n16643,n16644,n16645 );
   nor U9649 ( n16645,n16646,n16647,n16648 );
   buf U9650 ( p2_u3268,n19048 );
   nand U9651 ( n19048,n11769,n11770,n11771,n11772 );
   buf U9652 ( p1_u3250,n18951 );
   nand U9653 ( n18951,n16613,n16614,n16615 );
   nor U9654 ( n16615,n16616,n16617,n16618 );
   buf U9655 ( p2_u3267,n19049 );
   nand U9656 ( n19049,n11779,n11780,n11781,n11782 );
   buf U9657 ( p1_u3251,n18950 );
   nand U9658 ( n18950,n16591,n16592,n16593,n16594 );
   buf U9659 ( p2_u3266,n19050 );
   nand U9660 ( n19050,n11789,n11790,n11791,n11792 );
   buf U9661 ( p1_u3252,n18949 );
   nand U9662 ( n18949,n16567,n16568,n16569 );
   nor U9663 ( n16569,n16570,n16571,n16572 );
   buf U9664 ( p2_u3265,n19051 );
   nand U9665 ( n19051,n11796,n11797,n11798,n11799 );
   buf U9666 ( p1_u3253,n18948 );
   nand U9667 ( n18948,n16542,n16543,n16544,n16545 );
   buf U9668 ( p2_u3264,n19052 );
   nand U9669 ( n19052,n11805,n11806,n11807 );
   buf U9670 ( p1_u3254,n18947 );
   nand U9671 ( n18947,n16513,n16514,n16515,n16516 );
   nand U9672 ( n16516,n16506,n16517 );
   buf U9673 ( p2_u3263,n19055 );
   nor U9674 ( n19055,n11035,n11813 );
   buf U9675 ( p1_u3255,n18946 );
   nand U9676 ( n18946,n16484,n16485,n16486 );
   nor U9677 ( n16486,n16487,n16488,n16489 );
   nand U9678 ( n10003,n11034,p2_d_reg_3_ );
   not U9679 ( p2_u3262,n10003 );
   buf U9680 ( p1_u3256,n18945 );
   nand U9681 ( n18945,n16461,n16462,n16463,n16464 );
   nand U9682 ( n10006,n11034,p2_d_reg_4_ );
   not U9683 ( p2_u3261,n10006 );
   buf U9684 ( p1_u3257,n18944 );
   nand U9685 ( n18944,n16431,n16432,n16433,n16434 );
   nand U9686 ( n10009,n11034,p2_d_reg_5_ );
   not U9687 ( p2_u3260,n10009 );
   buf U9688 ( p1_u3258,n18943 );
   nand U9689 ( n18943,n16405,n16406,n16407,n16408 );
   nand U9690 ( n16408,n16409,n16410 );
   buf U9691 ( p2_u3259,n19056 );
   nor U9692 ( n19056,n11035,n11814 );
   buf U9693 ( p1_u3259,n18942 );
   nand U9694 ( n18942,n16381,n16382,n16383,n16384 );
   nand U9695 ( n16384,n16366,n16385 );
   nand U9696 ( n10014,n11034,p2_d_reg_7_ );
   not U9697 ( p2_u3258,n10014 );
   buf U9698 ( p1_u3260,n18941 );
   nand U9699 ( n18941,n16350,n16351,n16352,n16353 );
   nand U9700 ( n10017,n11034,p2_d_reg_8_ );
   not U9701 ( p2_u3257,n10017 );
   buf U9702 ( p1_u3261,n18940 );
   nand U9703 ( n18940,n16318,n16319,n16320,n16321 );
   nand U9704 ( n16321,n16300,n16322 );
   nand U9705 ( n10020,n11034,p2_d_reg_9_ );
   not U9706 ( p2_u3256,n10020 );
   buf U9707 ( p1_u3262,n18939 );
   nand U9708 ( n18939,n16283,n16284,n16285,n16286 );
   buf U9709 ( p2_u3255,n19057 );
   nor U9710 ( n19057,n11035,n11815 );
   buf U9711 ( p1_u3276,n18924 );
   nand U9712 ( n18924,n15775,n15776,n15777,n15778 );
   nor U9713 ( n15778,n15779,n15780,n15781,n15782 );
   nand U9714 ( n10025,n11034,p2_d_reg_11_ );
   not U9715 ( p2_u3254,n10025 );
   buf U9716 ( p1_u3277,n18923 );
   nand U9717 ( n18923,n15732,n15733,n15734,n15735 );
   nor U9718 ( n15735,n15736,n15737,n15738,n15739 );
   nand U9719 ( n10028,n11034,p2_d_reg_12_ );
   not U9720 ( p2_u3253,n10028 );
   buf U9721 ( p1_u3280,n18920 );
   nand U9722 ( n18920,n15648,n15649,n15650,n15651 );
   nor U9723 ( n15651,n15652,n15653,n15654,n15655 );
   buf U9724 ( p2_u3252,n19058 );
   nor U9725 ( n19058,n11035,n11816 );
   buf U9726 ( p1_u3281,n18919 );
   nand U9727 ( n18919,n15629,n15630,n15631,n15632 );
   nor U9728 ( n15632,n15633,n15634,n15635,n15636 );
   nand U9729 ( n10033,n11034,p2_d_reg_14_ );
   not U9730 ( p2_u3251,n10033 );
   buf U9731 ( p1_u3282,n18918 );
   nand U9732 ( n18918,n15585,n15586,n15587,n15588 );
   nor U9733 ( n15588,n15589,n15590,n15591,n15592 );
   nand U9734 ( n10036,n11034,p2_d_reg_15_ );
   not U9735 ( p2_u3250,n10036 );
   buf U9736 ( p1_u3283,n18917 );
   nand U9737 ( n18917,n15545,n15546,n15547,n15548 );
   nor U9738 ( n15548,n15549,n15550,n15551,n15552 );
   buf U9739 ( p2_u3249,n19059 );
   nor U9740 ( n19059,n11035,n11817 );
   buf U9741 ( p1_u3285,n18915 );
   nand U9742 ( n18915,n15482,n15483,n15484,n15485 );
   nor U9743 ( n15485,n15486,n15487,n15488,n15489 );
   buf U9744 ( p2_u3248,n19060 );
   nor U9745 ( n19060,n11035,n11818 );
   buf U9746 ( p1_u3286,n18914 );
   nand U9747 ( n18914,n15444,n15445,n15446,n15447 );
   nor U9748 ( n15447,n15448,n15449,n15450,n15451 );
   buf U9749 ( p2_u3247,n19061 );
   nor U9750 ( n19061,n11035,n11819 );
   buf U9751 ( p1_u3287,n18913 );
   nand U9752 ( n18913,n15403,n15404,n15405,n15406 );
   nor U9753 ( n15406,n15407,n15408,n15409,n15410 );
   buf U9754 ( p2_u3246,n19062 );
   nor U9755 ( n19062,n11035,n11820 );
   buf U9756 ( p1_u3296,n18842 );
   nor U9757 ( n18842,n14974,n15251 );
   nand U9758 ( n10047,n11034,p2_d_reg_20_ );
   not U9759 ( p2_u3245,n10047 );
   buf U9760 ( p1_u3298,n18841 );
   nor U9761 ( n18841,n14974,n15250 );
   nand U9762 ( n10050,n11034,p2_d_reg_21_ );
   not U9763 ( p2_u3244,n10050 );
   buf U9764 ( p1_u3306,n18840 );
   nor U9765 ( n18840,n14974,n15249 );
   nand U9766 ( n10053,n11034,p2_d_reg_22_ );
   not U9767 ( p2_u3243,n10053 );
   buf U9768 ( p1_u3307,n18839 );
   nor U9769 ( n18839,n14974,n15248 );
   nand U9770 ( n10056,n11034,p2_d_reg_23_ );
   not U9771 ( p2_u3242,n10056 );
   buf U9772 ( p1_u3308,n18838 );
   nor U9773 ( n18838,n14974,n15247 );
   nand U9774 ( n10059,n11034,p2_d_reg_24_ );
   not U9775 ( p2_u3241,n10059 );
   buf U9776 ( p1_u3309,n18837 );
   nor U9777 ( n18837,n14974,n15246 );
   nand U9778 ( n10062,n11034,p2_d_reg_25_ );
   not U9779 ( p2_u3240,n10062 );
   buf U9780 ( p1_u3312,n18836 );
   nor U9781 ( n18836,n14974,n15245 );
   nand U9782 ( n10065,n11034,p2_d_reg_26_ );
   not U9783 ( p2_u3239,n10065 );
   buf U9784 ( p1_u3315,n18835 );
   nor U9785 ( n18835,n14974,n15244 );
   buf U9786 ( p2_u3238,n19063 );
   nor U9787 ( n19063,n11035,n11821 );
   buf U9788 ( p1_u3319,n18834 );
   nor U9789 ( n18834,n14974,n15243 );
   nand U9790 ( n10070,n11034,p2_d_reg_28_ );
   not U9791 ( p2_u3237,n10070 );
   buf U9792 ( p1_u3323,n18833 );
   nor U9793 ( n18833,n14974,n15242 );
   buf U9794 ( p2_u3236,n19064 );
   nor U9795 ( n19064,n11035,n11822 );
   not U9796 ( n11035,n11034 );
   buf U9797 ( p1_u3440,n18832 );
   nand U9798 ( n18832,n14971,n14972 );
   nand U9799 ( n14972,p1_d_reg_1_,n10281 );
   nand U9800 ( n10075,n11034,p2_d_reg_30_ );
   not U9801 ( p2_u3235,n10075 );
   buf U9802 ( p1_u3439,n18831 );
   nand U9803 ( n18831,n14976,n14977 );
   nand U9804 ( n14977,p1_d_reg_0_,n10281 );
   nand U9805 ( n10078,n11034,p2_d_reg_31_ );
   not U9806 ( p2_u3234,n10078 );
   buf U9807 ( p1_u3324,n18830 );
   nand U9808 ( n18830,n15238,n15239,n15240 );
   buf U9809 ( p2_u3232,n19130 );
   nand U9810 ( n19130,n11842,n11843,n11844,n11845 );
   nand U9811 ( n11843,n11856,p2_reg3_reg_1_ );
   nor U9812 ( n11845,n11846,n11847,n11848,n11849 );
   buf U9813 ( p1_u3325,n18829 );
   nand U9814 ( n18829,n15229,n15230,n15231,n15232 );
   buf U9815 ( p2_u3229,n19133 );
   nand U9816 ( n19133,n11911,n11912,n11913,n11914 );
   nand U9817 ( n11912,n11856,n11931 );
   nor U9818 ( n11914,n11915,n11916,n11917,n11918 );
   buf U9819 ( p1_u3326,n18828 );
   nand U9820 ( n18828,n15221,n15222,n15223,n15224 );
   buf U9821 ( p2_u3228,n19134 );
   nand U9822 ( n19134,n11932,n11933,n11934,n11935 );
   nand U9823 ( n11933,n11856,n11953 );
   nor U9824 ( n11935,n11936,n11937,n11938,n11939 );
   buf U9825 ( p1_u3327,n18827 );
   nand U9826 ( n18827,n15215,n15216,n15217,n15218 );
   buf U9827 ( p2_u3224,n19138 );
   nand U9828 ( n19138,n12038,n12039,n12040,n12041 );
   nor U9829 ( n12041,n12042,n12043,n12044,n12045 );
   buf U9830 ( p1_u3328,n18826 );
   nand U9831 ( n18826,n15207,n15208,n15209,n15210 );
   buf U9832 ( p2_u3223,n19139 );
   nand U9833 ( n19139,n12051,n12052,n12053,n12054 );
   nor U9834 ( n12054,n12055,n12056,n12057,n12058 );
   buf U9835 ( p1_u3329,n18825 );
   nand U9836 ( n18825,n15201,n15202,n15203,n15204 );
   buf U9837 ( p2_u3222,n19140 );
   nand U9838 ( n19140,n12073,n12074,n12075,n12076 );
   nor U9839 ( n12076,n12077,n12078,n12079,n12080 );
   buf U9840 ( p1_u3330,n18824 );
   nand U9841 ( n18824,n15193,n15194,n15195,n15196 );
   buf U9842 ( p2_u3216,n19146 );
   nand U9843 ( n19146,n12215,n12216,n12217,n12218 );
   nor U9844 ( n12218,n12219,n12220,n12221,n12222 );
   buf U9845 ( p1_u3331,n18823 );
   nand U9846 ( n18823,n15187,n15188,n15189,n15190 );
   buf U9847 ( p2_u3215,n19147 );
   nand U9848 ( n19147,n12228,n12229,n12230,n12231 );
   nor U9849 ( n12231,n12232,n12233,n12234,n12235 );
   buf U9850 ( p1_u3332,n18822 );
   nand U9851 ( n18822,n15179,n15180,n15181,n15182 );
   buf U9852 ( p2_u3207,n19155 );
   nand U9853 ( n19155,n12409,n12410,n12411,n12412 );
   nand U9854 ( n12409,n11837,n10716 );
   buf U9855 ( p1_u3333,n18821 );
   nand U9856 ( n18821,n15173,n15174,n15175,n15176 );
   buf U9857 ( p2_u3203,n19159 );
   nand U9858 ( n19159,n12647,n12648,n12649 );
   buf U9859 ( p1_u3334,n18820 );
   nand U9860 ( n18820,n15165,n15166,n15167,n15168 );
   buf U9861 ( p2_u3202,n19160 );
   nand U9862 ( n19160,n12652,n12653,n12649 );
   buf U9863 ( p1_u3335,n18819 );
   nand U9864 ( n18819,n15159,n15160,n15161,n15162 );
   buf U9865 ( p2_u3200,n19162 );
   nand U9866 ( n19162,n12724,n12725,n12726,n12727 );
   nand U9867 ( n12727,n12706,n12728 );
   buf U9868 ( p1_u3336,n18818 );
   nand U9869 ( n18818,n15153,n15154,n15155,n15156 );
   buf U9870 ( p2_u3199,n19163 );
   nand U9871 ( n19163,n12759,n12760,n12761,n12762 );
   nand U9872 ( n12762,n12748,n12763 );
   buf U9873 ( p1_u3337,n18817 );
   nand U9874 ( n18817,n15144,n15145,n15146,n15147 );
   buf U9875 ( p2_u3197,n19165 );
   nand U9876 ( n19165,n12837,n12838,n12839,n12840 );
   buf U9877 ( p1_u3338,n18816 );
   nand U9878 ( n18816,n15136,n15137,n15138,n15139 );
   buf U9879 ( p2_u3196,n19166 );
   nand U9880 ( n19166,n12879,n12880,n12881,n12882 );
   buf U9881 ( p1_u3339,n18815 );
   nand U9882 ( n18815,n15130,n15131,n15132,n15133 );
   buf U9883 ( p2_u3195,n19167 );
   nand U9884 ( n19167,n12916,n12917,n12918,n12919 );
   nand U9885 ( n12919,n12897,n12920 );
   buf U9886 ( p1_u3340,n18814 );
   nand U9887 ( n18814,n15121,n15122,n15123,n15124 );
   buf U9888 ( p2_u3194,n19168 );
   nand U9889 ( n19168,n12952,n12953,n12954,n12955 );
   buf U9890 ( p1_u3341,n18813 );
   nand U9891 ( n18813,n15115,n15116,n15117,n15118 );
   buf U9892 ( p2_u3192,n19170 );
   nand U9893 ( n19170,n13037,n13038,n13039,n13040 );
   buf U9894 ( p1_u3342,n18812 );
   nand U9895 ( n18812,n15107,n15108,n15109,n15110 );
   buf U9896 ( p2_u3191,n19171 );
   nand U9897 ( n19171,n13074,n13075,n13076,n13077 );
   nand U9898 ( n13077,n12978,n13078 );
   buf U9899 ( p1_u3343,n18811 );
   nand U9900 ( n18811,n15101,n15102,n15103,n15104 );
   buf U9901 ( p2_u3190,n19172 );
   nand U9902 ( n19172,n13111,n13112,n13113,n13114 );
   buf U9903 ( p1_u3344,n18810 );
   nand U9904 ( n18810,n15096,n15097,n15098,n15099 );
   buf U9905 ( p2_u3189,n19173 );
   nand U9906 ( n19173,n13155,n13156,n13157,n13158 );
   buf U9907 ( p1_u3345,n18809 );
   nand U9908 ( n18809,n15090,n15091,n15092,n15093 );
   buf U9909 ( p2_u3188,n19174 );
   nand U9910 ( n19174,n13190,n13191,n13192,n13193 );
   buf U9911 ( p1_u3346,n18808 );
   nand U9912 ( n18808,n15085,n15086,n15087,n15088 );
   buf U9913 ( p2_u3187,n19175 );
   nand U9914 ( n19175,n13231,n13232,n13233,n13234 );
   nand U9915 ( n13234,n13235,n13204,n12701 );
   buf U9916 ( p1_u3347,n18807 );
   nand U9917 ( n18807,n15079,n15080,n15081,n15082 );
   buf U9918 ( p2_u3183,n19179 );
   nand U9919 ( n19179,n13392,n13393,n13394,n13395 );
   nand U9920 ( n13395,n13373,n13396 );
   buf U9921 ( p1_u3348,n18806 );
   nand U9922 ( n18806,n15071,n15072,n15073,n15074 );
   buf U9923 ( p2_u3296,n19213 );
   nor U9924 ( n19213,n11040,n11041 );
   buf U9925 ( p1_u3349,n18805 );
   nand U9926 ( n18805,n15065,n15066,n15067,n15068 );
   buf U9927 ( p2_u3181,n19214 );
   nand U9928 ( n19214,n13443,n13444,n13445,n13446 );
   buf U9929 ( p1_u3350,n18804 );
   nand U9930 ( n18804,n15056,n15057,n15058,n15059 );
   buf U9931 ( p2_u3180,n19215 );
   nand U9932 ( n19215,n13460,n13461,n13462,n13463 );
   buf U9933 ( p1_u3351,n18803 );
   nand U9934 ( n18803,n15050,n15051,n15052,n15053 );
   buf U9935 ( p2_u3179,n19216 );
   nand U9936 ( n19216,n13481,n13482,n13483,n13484 );
   buf U9937 ( p1_u3352,n18802 );
   nand U9938 ( n18802,n15045,n15046,n15047,n15048 );
   buf U9939 ( p2_u3178,n19217 );
   nand U9940 ( n19217,n13498,n13499,n13500,n13501 );
   buf U9941 ( p1_u3353,n18801 );
   nand U9942 ( n18801,n15039,n15040,n15041,n15042 );
   buf U9943 ( p2_u3177,n19218 );
   nand U9944 ( n19218,n13510,n13511,n13512,n13513 );
   buf U9945 ( p1_u3354,n18800 );
   nand U9946 ( n18800,n15034,n15035,n15036,n15037 );
   buf U9947 ( p2_u3175,n19220 );
   nand U9948 ( n19220,n13543,n13544,n13545,n13546 );
   buf U9949 ( p1_u3355,n18799 );
   nand U9950 ( n18799,n15026,n15027,n15028 );
   buf U9951 ( p2_u3171,n19224 );
   nand U9952 ( n19224,n13591,n13592,n13593,n13594 );
   buf U9953 ( u123,n18798 );
   xor U9954 ( n18798,n10453,p1_wr_reg );
   buf U9955 ( p2_u3170,n19225 );
   nand U9956 ( n19225,n13602,n13603,n13604,n13605 );
   buf U9957 ( u126,n18797 );
   xor U9958 ( n18797,n10452,p1_rd_reg );
   buf U9959 ( p2_u3169,n19226 );
   nand U9960 ( n19226,n13613,n13614,n13615,n13616 );
   buf U9961 ( add_1068_u46,n18796 );
   xor U9962 ( n18796,p2_addr_reg_0_,p1_addr_reg_0_ );
   buf U9963 ( p2_u3158,n19237 );
   nand U9964 ( n19237,n13770,n13771,n13772,n13773 );
   and U9965 ( n17676,n18545,n18546 );
   nand U9966 ( n15292,n16277,n14996 );
   and U9967 ( n13758,n14269,n14270 );
   nor U9968 ( n15032,n15031,p1_u3086 );
   nor U9969 ( n11549,n11548,p2_u3151 );
   not U9970 ( n16884,n16883 );
   nand U9971 ( n16883,n14968,n16288 );
   nand U9972 ( n11186,n11492,n11368 );
   nand U9973 ( n11187,n11493,n11494 );
   not U9974 ( p1_u3086,p1_state_reg );
   not U9975 ( p2_u3151,p2_state_reg );
   buf U9976 ( p1_u3237,n18996 );
   nand U9977 ( n18996,n17404,n17405,n17406 );
   buf U9978 ( p1_u3264,n18937 );
   nand U9979 ( n18937,n16260,n16261,n16262,n16263 );
   buf U9980 ( p2_u3226,n19136 );
   nand U9981 ( n19136,n11981,n11982,n11983,n11984 );
   nor U9982 ( n11984,n11985,n11986,n11987,n11988 );
   buf U9983 ( p1_u3273,n18927 );
   nand U9984 ( n18927,n15846,n15847,n15848,n15849 );
   nor U9985 ( n15849,n15850,n15851,n15852,n15853 );
   buf U9986 ( p2_u3230,n19132 );
   nand U9987 ( n19132,n11890,n11891,n11892,n11893 );
   nand U9988 ( n11891,n11856,n11910 );
   nor U9989 ( n11893,n11894,n11895,n11896,n11897 );
   buf U9990 ( p1_u3227,n19006 );
   nand U9991 ( n19006,n17534,n17535,n17536,n17537 );
   buf U9992 ( p2_u3176,n19219 );
   nand U9993 ( n19219,n13527,n13528,n13529,n13530 );
   buf U9994 ( p2_u3168,n19227 );
   nand U9995 ( n19227,n13626,n13627,n13628,n13629 );
   buf U9996 ( p2_u3217,n19145 );
   nand U9997 ( n19145,n12195,n12196,n12197,n12198 );
   nor U9998 ( n12198,n12199,n12200,n12201,n12202 );
   buf U9999 ( p1_u3290,n18910 );
   nand U10000 ( n18910,n15324,n15325,n15326,n15327 );
   nor U10001 ( n15327,n15328,n15329,n15330,n15331 );
   buf U10002 ( p1_u3267,n18933 );
   nand U10003 ( n18933,n16022,n16023,n16024,n16025 );
   nor U10004 ( n16025,n16026,n16027,n16028,n16029 );
   buf U10005 ( p1_u3226,n19007 );
   nand U10006 ( n19007,n17546,n17547,n17548,n17549 );
   nand U10007 ( n17547,n17555,n17366 );
   buf U10008 ( p2_u3233,n19129 );
   nand U10009 ( n19129,n11823,n11824,n11825,n11826 );
   nor U10010 ( n11826,n11827,n11828,n11829 );
   buf U10011 ( p2_u3173,n19222 );
   nand U10012 ( n19222,n13574,n13575,n13576,n13577 );
   buf U10013 ( p2_u3164,n19231 );
   nand U10014 ( n19231,n13678,n13679,n13680,n13681 );
   buf U10015 ( p1_u3222,n19011 );
   nand U10016 ( n19011,n17604,n17605,n17606 );
   buf U10017 ( p2_u3210,n19152 );
   nand U10018 ( n19152,n12358,n12359,n12360,n12361 );
   nor U10019 ( n12361,n12362,n12363,n12364,n12365 );
   buf U10020 ( p1_u3278,n18922 );
   nand U10021 ( n18922,n15712,n15713,n15714,n15715 );
   buf U10022 ( p1_u3270,n18930 );
   nand U10023 ( n18930,n15946,n15947,n15948,n15949 );
   nor U10024 ( n15949,n15950,n15951,n15952,n15953 );
   buf U10025 ( p1_u3224,n19009 );
   nand U10026 ( n19009,n17576,n17577,n17578,n17579 );
   buf U10027 ( p2_u3231,n19131 );
   nand U10028 ( n19131,n11857,n11858,n11859,n11860 );
   nor U10029 ( n11860,n11861,n11862,n11863 );
   buf U10030 ( p2_u3174,n19221 );
   nand U10031 ( n19221,n13555,n13556,n13557,n13558 );
   buf U10032 ( p2_u3163,n19232 );
   nand U10033 ( n19232,n13695,n13696,n13697,n13698 );
   not U10034 ( n11856,n11834 );
   buf U10035 ( p1_u3266,n18934 );
   nand U10036 ( n18934,n16065,n16066,n16067,n16068 );
   nor U10037 ( n16068,n16069,n16070,n16071,n16072 );
   buf U10038 ( p1_u3291,n18909 );
   nand U10039 ( n18909,n15294,n15295,n15296,n15297 );
   nor U10040 ( n15297,n15298,n15299,n15300,n15301 );
   buf U10041 ( p2_u3212,n19150 );
   nand U10042 ( n19150,n12301,n12302,n12303,n12304 );
   nor U10043 ( n12304,n12305,n12306,n12307,n12308 );
   buf U10044 ( p1_u3225,n19008 );
   nand U10045 ( n19008,n17560,n17561,n17562,n17563 );
   buf U10046 ( p1_u3221,n19012 );
   nand U10047 ( n19012,n17615,n17616,n17617,n17618 );
   buf U10048 ( p2_u3227,n19135 );
   nand U10049 ( n19135,n11954,n11955,n11956,n11957 );
   nor U10050 ( n11957,n11958,n11959,n11960 );
   buf U10051 ( p2_u3166,n19229 );
   nand U10052 ( n19229,n13655,n13656,n13657,n13658 );
   buf U10053 ( p2_u3161,n19234 );
   nand U10054 ( n19234,n13720,n13721,n13722,n13723 );
   not U10055 ( n16273,n18592 );
   nand U10056 ( n15320,n18360,n17135,n16288 );
   nor U10057 ( n12666,n11808,n13907 );
   not U10058 ( n13907,n12644 );
   buf U10059 ( p2_u3198,n19164 );
   nand U10060 ( n19164,n12793,n12794,n12795 );
   buf U10061 ( p1_u3272,n18928 );
   nand U10062 ( n18928,n15884,n15885,n15886,n15887 );
   nor U10063 ( n15887,n15888,n15889,n15890,n15891 );
   buf U10064 ( p1_u3271,n18929 );
   nand U10065 ( n18929,n15922,n15923,n15924,n15925 );
   buf U10066 ( p1_u3220,n19013 );
   nand U10067 ( n19013,n17629,n17630,n17631,n17632 );
   nand U10068 ( n17630,n17637,n17638,n17366 );
   buf U10069 ( p2_u3225,n19137 );
   nand U10070 ( n19137,n12004,n12005,n12006,n12007 );
   nand U10071 ( n12004,n11837,n10925 );
   buf U10072 ( p2_u3214,n19148 );
   nand U10073 ( n19148,n12244,n12245,n12246,n12247 );
   nor U10074 ( n12247,n12248,n12249,n12250 );
   buf U10075 ( p2_u3165,n19230 );
   nand U10076 ( n19230,n13666,n13667,n13668,n13669 );
   buf U10077 ( p2_u3160,n19235 );
   nand U10078 ( n19235,n13732,n13733,n13734,n13735 );
   not U10079 ( n15241,p1_ir_reg_31_ );
   nand U10080 ( n11831,n11837,n10696 );
   not U10081 ( n10696,n10729 );
   nand U10082 ( n14596,n16187,n16272 );
   buf U10083 ( p2_u3519,n19209 );
   nand U10084 ( n19209,n10464,n10465 );
   buf U10085 ( p2_u3193,n19169 );
   nand U10086 ( n19169,n12996,n12997,n12998 );
   buf U10087 ( p1_u3263,n18938 );
   nand U10088 ( n18938,n16265,n16266,n16262,n16267 );
   buf U10089 ( p1_u3275,n18925 );
   nand U10090 ( n18925,n15807,n15808,n15809,n15810 );
   buf U10091 ( p1_u3292,n18908 );
   nand U10092 ( n18908,n15269,n15270,n15271,n15272 );
   nor U10093 ( n15272,n15273,n15274,n15275,n15276 );
   buf U10094 ( p1_u3223,n19010 );
   nand U10095 ( n19010,n17589,n17590,n17591,n17592 );
   buf U10096 ( p1_u3217,n19016 );
   nand U10097 ( n19016,n17704,n17705,n17706,n17707 );
   or U10098 ( n17705,n17712,n17351 );
   buf U10099 ( p2_u3220,n19142 );
   nand U10100 ( n19142,n12116,n12117,n12118,n12119 );
   nand U10101 ( n12116,n11837,n10862 );
   buf U10102 ( p2_u3218,n19144 );
   nand U10103 ( n19144,n12167,n12168,n12169,n12170 );
   nor U10104 ( n12170,n12171,n12172,n12173 );
   buf U10105 ( p2_u3167,n19228 );
   nand U10106 ( n19228,n13640,n13641,n13642,n13643 );
   buf U10107 ( p2_u3159,n19236 );
   nand U10108 ( n19236,n13759,n13760,n13761,n13762 );
   nand U10109 ( n16288,n18634,n18635 );
   nand U10110 ( n15013,n18359,n17135 );
   nand U10111 ( n16291,n16774,n16188,n16805 );
   not U10112 ( n12716,n12806 );
   nor U10113 ( n12527,n14270,n14269 );
   nor U10114 ( n17286,n18546,n18547 );
   nand U10115 ( n17660,n18192,n18538 );
   buf U10116 ( p2_u3390,n19065 );
   nand U10117 ( n19065,n11010,n11011 );
   nand U10118 ( n11010,n10671,n10648 );
   nand U10119 ( n11011,n10670,p2_reg0_reg_0_ );
   buf U10120 ( p2_u3393,n19066 );
   nand U10121 ( n19066,n10997,n10998 );
   nand U10122 ( n10998,n10670,p2_reg0_reg_1_ );
   buf U10123 ( p2_u3396,n19067 );
   nand U10124 ( n19067,n10988,n10989 );
   nand U10125 ( n10989,n10670,p2_reg0_reg_2_ );
   buf U10126 ( p2_u3399,n19068 );
   nand U10127 ( n19068,n10974,n10975 );
   nand U10128 ( n10975,n10670,p2_reg0_reg_3_ );
   buf U10129 ( p2_u3402,n19069 );
   nand U10130 ( n19069,n10962,n10963 );
   buf U10131 ( p2_u3405,n19070 );
   nand U10132 ( n19070,n10949,n10950 );
   buf U10133 ( p2_u3408,n19071 );
   nand U10134 ( n19071,n10940,n10941 );
   buf U10135 ( p2_u3411,n19072 );
   nand U10136 ( n19072,n10926,n10927 );
   buf U10137 ( p2_u3414,n19073 );
   nand U10138 ( n19073,n10917,n10918 );
   buf U10139 ( p2_u3417,n19074 );
   nand U10140 ( n19074,n10905,n10906 );
   buf U10141 ( p2_u3420,n19075 );
   nand U10142 ( n19075,n10892,n10893 );
   buf U10143 ( p2_u3423,n19076 );
   nand U10144 ( n19076,n10878,n10879 );
   buf U10145 ( p2_u3426,n19077 );
   nand U10146 ( n19077,n10863,n10864 );
   buf U10147 ( p2_u3429,n19078 );
   nand U10148 ( n19078,n10854,n10855 );
   buf U10149 ( p2_u3432,n19079 );
   nand U10150 ( n19079,n10845,n10846 );
   buf U10151 ( p2_u3435,n19080 );
   nand U10152 ( n19080,n10837,n10838 );
   buf U10153 ( p2_u3438,n19081 );
   nand U10154 ( n19081,n10826,n10827 );
   buf U10155 ( p2_u3441,n19082 );
   nand U10156 ( n19082,n10813,n10814 );
   buf U10157 ( p2_u3444,n19083 );
   nand U10158 ( n19083,n10799,n10800 );
   buf U10159 ( p2_u3446,n19084 );
   nand U10160 ( n19084,n10791,n10792 );
   buf U10161 ( p2_u3447,n19085 );
   nand U10162 ( n19085,n10783,n10784 );
   buf U10163 ( p2_u3448,n19086 );
   nand U10164 ( n19086,n10772,n10773 );
   buf U10165 ( p2_u3449,n19087 );
   nand U10166 ( n19087,n10763,n10764 );
   buf U10167 ( p2_u3450,n19088 );
   nand U10168 ( n19088,n10750,n10751 );
   buf U10169 ( p2_u3451,n19089 );
   nand U10170 ( n19089,n10736,n10737 );
   buf U10171 ( p2_u3452,n19090 );
   nand U10172 ( n19090,n10717,n10718 );
   buf U10173 ( p2_u3453,n19091 );
   nand U10174 ( n19091,n10706,n10707 );
   buf U10175 ( p2_u3454,n19092 );
   nand U10176 ( n19092,n10698,n10699 );
   buf U10177 ( p2_u3455,n19093 );
   nand U10178 ( n19093,n10689,n10690 );
   buf U10179 ( p2_u3456,n19094 );
   nand U10180 ( n19094,n10680,n10681 );
   buf U10181 ( p2_u3457,n19095 );
   nand U10182 ( n19095,n10676,n10677 );
   buf U10183 ( p2_u3458,n19096 );
   nand U10184 ( n19096,n10668,n10669 );
   buf U10185 ( p1_u3553,n18906 );
   nand U10186 ( n18906,n14442,n14443 );
   nand U10187 ( n14443,n14444,n14445 );
   buf U10188 ( p1_u3453,n18843 );
   nand U10189 ( n18843,n14949,n14950 );
   nand U10190 ( n14950,n14545,n14539 );
   buf U10191 ( p1_u3456,n18844 );
   nand U10192 ( n18844,n14932,n14933 );
   nand U10193 ( n14933,n14545,n14536 );
   buf U10194 ( p1_u3459,n18845 );
   nand U10195 ( n18845,n14918,n14919 );
   nand U10196 ( n14919,n14545,n14533 );
   buf U10197 ( p1_u3462,n18846 );
   nand U10198 ( n18846,n14906,n14907 );
   nand U10199 ( n14907,n14545,n14530 );
   buf U10200 ( p1_u3465,n18847 );
   nand U10201 ( n18847,n14890,n14891 );
   nand U10202 ( n14891,n14545,n14527 );
   buf U10203 ( p1_u3468,n18848 );
   nand U10204 ( n18848,n14874,n14875 );
   nand U10205 ( n14875,n14545,n14524 );
   buf U10206 ( p1_u3471,n18849 );
   nand U10207 ( n18849,n14862,n14863 );
   nand U10208 ( n14863,n14545,n14521 );
   buf U10209 ( p1_u3474,n18850 );
   nand U10210 ( n18850,n14851,n14852 );
   nand U10211 ( n14852,n14545,n14518 );
   buf U10212 ( p1_u3477,n18851 );
   nand U10213 ( n18851,n14839,n14840 );
   nand U10214 ( n14840,n14545,n14515 );
   buf U10215 ( p1_u3480,n18852 );
   nand U10216 ( n18852,n14824,n14825 );
   nand U10217 ( n14825,n14545,n14512 );
   buf U10218 ( p1_u3483,n18853 );
   nand U10219 ( n18853,n14813,n14814 );
   nand U10220 ( n14814,n14545,n14509 );
   buf U10221 ( p1_u3486,n18854 );
   nand U10222 ( n18854,n14801,n14802 );
   nand U10223 ( n14802,n14545,n14506 );
   buf U10224 ( p1_u3489,n18855 );
   nand U10225 ( n18855,n14785,n14786 );
   nand U10226 ( n14786,n14545,n14503 );
   buf U10227 ( p1_u3492,n18856 );
   nand U10228 ( n18856,n14774,n14775 );
   nand U10229 ( n14775,n14545,n14500 );
   buf U10230 ( p1_u3495,n18857 );
   nand U10231 ( n18857,n14760,n14761 );
   nand U10232 ( n14761,n14545,n14497 );
   buf U10233 ( p1_u3498,n18858 );
   nand U10234 ( n18858,n14746,n14747 );
   nand U10235 ( n14747,n14545,n14494 );
   buf U10236 ( p1_u3501,n18859 );
   nand U10237 ( n18859,n14735,n14736 );
   nand U10238 ( n14736,n14545,n14491 );
   buf U10239 ( p1_u3504,n18860 );
   nand U10240 ( n18860,n14724,n14725 );
   nand U10241 ( n14725,n14545,n14488 );
   buf U10242 ( p1_u3507,n18861 );
   nand U10243 ( n18861,n14709,n14710 );
   nand U10244 ( n14710,n14545,n14485 );
   buf U10245 ( p1_u3509,n18862 );
   nand U10246 ( n18862,n14694,n14695 );
   nand U10247 ( n14695,n14545,n14482 );
   buf U10248 ( p1_u3510,n18863 );
   nand U10249 ( n18863,n14683,n14684 );
   nand U10250 ( n14684,n14545,n14479 );
   buf U10251 ( p1_u3511,n18864 );
   nand U10252 ( n18864,n14671,n14672 );
   nand U10253 ( n14672,n14545,n14476 );
   buf U10254 ( p1_u3512,n18865 );
   nand U10255 ( n18865,n14658,n14659 );
   nand U10256 ( n14659,n14545,n14473 );
   buf U10257 ( p1_u3513,n18866 );
   nand U10258 ( n18866,n14647,n14648 );
   nand U10259 ( n14648,n14545,n14470 );
   buf U10260 ( p1_u3514,n18867 );
   nand U10261 ( n18867,n14631,n14632 );
   nand U10262 ( n14632,n14545,n14467 );
   buf U10263 ( p1_u3515,n18868 );
   nand U10264 ( n18868,n14611,n14612 );
   nand U10265 ( n14612,n14545,n14464 );
   buf U10266 ( p1_u3516,n18869 );
   nand U10267 ( n18869,n14598,n14599 );
   nand U10268 ( n14599,n14545,n14461 );
   buf U10269 ( p1_u3517,n18870 );
   nand U10270 ( n18870,n14585,n14586 );
   nand U10271 ( n14586,n14545,n14458 );
   buf U10272 ( p1_u3518,n18871 );
   nand U10273 ( n18871,n14573,n14574 );
   nand U10274 ( n14574,n14545,n14455 );
   buf U10275 ( p1_u3519,n18872 );
   nand U10276 ( n18872,n14562,n14563 );
   nand U10277 ( n14563,n14545,n14452 );
   buf U10278 ( p1_u3520,n18873 );
   nand U10279 ( n18873,n14554,n14555 );
   nand U10280 ( n14555,n14545,n14449 );
   buf U10281 ( p2_u3376,n19053 );
   nand U10282 ( n19053,n11037,n11038 );
   buf U10283 ( p1_u3576,n18981 );
   nand U10284 ( n18981,n14373,n14374 );
   buf U10285 ( p1_u3583,n18988 );
   nand U10286 ( n18988,n14352,n14353 );
   buf U10287 ( p2_u3512,n19202 );
   nand U10288 ( n19202,n10485,n10486 );
   buf U10289 ( p2_u3514,n19204 );
   nand U10290 ( n19204,n10479,n10480 );
   buf U10291 ( p2_u3186,n19176 );
   nand U10292 ( n19176,n13270,n13271,n13272 );
   nor U10293 ( n13272,n13273,n13274,n13275 );
   buf U10294 ( p2_u3221,n19141 );
   nand U10295 ( n19141,n12094,n12095,n12096,n12097 );
   nand U10296 ( n12094,n11853,n10875 );
   nor U10297 ( n12097,n12098,n12099,n12100,n12101 );
   buf U10298 ( p1_u3289,n18911 );
   nand U10299 ( n18911,n15351,n15352,n15353,n15354 );
   nor U10300 ( n15354,n15355,n15356,n15357,n15358 );
   buf U10301 ( p1_u3274,n18926 );
   nand U10302 ( n18926,n15828,n15829,n15830,n15831 );
   buf U10303 ( p1_u3284,n18916 );
   nand U10304 ( n18916,n15522,n15523,n15524,n15525 );
   nor U10305 ( n15525,n15526,n15527,n15528,n15529 );
   buf U10306 ( p1_u3215,n19018 );
   nand U10307 ( n19018,n17730,n17731,n17732,n17733 );
   buf U10308 ( p1_u3214,n19019 );
   nand U10309 ( n19019,n17744,n17745,n17746,n17747 );
   buf U10310 ( p2_u3219,n19143 );
   nand U10311 ( n19143,n12138,n12139,n12140,n12141 );
   nand U10312 ( n12138,n11837,n10853 );
   buf U10313 ( p2_u3206,n19156 );
   nand U10314 ( n19156,n12438,n12439,n12440,n12441 );
   nor U10315 ( n12441,n12442,n12443,n12444 );
   buf U10316 ( p2_u3162,n19233 );
   nand U10317 ( n19233,n13709,n13710,n13711,n13712 );
   buf U10318 ( p2_u3157,n19238 );
   nand U10319 ( n19238,n13784,n13785,n13786,n13787 );
   buf U10320 ( p2_u3156,n19239 );
   nand U10321 ( n19239,n13799,n13800,n13801,n13802 );
   nor U10322 ( n15667,n15427,n15666 );
   nor U10323 ( n16036,n15427,n16040 );
   nor U10324 ( n15463,n15427,n15462 );
   not U10325 ( n16096,n15427 );
   nor U10326 ( n12665,n11812,n13907 );
   not U10327 ( n12690,n12804 );
   nand U10328 ( n12804,n12659,n13427 );
   not U10329 ( n14623,n14550 );
   nand U10330 ( n10730,n10660,n11030 );
   nor U10331 ( n12526,n14270,n14271 );
   nor U10332 ( n17285,n18546,n18545 );
   not U10333 ( n12713,n11159 );
   nand U10334 ( n12806,n11159,n13427 );
   nand U10335 ( n11159,n14341,n14342,n11786 );
   nand U10336 ( n10281,n14541,n15252 );
   not U10337 ( n14974,n10281 );
   nor U10338 ( n14541,n16820,p1_u3086,n16817 );
   nand U10339 ( n15252,n18629,n18630,n18631 );
   not U10340 ( n13850,n13751 );
   not U10341 ( n17655,n18192 );
   not U10342 ( n17479,n17657 );
   buf U10343 ( p2_u3490,n19128 );
   nand U10344 ( n19128,n10551,n10552 );
   nand U10345 ( n10552,n10553,n10554 );
   buf U10346 ( p1_u3521,n18874 );
   nand U10347 ( n18874,n14543,n14544 );
   nand U10348 ( n14544,n14545,n14445 );
   buf U10349 ( p2_u3377,n19054 );
   nand U10350 ( n19054,n11032,n11033 );
   buf U10351 ( p2_u3459,n19097 );
   nand U10352 ( n19097,n10646,n10647 );
   buf U10353 ( p2_u3460,n19098 );
   nand U10354 ( n19098,n10643,n10644 );
   buf U10355 ( p2_u3461,n19099 );
   nand U10356 ( n19099,n10640,n10641 );
   buf U10357 ( p2_u3462,n19100 );
   nand U10358 ( n19100,n10637,n10638 );
   buf U10359 ( p2_u3463,n19101 );
   nand U10360 ( n19101,n10634,n10635 );
   buf U10361 ( p2_u3464,n19102 );
   nand U10362 ( n19102,n10631,n10632 );
   buf U10363 ( p2_u3465,n19103 );
   nand U10364 ( n19103,n10628,n10629 );
   buf U10365 ( p2_u3466,n19104 );
   nand U10366 ( n19104,n10625,n10626 );
   buf U10367 ( p2_u3467,n19105 );
   nand U10368 ( n19105,n10622,n10623 );
   buf U10369 ( p2_u3468,n19106 );
   nand U10370 ( n19106,n10619,n10620 );
   buf U10371 ( p2_u3469,n19107 );
   nand U10372 ( n19107,n10616,n10617 );
   buf U10373 ( p2_u3470,n19108 );
   nand U10374 ( n19108,n10613,n10614 );
   buf U10375 ( p2_u3471,n19109 );
   nand U10376 ( n19109,n10610,n10611 );
   buf U10377 ( p2_u3472,n19110 );
   nand U10378 ( n19110,n10607,n10608 );
   buf U10379 ( p2_u3473,n19111 );
   nand U10380 ( n19111,n10604,n10605 );
   buf U10381 ( p2_u3474,n19112 );
   nand U10382 ( n19112,n10601,n10602 );
   buf U10383 ( p2_u3475,n19113 );
   nand U10384 ( n19113,n10598,n10599 );
   buf U10385 ( p2_u3476,n19114 );
   nand U10386 ( n19114,n10595,n10596 );
   buf U10387 ( p2_u3477,n19115 );
   nand U10388 ( n19115,n10592,n10593 );
   buf U10389 ( p2_u3478,n19116 );
   nand U10390 ( n19116,n10589,n10590 );
   buf U10391 ( p2_u3479,n19117 );
   nand U10392 ( n19117,n10586,n10587 );
   buf U10393 ( p2_u3480,n19118 );
   nand U10394 ( n19118,n10583,n10584 );
   buf U10395 ( p2_u3481,n19119 );
   nand U10396 ( n19119,n10580,n10581 );
   buf U10397 ( p2_u3482,n19120 );
   nand U10398 ( n19120,n10577,n10578 );
   buf U10399 ( p2_u3483,n19121 );
   nand U10400 ( n19121,n10574,n10575 );
   buf U10401 ( p2_u3484,n19122 );
   nand U10402 ( n19122,n10571,n10572 );
   buf U10403 ( p2_u3485,n19123 );
   nand U10404 ( n19123,n10568,n10569 );
   buf U10405 ( p2_u3486,n19124 );
   nand U10406 ( n19124,n10565,n10566 );
   buf U10407 ( p2_u3487,n19125 );
   nand U10408 ( n19125,n10562,n10563 );
   buf U10409 ( p2_u3488,n19126 );
   nand U10410 ( n19126,n10559,n10560 );
   buf U10411 ( p2_u3489,n19127 );
   nand U10412 ( n19127,n10556,n10557 );
   buf U10413 ( p1_u3522,n18875 );
   nand U10414 ( n18875,n14537,n14538 );
   buf U10415 ( p1_u3523,n18876 );
   nand U10416 ( n18876,n14534,n14535 );
   buf U10417 ( p1_u3524,n18877 );
   nand U10418 ( n18877,n14531,n14532 );
   buf U10419 ( p1_u3525,n18878 );
   nand U10420 ( n18878,n14528,n14529 );
   buf U10421 ( p1_u3526,n18879 );
   nand U10422 ( n18879,n14525,n14526 );
   buf U10423 ( p1_u3527,n18880 );
   nand U10424 ( n18880,n14522,n14523 );
   buf U10425 ( p1_u3528,n18881 );
   nand U10426 ( n18881,n14519,n14520 );
   buf U10427 ( p1_u3529,n18882 );
   nand U10428 ( n18882,n14516,n14517 );
   buf U10429 ( p1_u3530,n18883 );
   nand U10430 ( n18883,n14513,n14514 );
   buf U10431 ( p1_u3531,n18884 );
   nand U10432 ( n18884,n14510,n14511 );
   buf U10433 ( p1_u3532,n18885 );
   nand U10434 ( n18885,n14507,n14508 );
   buf U10435 ( p1_u3533,n18886 );
   nand U10436 ( n18886,n14504,n14505 );
   buf U10437 ( p1_u3534,n18887 );
   nand U10438 ( n18887,n14501,n14502 );
   buf U10439 ( p1_u3535,n18888 );
   nand U10440 ( n18888,n14498,n14499 );
   buf U10441 ( p1_u3536,n18889 );
   nand U10442 ( n18889,n14495,n14496 );
   buf U10443 ( p1_u3537,n18890 );
   nand U10444 ( n18890,n14492,n14493 );
   buf U10445 ( p1_u3538,n18891 );
   nand U10446 ( n18891,n14489,n14490 );
   buf U10447 ( p1_u3539,n18892 );
   nand U10448 ( n18892,n14486,n14487 );
   buf U10449 ( p1_u3540,n18893 );
   nand U10450 ( n18893,n14483,n14484 );
   buf U10451 ( p1_u3541,n18894 );
   nand U10452 ( n18894,n14480,n14481 );
   buf U10453 ( p1_u3542,n18895 );
   nand U10454 ( n18895,n14477,n14478 );
   buf U10455 ( p1_u3543,n18896 );
   nand U10456 ( n18896,n14474,n14475 );
   buf U10457 ( p1_u3544,n18897 );
   nand U10458 ( n18897,n14471,n14472 );
   buf U10459 ( p1_u3545,n18898 );
   nand U10460 ( n18898,n14468,n14469 );
   buf U10461 ( p1_u3546,n18899 );
   nand U10462 ( n18899,n14465,n14466 );
   buf U10463 ( p1_u3547,n18900 );
   nand U10464 ( n18900,n14462,n14463 );
   buf U10465 ( p1_u3548,n18901 );
   nand U10466 ( n18901,n14459,n14460 );
   buf U10467 ( p1_u3549,n18902 );
   nand U10468 ( n18902,n14456,n14457 );
   buf U10469 ( p1_u3550,n18903 );
   nand U10470 ( n18903,n14453,n14454 );
   buf U10471 ( p1_u3551,n18904 );
   nand U10472 ( n18904,n14450,n14451 );
   buf U10473 ( p1_u3552,n18905 );
   nand U10474 ( n18905,n14447,n14448 );
   buf U10475 ( p1_u3554,n18959 );
   nand U10476 ( n18959,n14439,n14440 );
   buf U10477 ( p1_u3555,n18960 );
   nand U10478 ( n18960,n14436,n14437 );
   buf U10479 ( p1_u3556,n18961 );
   nand U10480 ( n18961,n14433,n14434 );
   buf U10481 ( p1_u3557,n18962 );
   nand U10482 ( n18962,n14430,n14431 );
   buf U10483 ( p1_u3558,n18963 );
   nand U10484 ( n18963,n14427,n14428 );
   buf U10485 ( p1_u3559,n18964 );
   nand U10486 ( n18964,n14424,n14425 );
   buf U10487 ( p1_u3560,n18965 );
   nand U10488 ( n18965,n14421,n14422 );
   buf U10489 ( p1_u3561,n18966 );
   nand U10490 ( n18966,n14418,n14419 );
   buf U10491 ( p1_u3562,n18967 );
   nand U10492 ( n18967,n14415,n14416 );
   buf U10493 ( p1_u3563,n18968 );
   nand U10494 ( n18968,n14412,n14413 );
   buf U10495 ( p1_u3564,n18969 );
   nand U10496 ( n18969,n14409,n14410 );
   buf U10497 ( p1_u3565,n18970 );
   nand U10498 ( n18970,n14406,n14407 );
   buf U10499 ( p1_u3566,n18971 );
   nand U10500 ( n18971,n14403,n14404 );
   buf U10501 ( p1_u3567,n18972 );
   nand U10502 ( n18972,n14400,n14401 );
   buf U10503 ( p1_u3568,n18973 );
   nand U10504 ( n18973,n14397,n14398 );
   buf U10505 ( p1_u3569,n18974 );
   nand U10506 ( n18974,n14394,n14395 );
   buf U10507 ( p1_u3570,n18975 );
   nand U10508 ( n18975,n14391,n14392 );
   buf U10509 ( p1_u3571,n18976 );
   nand U10510 ( n18976,n14388,n14389 );
   buf U10511 ( p1_u3572,n18977 );
   nand U10512 ( n18977,n14385,n14386 );
   buf U10513 ( p1_u3573,n18978 );
   nand U10514 ( n18978,n14382,n14383 );
   buf U10515 ( p1_u3574,n18979 );
   nand U10516 ( n18979,n14379,n14380 );
   buf U10517 ( p1_u3575,n18980 );
   nand U10518 ( n18980,n14376,n14377 );
   buf U10519 ( p1_u3577,n18982 );
   nand U10520 ( n18982,n14370,n14371 );
   buf U10521 ( p1_u3578,n18983 );
   nand U10522 ( n18983,n14367,n14368 );
   buf U10523 ( p1_u3579,n18984 );
   nand U10524 ( n18984,n14364,n14365 );
   buf U10525 ( p1_u3580,n18985 );
   nand U10526 ( n18985,n14361,n14362 );
   buf U10527 ( p1_u3581,n18986 );
   nand U10528 ( n18986,n14358,n14359 );
   buf U10529 ( p1_u3582,n18987 );
   nand U10530 ( n18987,n14355,n14356 );
   buf U10531 ( p1_u3584,n18989 );
   nand U10532 ( n18989,n14349,n14350 );
   buf U10533 ( p1_u3585,n18990 );
   nand U10534 ( n18990,n14345,n14346 );
   buf U10535 ( p2_u3491,n19181 );
   nand U10536 ( n19181,n10548,n10549 );
   buf U10537 ( p2_u3492,n19182 );
   nand U10538 ( n19182,n10545,n10546 );
   buf U10539 ( p2_u3493,n19183 );
   nand U10540 ( n19183,n10542,n10543 );
   buf U10541 ( p2_u3494,n19184 );
   nand U10542 ( n19184,n10539,n10540 );
   buf U10543 ( p2_u3495,n19185 );
   nand U10544 ( n19185,n10536,n10537 );
   buf U10545 ( p2_u3496,n19186 );
   nand U10546 ( n19186,n10533,n10534 );
   buf U10547 ( p2_u3497,n19187 );
   nand U10548 ( n19187,n10530,n10531 );
   buf U10549 ( p2_u3498,n19188 );
   nand U10550 ( n19188,n10527,n10528 );
   buf U10551 ( p2_u3499,n19189 );
   nand U10552 ( n19189,n10524,n10525 );
   buf U10553 ( p2_u3500,n19190 );
   nand U10554 ( n19190,n10521,n10522 );
   buf U10555 ( p2_u3501,n19191 );
   nand U10556 ( n19191,n10518,n10519 );
   buf U10557 ( p2_u3502,n19192 );
   nand U10558 ( n19192,n10515,n10516 );
   buf U10559 ( p2_u3503,n19193 );
   nand U10560 ( n19193,n10512,n10513 );
   buf U10561 ( p2_u3504,n19194 );
   nand U10562 ( n19194,n10509,n10510 );
   buf U10563 ( p2_u3505,n19195 );
   nand U10564 ( n19195,n10506,n10507 );
   buf U10565 ( p2_u3506,n19196 );
   nand U10566 ( n19196,n10503,n10504 );
   buf U10567 ( p2_u3507,n19197 );
   nand U10568 ( n19197,n10500,n10501 );
   buf U10569 ( p2_u3508,n19198 );
   nand U10570 ( n19198,n10497,n10498 );
   buf U10571 ( p2_u3509,n19199 );
   nand U10572 ( n19199,n10494,n10495 );
   buf U10573 ( p2_u3510,n19200 );
   nand U10574 ( n19200,n10491,n10492 );
   buf U10575 ( p2_u3511,n19201 );
   nand U10576 ( n19201,n10488,n10489 );
   buf U10577 ( p2_u3513,n19203 );
   nand U10578 ( n19203,n10482,n10483 );
   buf U10579 ( p2_u3515,n19205 );
   nand U10580 ( n19205,n10476,n10477 );
   buf U10581 ( p2_u3516,n19206 );
   nand U10582 ( n19206,n10473,n10474 );
   buf U10583 ( p2_u3517,n19207 );
   nand U10584 ( n19207,n10470,n10471 );
   buf U10585 ( p2_u3518,n19208 );
   nand U10586 ( n19208,n10467,n10468 );
   buf U10587 ( p2_u3520,n19210 );
   nand U10588 ( n19210,n10461,n10462 );
   buf U10589 ( p2_u3521,n19211 );
   nand U10590 ( n19211,n10458,n10459 );
   buf U10591 ( p2_u3522,n19212 );
   nand U10592 ( n19212,n10454,n10455 );
   buf U10593 ( p2_u3185,n19177 );
   nand U10594 ( n19177,n13309,n13310,n13311 );
   nor U10595 ( n13311,n13312,n13313,n13314 );
   buf U10596 ( p1_u3279,n18921 );
   nand U10597 ( n18921,n15683,n15684,n15685,n15686 );
   nand U10598 ( n15683,n14996,n14766 );
   buf U10599 ( p1_u3265,n18935 );
   nand U10600 ( n18935,n16104,n16105,n16106,n16107 );
   nor U10601 ( n16107,n16108,n16109,n16110,n16111 );
   buf U10602 ( p1_u3269,n18931 );
   nand U10603 ( n18931,n15987,n15988,n15989,n15990 );
   buf U10604 ( p2_u3209,n19153 );
   nand U10605 ( n19153,n12379,n12380,n12381,n12382 );
   buf U10606 ( p1_u3293,n18907 );
   nand U10607 ( n18907,n15253,n15254,n15255,n15256 );
   nor U10608 ( n15256,n15257,n15258,n15259 );
   buf U10609 ( p1_u3216,n19017 );
   nand U10610 ( n19017,n17717,n17718,n17719,n17720 );
   buf U10611 ( p1_u3213,n19020 );
   nand U10612 ( n19020,n18328,n18329,n18330,n18331 );
   buf U10613 ( p2_u3213,n19149 );
   nand U10614 ( n19149,n12270,n12271,n12272,n12273 );
   nor U10615 ( n12273,n12274,n12275,n12276 );
   buf U10616 ( p2_u3211,n19151 );
   nand U10617 ( n19151,n12327,n12328,n12329,n12330 );
   nand U10618 ( n12327,n11837,n10771 );
   buf U10619 ( p2_u3154,n19241 );
   nand U10620 ( n19241,n13827,n13828,n13829,n13830 );
   buf U10621 ( p1_u3356,n18936 );
   nand U10622 ( n18936,n14979,n14980,n14981,n14982 );
   nand U10623 ( n14979,n14996,n14572 );
   buf U10624 ( p2_u3153,n19242 );
   nand U10625 ( n19242,n14137,n14138,n14139,n14140 );
   buf U10626 ( p2_u3204,n19158 );
   nand U10627 ( n19158,n12501,n12502,n12503,n12504 );
   nand U10628 ( n12501,n11837,n10685 );
   buf U10629 ( p1_u3247,n18954 );
   nand U10630 ( n18954,n16698,n16699,n16700,n16701 );
   buf U10631 ( add_1068_u4,n18777 );
   xor U10632 ( n18777,n18705,n18706 );
   nand U10633 ( n15437,n18359,n14966 );
   nand U10634 ( n16304,n16805,n16768 );
   nor U10635 ( n15300,n14929,n15302 );
   nor U10636 ( n15371,n14902,n15302 );
   nor U10637 ( n15928,n14669,n15302 );
   nor U10638 ( n15636,n14797,n15302 );
   nor U10639 ( n15689,n14773,n15302 );
   not U10640 ( n14991,n15302 );
   not U10641 ( n14551,n14607 );
   or U10642 ( n15030,n15031,n15032 );
   not U10643 ( n15031,n15061 );
   not U10644 ( n12701,n12745 );
   nand U10645 ( n12745,p2_u3893,n11164 );
   nand U10646 ( n14568,n14970,n16884 );
   not U10647 ( n11837,n11836 );
   nand U10648 ( n11836,n10650,n12668 );
   and U10649 ( n12525,n14271,n14270 );
   and U10650 ( n17284,n18547,n18546 );
   nand U10651 ( n11034,n10650,n9903 );
   nor U10652 ( n14287,n14291,n9903 );
   nor U10653 ( n14302,n14307,n9903 );
   nor U10654 ( n14301,n14308,n9903 );
   nor U10655 ( n14293,n14296,n9903 );
   nor U10656 ( n14304,n14305,n9903 );
   nor U10657 ( n14303,n14306,n9903 );
   nor U10658 ( n14297,n9903,n11819 );
   nor U10659 ( n14294,n9903,n11817 );
   nor U10660 ( n14300,n9903,n11822 );
   nor U10661 ( n14298,n9903,n11821 );
   nor U10662 ( n14289,n9903,n11816 );
   nor U10663 ( n14288,n9903,n11818 );
   nor U10664 ( n14290,n9903,n11814 );
   nor U10665 ( n14299,n9903,n11813 );
   nor U10666 ( n14295,n9903,n11820 );
   nor U10667 ( n14292,n9903,n11815 );
   or U10668 ( n14309,n9903,p2_d_reg_1_ );
   or U10669 ( n14312,n9903,p2_d_reg_0_ );
   nor U10670 ( n11550,n11812,p2_state_reg );
   not U10671 ( p1_u3973,n14347 );
   nand U10672 ( n14347,n16821,p1_state_reg,n16820 );
   not U10673 ( p2_u3893,n10456 );
   nand U10674 ( n10456,n11045,p2_state_reg,n13433 );
   nand U10675 ( n10727,n12646,n12499 );
   nor U10676 ( n12646,n12659,n13907 );
   nor U10677 ( n11546,n11808,p2_state_reg );
   nand U10678 ( n14622,n16187,n16188 );
   not U10679 ( n14545,n14553 );
   nand U10680 ( n14553,n14541,n14959,n14542 );
   not U10681 ( n14444,n14446 );
   nand U10682 ( n14446,n14540,n14541,n14542 );
   not U10683 ( n10553,n10555 );
   nand U10684 ( n10555,n10649,n10650,n10651,n10652 );
   nor U10685 ( n15029,n11808,p1_state_reg );
   nor U10686 ( n15033,n11812,p1_state_reg );
   nor U10687 ( n17294,n11812,n16273 );
   nor U10688 ( n17289,n11808,n16273 );
   nand U10689 ( n17657,n18536,n18537,n18538 );
   not U10690 ( n10670,n10671 );
   nand U10691 ( n10671,n11019,n11020 );
   nand U10692 ( n13751,n12594,n11163,n14255 );
   not U10693 ( n14996,n14995 );
   nand U10694 ( n14995,n14541,n16278 );
   not U10695 ( n11808,n11812 );
   nand U10696 ( n11812,n18593,n18594 );
   not U10697 ( n17654,n18185 );
   buf U10698 ( p2_u3150,n19243 );
   nand U10699 ( n19243,n13439,n14321 );
   buf U10700 ( p2_u3184,n19178 );
   nand U10701 ( n19178,n13351,n13352,n13353 );
   nor U10702 ( n13353,n13354,n13355,n13356 );
   buf U10703 ( p1_u3288,n18912 );
   nand U10704 ( n18912,n15378,n15379,n15380,n15381 );
   nor U10705 ( n15381,n15382,n15383,n15384,n15385 );
   buf U10706 ( p1_u3268,n18932 );
   nand U10707 ( n18932,n16006,n16007,n16008,n16009 );
   buf U10708 ( p2_u3208,n19154 );
   nand U10709 ( n19154,n12394,n12395,n12396,n12397 );
   buf U10710 ( p2_u3205,n19157 );
   nand U10711 ( n19157,n12474,n12475,n12476,n12477 );
   nor U10712 ( n12477,n12478,n12479,n12480 );
   buf U10713 ( p2_u3201,n19161 );
   nand U10714 ( n19161,n12679,n12680,n12681,n12682 );
   buf U10715 ( p2_u3155,n19240 );
   nand U10716 ( n19240,n13811,n13812,n13813,n13814 );
   buf U10717 ( p1_u3219,n19014 );
   nand U10718 ( n19014,n17679,n17680,n17681,n17682 );
   or U10719 ( n17680,n17686,n17351 );
   buf U10720 ( p2_u3182,n19180 );
   nand U10721 ( n19180,n13404,n13406,n13417,n13418 );
   buf U10722 ( p1_u3232,n19001 );
   nand U10723 ( n19001,n17472,n17473,n17474,n17475 );
   buf U10724 ( p2_u3172,n19223 );
   nand U10725 ( n19223,n13586,n13587,n13588,n13589 );
   nand U10726 ( n13589,p2_reg3_reg_0_,n13526 );
   buf U10727 ( add_1068_u55,n18778 );
   xor U10728 ( n18778,n18679,n18680 );
   buf U10729 ( add_1068_u56,n18779 );
   xor U10730 ( n18779,n18676,n18677 );
   buf U10731 ( add_1068_u57,n18780 );
   xor U10732 ( n18780,n18673,n18674 );
   buf U10733 ( add_1068_u58,n18781 );
   xor U10734 ( n18781,n18671,n18672 );
   buf U10735 ( add_1068_u59,n18782 );
   xor U10736 ( n18782,n18668,n18669 );
   buf U10737 ( add_1068_u60,n18783 );
   xor U10738 ( n18783,n18665,n18666 );
   buf U10739 ( add_1068_u61,n18784 );
   xor U10740 ( n18784,n18662,n18663 );
   buf U10741 ( add_1068_u62,n18785 );
   xor U10742 ( n18785,n18659,n18660 );
   buf U10743 ( add_1068_u63,n18786 );
   xor U10744 ( n18786,n18657,n18658 );
   buf U10745 ( add_1068_u47,n18787 );
   xor U10746 ( n18787,n18702,n18703 );
   buf U10747 ( add_1068_u48,n18788 );
   xor U10748 ( n18788,n18700,n18701 );
   buf U10749 ( add_1068_u49,n18789 );
   xor U10750 ( n18789,n18698,n18699 );
   buf U10751 ( add_1068_u50,n18790 );
   xor U10752 ( n18790,n18694,n18695 );
   buf U10753 ( add_1068_u51,n18791 );
   xor U10754 ( n18791,n18691,n18692 );
   buf U10755 ( add_1068_u52,n18792 );
   xor U10756 ( n18792,n18688,n18689 );
   buf U10757 ( add_1068_u53,n18793 );
   xor U10758 ( n18793,n18685,n18686 );
   buf U10759 ( add_1068_u54,n18794 );
   xor U10760 ( n18794,n18682,n18683 );
   buf U10761 ( add_1068_u5,n18795 );
   xor U10762 ( n18795,n18696,n18697 );
   xor U10763 ( n18697,p2_addr_reg_1_,p1_addr_reg_1_ );
   not U10764 ( n10453,p2_wr_reg );
   nand U10765 ( n10455,p2_datao_reg_31_,n10456 );
   nand U10766 ( n10454,p2_u3893,n10457 );
   nand U10767 ( n10459,p2_datao_reg_30_,n10456 );
   nand U10768 ( n10458,p2_u3893,n10460 );
   nand U10769 ( n10462,p2_datao_reg_29_,n10456 );
   nand U10770 ( n10461,p2_u3893,n10463 );
   nand U10771 ( n10465,p2_datao_reg_28_,n10456 );
   nand U10772 ( n10464,p2_u3893,n10466 );
   nand U10773 ( n10468,p2_datao_reg_27_,n10456 );
   nand U10774 ( n10467,p2_u3893,n10469 );
   nand U10775 ( n10471,p2_datao_reg_26_,n10456 );
   nand U10776 ( n10470,p2_u3893,n10472 );
   nand U10777 ( n10474,p2_datao_reg_25_,n10456 );
   nand U10778 ( n10473,p2_u3893,n10475 );
   nand U10779 ( n10477,p2_datao_reg_24_,n10456 );
   nand U10780 ( n10476,p2_u3893,n10478 );
   nand U10781 ( n10480,p2_datao_reg_23_,n10456 );
   nand U10782 ( n10479,p2_u3893,n10481 );
   nand U10783 ( n10483,p2_datao_reg_22_,n10456 );
   nand U10784 ( n10482,p2_u3893,n10484 );
   nand U10785 ( n10486,p2_datao_reg_21_,n10456 );
   nand U10786 ( n10485,p2_u3893,n10487 );
   nand U10787 ( n10489,p2_datao_reg_20_,n10456 );
   nand U10788 ( n10488,p2_u3893,n10490 );
   nand U10789 ( n10492,p2_datao_reg_19_,n10456 );
   nand U10790 ( n10491,p2_u3893,n10493 );
   nand U10791 ( n10495,p2_datao_reg_18_,n10456 );
   nand U10792 ( n10494,p2_u3893,n10496 );
   nand U10793 ( n10498,p2_datao_reg_17_,n10456 );
   nand U10794 ( n10497,p2_u3893,n10499 );
   nand U10795 ( n10501,p2_datao_reg_16_,n10456 );
   nand U10796 ( n10500,p2_u3893,n10502 );
   nand U10797 ( n10504,p2_datao_reg_15_,n10456 );
   nand U10798 ( n10503,p2_u3893,n10505 );
   nand U10799 ( n10507,p2_datao_reg_14_,n10456 );
   nand U10800 ( n10506,p2_u3893,n10508 );
   nand U10801 ( n10510,p2_datao_reg_13_,n10456 );
   nand U10802 ( n10509,p2_u3893,n10511 );
   nand U10803 ( n10513,p2_datao_reg_12_,n10456 );
   nand U10804 ( n10512,p2_u3893,n10514 );
   nand U10805 ( n10516,p2_datao_reg_11_,n10456 );
   nand U10806 ( n10515,p2_u3893,n10517 );
   nand U10807 ( n10519,p2_datao_reg_10_,n10456 );
   nand U10808 ( n10518,p2_u3893,n10520 );
   nand U10809 ( n10522,p2_datao_reg_9_,n10456 );
   nand U10810 ( n10521,p2_u3893,n10523 );
   nand U10811 ( n10525,p2_datao_reg_8_,n10456 );
   nand U10812 ( n10524,p2_u3893,n10526 );
   nand U10813 ( n10528,p2_datao_reg_7_,n10456 );
   nand U10814 ( n10527,p2_u3893,n10529 );
   nand U10815 ( n10531,p2_datao_reg_6_,n10456 );
   nand U10816 ( n10530,p2_u3893,n10532 );
   nand U10817 ( n10534,p2_datao_reg_5_,n10456 );
   nand U10818 ( n10533,p2_u3893,n10535 );
   nand U10819 ( n10537,p2_datao_reg_4_,n10456 );
   nand U10820 ( n10536,p2_u3893,n10538 );
   nand U10821 ( n10540,p2_datao_reg_3_,n10456 );
   nand U10822 ( n10539,p2_u3893,n10541 );
   nand U10823 ( n10543,p2_datao_reg_2_,n10456 );
   nand U10824 ( n10542,p2_u3893,n10544 );
   nand U10825 ( n10546,p2_datao_reg_1_,n10456 );
   nand U10826 ( n10545,p2_u3893,n10547 );
   nand U10827 ( n10549,p2_datao_reg_0_,n10456 );
   nand U10828 ( n10548,p2_u3893,n10550 );
   nand U10829 ( n10551,p2_reg1_reg_31_,n10555 );
   nand U10830 ( n10557,p2_reg1_reg_30_,n10555 );
   nand U10831 ( n10556,n10553,n10558 );
   nand U10832 ( n10560,p2_reg1_reg_29_,n10555 );
   nand U10833 ( n10559,n10553,n10561 );
   nand U10834 ( n10563,p2_reg1_reg_28_,n10555 );
   nand U10835 ( n10562,n10553,n10564 );
   nand U10836 ( n10566,p2_reg1_reg_27_,n10555 );
   nand U10837 ( n10565,n10553,n10567 );
   nand U10838 ( n10569,p2_reg1_reg_26_,n10555 );
   nand U10839 ( n10568,n10553,n10570 );
   nand U10840 ( n10572,p2_reg1_reg_25_,n10555 );
   nand U10841 ( n10571,n10553,n10573 );
   nand U10842 ( n10575,p2_reg1_reg_24_,n10555 );
   nand U10843 ( n10574,n10553,n10576 );
   nand U10844 ( n10578,p2_reg1_reg_23_,n10555 );
   nand U10845 ( n10577,n10553,n10579 );
   nand U10846 ( n10581,p2_reg1_reg_22_,n10555 );
   nand U10847 ( n10580,n10553,n10582 );
   nand U10848 ( n10584,p2_reg1_reg_21_,n10555 );
   nand U10849 ( n10583,n10553,n10585 );
   nand U10850 ( n10587,p2_reg1_reg_20_,n10555 );
   nand U10851 ( n10586,n10553,n10588 );
   nand U10852 ( n10590,p2_reg1_reg_19_,n10555 );
   nand U10853 ( n10589,n10553,n10591 );
   nand U10854 ( n10593,p2_reg1_reg_18_,n10555 );
   nand U10855 ( n10592,n10553,n10594 );
   nand U10856 ( n10596,p2_reg1_reg_17_,n10555 );
   nand U10857 ( n10595,n10553,n10597 );
   nand U10858 ( n10599,p2_reg1_reg_16_,n10555 );
   nand U10859 ( n10598,n10553,n10600 );
   nand U10860 ( n10602,p2_reg1_reg_15_,n10555 );
   nand U10861 ( n10601,n10553,n10603 );
   nand U10862 ( n10605,p2_reg1_reg_14_,n10555 );
   nand U10863 ( n10604,n10553,n10606 );
   nand U10864 ( n10608,p2_reg1_reg_13_,n10555 );
   nand U10865 ( n10607,n10553,n10609 );
   nand U10866 ( n10611,p2_reg1_reg_12_,n10555 );
   nand U10867 ( n10610,n10553,n10612 );
   nand U10868 ( n10614,p2_reg1_reg_11_,n10555 );
   nand U10869 ( n10613,n10553,n10615 );
   nand U10870 ( n10617,p2_reg1_reg_10_,n10555 );
   nand U10871 ( n10616,n10553,n10618 );
   nand U10872 ( n10620,p2_reg1_reg_9_,n10555 );
   nand U10873 ( n10619,n10553,n10621 );
   nand U10874 ( n10623,p2_reg1_reg_8_,n10555 );
   nand U10875 ( n10622,n10553,n10624 );
   nand U10876 ( n10626,p2_reg1_reg_7_,n10555 );
   nand U10877 ( n10625,n10553,n10627 );
   nand U10878 ( n10629,p2_reg1_reg_6_,n10555 );
   nand U10879 ( n10628,n10553,n10630 );
   nand U10880 ( n10632,p2_reg1_reg_5_,n10555 );
   nand U10881 ( n10631,n10553,n10633 );
   nand U10882 ( n10635,p2_reg1_reg_4_,n10555 );
   nand U10883 ( n10634,n10553,n10636 );
   nand U10884 ( n10638,p2_reg1_reg_3_,n10555 );
   nand U10885 ( n10637,n10553,n10639 );
   nand U10886 ( n10641,p2_reg1_reg_2_,n10555 );
   nand U10887 ( n10640,n10553,n10642 );
   nand U10888 ( n10644,p2_reg1_reg_1_,n10555 );
   nand U10889 ( n10643,n10553,n10645 );
   nand U10890 ( n10647,p2_reg1_reg_0_,n10555 );
   nand U10891 ( n10646,n10553,n10648 );
   nand U10892 ( n10652,n10653,n10654 );
   nand U10893 ( n10654,n10655,n10656 );
   nand U10894 ( n10656,n10657,n10658,n10659 );
   nand U10895 ( n10658,n10660,n10661 );
   nand U10896 ( n10657,n10662,n10663 );
   nand U10897 ( n10651,n10664,n10665 );
   nand U10898 ( n10664,n10666,n10667 );
   nand U10899 ( n10669,n10670,p2_reg0_reg_31_ );
   nand U10900 ( n10668,n10671,n10554 );
   nand U10901 ( n10554,n10672,n10673 );
   nand U10902 ( n10673,n10674,n10675 );
   nand U10903 ( n10677,n10670,p2_reg0_reg_30_ );
   nand U10904 ( n10676,n10671,n10558 );
   nand U10905 ( n10558,n10672,n10678 );
   nand U10906 ( n10678,n10679,n10675 );
   nand U10907 ( n10681,n10670,p2_reg0_reg_29_ );
   nand U10908 ( n10680,n10671,n10561 );
   nand U10909 ( n10561,n10682,n10683,n10684 );
   not U10910 ( n10684,n10685 );
   nand U10911 ( n10683,n10686,n10687 );
   nand U10912 ( n10682,n10688,n10675 );
   nand U10913 ( n10690,n10670,p2_reg0_reg_28_ );
   nand U10914 ( n10689,n10671,n10564 );
   nand U10915 ( n10564,n10691,n10692,n10693,n10694 );
   nand U10916 ( n10694,n10695,n10686 );
   nand U10917 ( n10693,n10696,n10463 );
   nand U10918 ( n10692,n10697,n10675 );
   nand U10919 ( n10699,n10670,p2_reg0_reg_27_ );
   nand U10920 ( n10698,n10671,n10567 );
   nand U10921 ( n10567,n10700,n10701,n10702,n10703 );
   nand U10922 ( n10703,n10686,n10704 );
   nand U10923 ( n10702,n10696,n10466 );
   nand U10924 ( n10701,n10705,n10675 );
   nand U10925 ( n10707,n10670,p2_reg0_reg_26_ );
   nand U10926 ( n10706,n10671,n10570 );
   nand U10927 ( n10570,n10708,n10709,n10710,n10711 );
   or U10928 ( n10711,n10712,n10713,n10714 );
   nand U10929 ( n10710,n10696,n10469 );
   nand U10930 ( n10709,n10715,n10675 );
   not U10931 ( n10708,n10716 );
   nand U10932 ( n10718,n10670,p2_reg0_reg_25_ );
   nand U10933 ( n10717,n10671,n10573 );
   nand U10934 ( n10573,n10719,n10720,n10721,n10722 );
   nor U10935 ( n10722,n10723,n10724,n10725 );
   nor U10936 ( n10725,n10726,n10727 );
   nor U10937 ( n10724,n10728,n10729 );
   nor U10938 ( n10723,n10730,n10731 );
   nand U10939 ( n10721,n10732,n10733 );
   or U10940 ( n10720,n10734,n10714 );
   or U10941 ( n10719,n10734,n10735 );
   nand U10942 ( n10737,n10670,p2_reg0_reg_24_ );
   nand U10943 ( n10736,n10671,n10576 );
   nand U10944 ( n10576,n10738,n10739,n10740,n10741 );
   nor U10945 ( n10741,n10742,n10743,n10744 );
   nor U10946 ( n10744,n10745,n10727 );
   nor U10947 ( n10743,n10746,n10729 );
   nor U10948 ( n10742,n10730,n10747 );
   nand U10949 ( n10740,n10748,n10733 );
   or U10950 ( n10739,n10714,n10749 );
   or U10951 ( n10738,n10749,n10735 );
   nand U10952 ( n10751,n10670,p2_reg0_reg_23_ );
   nand U10953 ( n10750,n10671,n10579 );
   nand U10954 ( n10579,n10752,n10753,n10754,n10755 );
   nor U10955 ( n10755,n10756,n10757,n10758 );
   nor U10956 ( n10758,n10759,n10727 );
   nor U10957 ( n10757,n10726,n10729 );
   nor U10958 ( n10756,n10730,n10760 );
   nand U10959 ( n10754,n10686,n10761 );
   nand U10960 ( n10752,n10762,n10733 );
   nand U10961 ( n10764,n10670,p2_reg0_reg_22_ );
   nand U10962 ( n10763,n10671,n10582 );
   nand U10963 ( n10582,n10765,n10766,n10767,n10768 );
   nand U10964 ( n10768,n10686,n10769 );
   nand U10965 ( n10767,n10696,n10481 );
   nand U10966 ( n10766,n10770,n10675 );
   not U10967 ( n10765,n10771 );
   nand U10968 ( n10773,n10670,p2_reg0_reg_21_ );
   nand U10969 ( n10772,n10671,n10585 );
   nand U10970 ( n10585,n10774,n10775,n10776,n10777 );
   nor U10971 ( n10777,n10778,n10779 );
   nor U10972 ( n10778,n10730,n10780 );
   nand U10973 ( n10776,n10781,n10490 );
   nand U10974 ( n10775,n10782,n10686 );
   nand U10975 ( n10774,n10696,n10484 );
   nand U10976 ( n10784,n10670,p2_reg0_reg_20_ );
   nand U10977 ( n10783,n10671,n10588 );
   nand U10978 ( n10588,n10785,n10786,n10787,n10788 );
   nand U10979 ( n10788,n10789,n10686 );
   nand U10980 ( n10787,n10696,n10487 );
   nand U10981 ( n10786,n10790,n10675 );
   nand U10982 ( n10792,n10670,p2_reg0_reg_19_ );
   nand U10983 ( n10791,n10671,n10591 );
   nand U10984 ( n10591,n10793,n10794,n10795,n10796 );
   nand U10985 ( n10796,n10797,n10686 );
   nand U10986 ( n10795,n10696,n10490 );
   nand U10987 ( n10794,n10798,n10675 );
   nand U10988 ( n10800,n10670,p2_reg0_reg_18_ );
   nand U10989 ( n10799,n10671,n10594 );
   nand U10990 ( n10594,n10801,n10802,n10803,n10804 );
   nor U10991 ( n10804,n10805,n10806 );
   nor U10992 ( n10806,n10730,n10807 );
   nor U10993 ( n10805,n10808,n10727 );
   nand U10994 ( n10803,n10696,n10493 );
   nand U10995 ( n10802,n10809,n10810 );
   or U10996 ( n10801,n10811,n10812 );
   nand U10997 ( n10814,n10670,p2_reg0_reg_17_ );
   nand U10998 ( n10813,n10671,n10597 );
   nand U10999 ( n10597,n10815,n10816,n10817,n10818 );
   nor U11000 ( n10818,n10819,n10820 );
   nor U11001 ( n10820,n10730,n10821 );
   nor U11002 ( n10819,n10822,n10727 );
   nand U11003 ( n10817,n10696,n10496 );
   or U11004 ( n10816,n10823,n10812,n10824 );
   nand U11005 ( n10815,n10825,n10810 );
   nand U11006 ( n10827,n10670,p2_reg0_reg_16_ );
   nand U11007 ( n10826,n10671,n10600 );
   nand U11008 ( n10600,n10828,n10829,n10830,n10831 );
   nor U11009 ( n10831,n10832,n10833 );
   nor U11010 ( n10833,n10730,n10834 );
   nor U11011 ( n10832,n10835,n10727 );
   nand U11012 ( n10830,n10696,n10499 );
   nand U11013 ( n10828,n10836,n10810 );
   nand U11014 ( n10838,n10670,p2_reg0_reg_15_ );
   nand U11015 ( n10837,n10671,n10603 );
   nand U11016 ( n10603,n10839,n10840,n10841,n10842 );
   nand U11017 ( n10842,n10843,n10686 );
   nand U11018 ( n10841,n10696,n10502 );
   nand U11019 ( n10840,n10844,n10675 );
   nand U11020 ( n10846,n10670,p2_reg0_reg_14_ );
   nand U11021 ( n10845,n10671,n10606 );
   nand U11022 ( n10606,n10847,n10848,n10849,n10850 );
   or U11023 ( n10850,n10851,n10714 );
   nand U11024 ( n10849,n10696,n10505 );
   nand U11025 ( n10848,n10852,n10675 );
   not U11026 ( n10847,n10853 );
   nand U11027 ( n10855,n10670,p2_reg0_reg_13_ );
   nand U11028 ( n10854,n10671,n10609 );
   nand U11029 ( n10609,n10856,n10857,n10858,n10859 );
   nand U11030 ( n10859,n10860,n10686 );
   nand U11031 ( n10858,n10696,n10508 );
   nand U11032 ( n10857,n10861,n10675 );
   not U11033 ( n10856,n10862 );
   nand U11034 ( n10864,n10670,p2_reg0_reg_12_ );
   nand U11035 ( n10863,n10671,n10612 );
   nand U11036 ( n10612,n10865,n10866,n10867,n10868 );
   nor U11037 ( n10868,n10869,n10870,n10871 );
   nor U11038 ( n10871,n10872,n10727 );
   nor U11039 ( n10870,n10873,n10729 );
   nor U11040 ( n10869,n10730,n10874 );
   nand U11041 ( n10867,n10875,n10733 );
   nand U11042 ( n10865,n10876,n10877 );
   nand U11043 ( n10879,n10670,p2_reg0_reg_11_ );
   nand U11044 ( n10878,n10671,n10615 );
   nand U11045 ( n10615,n10880,n10881,n10882,n10883 );
   nor U11046 ( n10883,n10884,n10885,n10886 );
   nor U11047 ( n10886,n10887,n10727 );
   nor U11048 ( n10885,n10888,n10729 );
   nor U11049 ( n10884,n10730,n10889 );
   or U11050 ( n10882,n10890,n10812 );
   nand U11051 ( n10880,n10891,n10877 );
   nand U11052 ( n10893,n10670,p2_reg0_reg_10_ );
   nand U11053 ( n10892,n10671,n10618 );
   nand U11054 ( n10618,n10894,n10895,n10896,n10897 );
   nor U11055 ( n10897,n10898,n10899 );
   nor U11056 ( n10899,n10730,n10900 );
   nor U11057 ( n10898,n10901,n10727 );
   nand U11058 ( n10896,n10696,n10517 );
   nand U11059 ( n10895,n10902,n10903,n10733 );
   nand U11060 ( n10894,n10904,n10810 );
   nand U11061 ( n10906,n10670,p2_reg0_reg_9_ );
   nand U11062 ( n10905,n10671,n10621 );
   nand U11063 ( n10621,n10907,n10908,n10909,n10910 );
   nor U11064 ( n10910,n10911,n10912 );
   nor U11065 ( n10912,n10730,n10913 );
   nor U11066 ( n10911,n10914,n10727 );
   nand U11067 ( n10909,n10696,n10520 );
   nand U11068 ( n10908,n10915,n10810 );
   or U11069 ( n10907,n10916,n10812 );
   nand U11070 ( n10918,n10670,p2_reg0_reg_8_ );
   nand U11071 ( n10917,n10671,n10624 );
   nand U11072 ( n10624,n10919,n10920,n10921,n10922 );
   nand U11073 ( n10922,n10686,n10923 );
   nand U11074 ( n10921,n10696,n10523 );
   nand U11075 ( n10920,n10924,n10675 );
   not U11076 ( n10919,n10925 );
   nand U11077 ( n10927,n10670,p2_reg0_reg_7_ );
   nand U11078 ( n10926,n10671,n10627 );
   nand U11079 ( n10627,n10928,n10929,n10930,n10931 );
   nor U11080 ( n10931,n10932,n10933,n10934 );
   nor U11081 ( n10934,n10935,n10727 );
   nor U11082 ( n10933,n10914,n10729 );
   nor U11083 ( n10932,n10730,n10936 );
   nand U11084 ( n10930,n10937,n10877 );
   nand U11085 ( n10928,n10938,n10733,n10939 );
   nand U11086 ( n10941,n10670,p2_reg0_reg_6_ );
   nand U11087 ( n10940,n10671,n10630 );
   nand U11088 ( n10630,n10942,n10943,n10944,n10945 );
   nand U11089 ( n10945,n10686,n10946 );
   nand U11090 ( n10944,n10696,n10529 );
   nand U11091 ( n10943,n10947,n10675 );
   not U11092 ( n10942,n10948 );
   nand U11093 ( n10950,n10670,p2_reg0_reg_5_ );
   nand U11094 ( n10949,n10671,n10633 );
   nand U11095 ( n10633,n10951,n10952,n10953,n10954 );
   nor U11096 ( n10954,n10955,n10956 );
   nor U11097 ( n10956,n10730,n10957 );
   nor U11098 ( n10955,n10958,n10727 );
   nand U11099 ( n10953,n10696,n10532 );
   nand U11100 ( n10952,n10959,n10960,n10733 );
   nand U11101 ( n10951,n10961,n10810 );
   nand U11102 ( n10963,n10670,p2_reg0_reg_4_ );
   nand U11103 ( n10962,n10671,n10636 );
   nand U11104 ( n10636,n10964,n10965,n10966,n10967 );
   nor U11105 ( n10967,n10968,n10969 );
   nor U11106 ( n10969,n10730,n10970 );
   nor U11107 ( n10968,n10971,n10727 );
   nand U11108 ( n10966,n10696,n10535 );
   nand U11109 ( n10965,n10972,n10810 );
   or U11110 ( n10964,n10973,n10812 );
   nand U11111 ( n10974,n10671,n10639 );
   nand U11112 ( n10639,n10976,n10977,n10978,n10979 );
   nor U11113 ( n10979,n10980,n10981,n10982 );
   nor U11114 ( n10982,n10983,n10727 );
   nor U11115 ( n10981,n10958,n10729 );
   nor U11116 ( n10980,n10730,n10984 );
   nand U11117 ( n10978,n10985,n10733 );
   nand U11118 ( n10976,n10877,n10986 );
   nand U11119 ( n10877,n10987,n10714 );
   nand U11120 ( n10988,n10671,n10642 );
   nand U11121 ( n10642,n10990,n10991,n10992,n10993 );
   nand U11122 ( n10993,n10994,n10686 );
   nand U11123 ( n10992,n10696,n10541 );
   nand U11124 ( n10991,n10995,n10675 );
   not U11125 ( n10990,n10996 );
   nand U11126 ( n10997,n10671,n10645 );
   nand U11127 ( n10645,n10999,n11000,n11001,n11002 );
   nor U11128 ( n11002,n11003,n11004 );
   nor U11129 ( n11004,n10730,n11005 );
   nor U11130 ( n11003,n11006,n10727 );
   nand U11131 ( n11001,n10696,n10544 );
   nand U11132 ( n11000,n11007,n10810 );
   nand U11133 ( n10810,n10735,n10714 );
   not U11134 ( n10735,n11008 );
   nand U11135 ( n10999,n11009,n10733 );
   nand U11136 ( n10648,n11012,n11013,n11014,n11015 );
   nand U11137 ( n11015,n10686,n11016 );
   nand U11138 ( n11014,n10696,n10547 );
   nand U11139 ( n11013,n11017,n10675 );
   not U11140 ( n11012,n11018 );
   nand U11141 ( n11020,n10650,n11021 );
   nand U11142 ( n11021,n11022,n11023 );
   nand U11143 ( n11023,n11024,n11025 );
   nand U11144 ( n11022,n11026,n11027 );
   nand U11145 ( n11027,n11028,n11029 );
   nand U11146 ( n11029,n10662,n11030 );
   xor U11147 ( n11028,n10660,n10661 );
   nand U11148 ( n11019,n11031,n11025 );
   nand U11149 ( n11033,p2_d_reg_1_,n11034 );
   nand U11150 ( n11032,n11035,n11036 );
   nand U11151 ( n11038,p2_d_reg_0_,n11034 );
   nand U11152 ( n11037,n11035,n11039 );
   nor U11153 ( n11041,n11042,n11043 );
   not U11154 ( n11043,n11044 );
   nor U11155 ( n11042,p2_u3151,n11045 );
   nor U11156 ( n11048,n11049,n11050 );
   and U11157 ( n11047,n11050,n11051 );
   nand U11158 ( n11050,n11052,n11053 );
   nand U11159 ( n11053,n11054,n11055 );
   nand U11160 ( n11055,n11056,n11057 );
   nand U11161 ( n11057,n11058,n10674 );
   or U11162 ( n11058,n11059,n10460 );
   or U11163 ( n11056,n10457,n10679 );
   nand U11164 ( n11054,n11060,n11061 );
   nand U11165 ( n11061,n11062,n11063 );
   or U11166 ( n11063,n11064,n10463 );
   nand U11167 ( n11062,n11065,n11066 );
   nand U11168 ( n11066,n11067,n11068 );
   nand U11169 ( n11067,n11069,n11070 );
   nand U11170 ( n11070,n11071,n11072,n11073,n11074 );
   nor U11171 ( n11074,n11075,n11076 );
   nor U11172 ( n11076,n11077,n11078,n11079 );
   not U11173 ( n11079,n11080 );
   nor U11174 ( n11078,n11081,n11082 );
   nor U11175 ( n11082,n11083,n11084 );
   nor U11176 ( n11083,n11085,n11086 );
   not U11177 ( n11085,n11087 );
   nand U11178 ( n11077,n11088,n11089,n11090 );
   nand U11179 ( n11090,n11091,n11087,n11092,n11093 );
   nor U11180 ( n11093,n11094,n11081,n11095 );
   not U11181 ( n11095,n11096 );
   nand U11182 ( n11092,n11097,n11098,n11099 );
   nand U11183 ( n11099,n11100,n11101 );
   nand U11184 ( n11101,n11102,n11103,n11104 );
   nand U11185 ( n11102,n11105,n11106 );
   nand U11186 ( n11105,n11107,n11108 );
   nand U11187 ( n11108,n11109,n11110,n11111,n11112 );
   nor U11188 ( n11112,n11113,n11114,n11115 );
   nor U11189 ( n11115,n11116,n10511 );
   nor U11190 ( n11114,n11117,n11118,n11119 );
   nor U11191 ( n11113,n11118,n11120 );
   nand U11192 ( n11109,n11121,n11122,n11123,n11124 );
   nor U11193 ( n11124,n11118,n11125,n11119,n11126 );
   nor U11194 ( n11126,n11127,n11128,n11129,n11130 );
   nand U11195 ( n11128,n11131,n11132 );
   nand U11196 ( n11131,n10971,n11133 );
   not U11197 ( n11119,n11134 );
   nor U11198 ( n11125,n11135,n11130 );
   nor U11199 ( n11135,n11136,n11137 );
   nor U11200 ( n11136,n10914,n10924 );
   not U11201 ( n11118,n11138 );
   nand U11202 ( n11122,n11139,n11140,n11141 );
   nor U11203 ( n11141,n11127,n10971,n11133 );
   nand U11204 ( n11121,n11140,n11142,n11139 );
   nand U11205 ( n11142,n11143,n11144,n11145 );
   nand U11206 ( n11097,n10807,n10496 );
   nand U11207 ( n11091,n11146,n11098,n11147 );
   nand U11208 ( n11073,n11088,n11089,n11148 );
   nand U11209 ( n11148,n11149,n11150 );
   nand U11210 ( n11060,n11064,n10463 );
   nand U11211 ( n11052,n11151,n10674 );
   nand U11212 ( n11151,n10457,n11152 );
   nand U11213 ( n11152,n11059,n10460 );
   nand U11214 ( n11046,n11153,n11154,n11044 );
   nand U11215 ( n11044,p2_b_reg,n11155 );
   nand U11216 ( n11155,n11156,n11157,p2_state_reg );
   nand U11217 ( n11157,n11158,n11045 );
   nand U11218 ( n11158,n11159,n11160,n11161,n11162 );
   nor U11219 ( n11162,n11163,n11164 );
   nand U11220 ( n11156,n11165,n11166 );
   nand U11221 ( n11154,n11167,n11168 );
   xor U11222 ( n11167,n11169,n11170 );
   nand U11223 ( n11170,n11171,n11172,n11173,n11174 );
   nand U11224 ( n11174,n11175,n11176,n11177 );
   nand U11225 ( n11173,n11178,n11179,n11180 );
   nand U11226 ( n11172,n11181,n11182,n11178 );
   and U11227 ( n11178,n11175,n11183 );
   or U11228 ( n11183,n11176,n11177 );
   and U11229 ( n11177,n11184,n11185 );
   nand U11230 ( n11185,n10679,n11186 );
   nand U11231 ( n11184,n11187,n10460 );
   nand U11232 ( n11176,n11188,n11189 );
   nand U11233 ( n11189,n11186,n10460 );
   nand U11234 ( n11188,n10679,n11187 );
   nand U11235 ( n11175,n11190,n11191 );
   or U11236 ( n11182,n11179,n11180 );
   and U11237 ( n11180,n11192,n11193 );
   nand U11238 ( n11193,n10688,n11186 );
   nand U11239 ( n11192,n11187,n10463 );
   nand U11240 ( n11179,n11194,n11195 );
   nand U11241 ( n11195,n11186,n10463 );
   nand U11242 ( n11194,n10688,n11187 );
   nand U11243 ( n11181,n11196,n11197,n11198 );
   nand U11244 ( n11198,n11199,n11200,n11201,n11202 );
   nand U11245 ( n11201,n11203,n11204 );
   or U11246 ( n11200,n11205,n11206 );
   nand U11247 ( n11199,n11207,n11208,n11209 );
   or U11248 ( n11209,n11204,n11203 );
   and U11249 ( n11203,n11210,n11211 );
   nand U11250 ( n11211,n11186,n10472 );
   nand U11251 ( n11210,n10715,n11187 );
   nand U11252 ( n11204,n11212,n11213 );
   nand U11253 ( n11213,n10715,n11186 );
   nand U11254 ( n11212,n11187,n10472 );
   nand U11255 ( n11208,n11214,n11215,n11216,n11217 );
   nand U11256 ( n11217,n11218,n11219 );
   nand U11257 ( n11216,n11220,n11221,n11222,n11223 );
   nor U11258 ( n11223,n11224,n11225,n11226,n11227 );
   nor U11259 ( n11227,n11228,n11229 );
   nor U11260 ( n11226,n11230,n11231,n11232 );
   not U11261 ( n11231,n11233 );
   nor U11262 ( n11225,n11234,n11235,n11236 );
   nand U11263 ( n11222,n11237,n11238,n11239 );
   nor U11264 ( n11239,n11240,n11241,n11242 );
   nor U11265 ( n11242,n11243,n11244 );
   nor U11266 ( n11244,n11245,n11246 );
   nor U11267 ( n11246,n11247,n11248 );
   and U11268 ( n11245,n11249,n11250 );
   nor U11269 ( n11241,n11243,n11251,n11252,n11253 );
   not U11270 ( n11243,n11254 );
   and U11271 ( n11240,n11236,n11235 );
   and U11272 ( n11235,n11255,n11256 );
   nand U11273 ( n11256,n11186,n10493 );
   nand U11274 ( n11255,n10798,n11187 );
   nand U11275 ( n11236,n11257,n11258 );
   nand U11276 ( n11258,n10798,n11186 );
   nand U11277 ( n11257,n11187,n10493 );
   nand U11278 ( n11238,n11259,n11254,n11260,n11261 );
   nor U11279 ( n11261,n11252,n11262 );
   and U11280 ( n11262,n11253,n11251 );
   and U11281 ( n11251,n11263,n11264 );
   nand U11282 ( n11264,n11265,n11186 );
   nand U11283 ( n11263,n11187,n10502 );
   nand U11284 ( n11253,n11266,n11267 );
   nand U11285 ( n11267,n11186,n10502 );
   nand U11286 ( n11266,n11265,n11187 );
   nor U11287 ( n11252,n11250,n11249 );
   nand U11288 ( n11249,n11268,n11269 );
   nand U11289 ( n11269,n11270,n11186 );
   nand U11290 ( n11268,n11187,n10499 );
   and U11291 ( n11250,n11271,n11272 );
   nand U11292 ( n11272,n11186,n10499 );
   nand U11293 ( n11271,n11270,n11187 );
   nand U11294 ( n11260,n11273,n11274 );
   nand U11295 ( n11254,n11247,n11248 );
   nand U11296 ( n11248,n11275,n11276 );
   nand U11297 ( n11276,n11186,n10496 );
   nand U11298 ( n11275,n11147,n11187 );
   and U11299 ( n11247,n11277,n11278 );
   nand U11300 ( n11278,n11147,n11186 );
   nand U11301 ( n11277,n11187,n10496 );
   nand U11302 ( n11259,n11279,n11280 );
   nand U11303 ( n11280,n11281,n11282 );
   nand U11304 ( n11282,n11186,n10505 );
   nand U11305 ( n11281,n10844,n11187 );
   or U11306 ( n11279,n11274,n11273 );
   and U11307 ( n11273,n11283,n11284 );
   nand U11308 ( n11284,n10844,n11186 );
   nand U11309 ( n11283,n11187,n10505 );
   nand U11310 ( n11274,n11285,n11286 );
   nand U11311 ( n11286,n11287,n11288 );
   nand U11312 ( n11288,n11289,n11290 );
   nand U11313 ( n11287,n11291,n11292 );
   nand U11314 ( n11292,n11186,n10508 );
   nand U11315 ( n11291,n11187,n10852 );
   or U11316 ( n11285,n11290,n11289 );
   and U11317 ( n11289,n11293,n11294 );
   nand U11318 ( n11294,n11295,n11296,n11297,n11298 );
   nor U11319 ( n11298,n11299,n11300 );
   nor U11320 ( n11300,n11301,n11302 );
   nor U11321 ( n11299,n11303,n11304 );
   nand U11322 ( n11297,n11305,n11306,n11307 );
   nand U11323 ( n11296,n11308,n11309,n11310,n11311 );
   nor U11324 ( n11311,n11312,n11313 );
   nor U11325 ( n11312,n11314,n11315 );
   nand U11326 ( n11310,n11316,n11317 );
   nand U11327 ( n11309,n11318,n11319 );
   not U11328 ( n11319,n11320 );
   nand U11329 ( n11318,n11321,n11322 );
   nand U11330 ( n11322,n11323,n11324,n11325 );
   not U11331 ( n11324,n11326 );
   nand U11332 ( n11321,n11327,n11328 );
   nand U11333 ( n11308,n11329,n11330,n11331,n11332 );
   nor U11334 ( n11332,n11333,n11320,n11326 );
   nor U11335 ( n11326,n11328,n11327 );
   and U11336 ( n11327,n11334,n11335 );
   nand U11337 ( n11335,n10924,n11186 );
   nand U11338 ( n11334,n11187,n10526 );
   nand U11339 ( n11328,n11336,n11337 );
   nand U11340 ( n11337,n11186,n10526 );
   nand U11341 ( n11336,n10924,n11187 );
   nor U11342 ( n11320,n11317,n11316 );
   and U11343 ( n11316,n11338,n11339 );
   nand U11344 ( n11339,n11340,n11186 );
   nand U11345 ( n11338,n11187,n10523 );
   nand U11346 ( n11317,n11341,n11342 );
   nand U11347 ( n11342,n11186,n10523 );
   nand U11348 ( n11341,n11340,n11187 );
   nor U11349 ( n11333,n11343,n11344,n11345 );
   nand U11350 ( n11331,n11346,n11347,n11348,n11349 );
   nand U11351 ( n11349,n11350,n11351 );
   nand U11352 ( n11351,n11352,n11353 );
   nand U11353 ( n11350,n11354,n11355 );
   nand U11354 ( n11355,n11356,n11357 );
   nand U11355 ( n11357,n11358,n11359 );
   nand U11356 ( n11356,n11360,n11361 );
   nand U11357 ( n11361,n11186,n10544 );
   nand U11358 ( n11360,n10995,n11187 );
   or U11359 ( n11354,n11359,n11358 );
   and U11360 ( n11358,n11362,n11363 );
   nand U11361 ( n11363,n11364,n11365,n11366 );
   or U11362 ( n11366,n11367,n11368 );
   nand U11363 ( n11365,n11369,n11370 );
   nand U11364 ( n11370,n11368,n11367 );
   nand U11365 ( n11367,n11371,n11372 );
   nand U11366 ( n11372,n11186,n10550 );
   nand U11367 ( n11371,n11187,n11017 );
   nand U11368 ( n11369,n11373,n11374 );
   nand U11369 ( n11374,n11187,n10550 );
   nand U11370 ( n11364,n11375,n11376 );
   or U11371 ( n11362,n11376,n11375 );
   and U11372 ( n11375,n11377,n11378 );
   nand U11373 ( n11378,n10547,n11186 );
   nand U11374 ( n11377,n11379,n11187 );
   nand U11375 ( n11376,n11380,n11381 );
   nand U11376 ( n11381,n11186,n11379 );
   nand U11377 ( n11380,n11187,n10547 );
   nand U11378 ( n11359,n11382,n11383 );
   nand U11379 ( n11383,n10995,n11186 );
   nand U11380 ( n11382,n11187,n10544 );
   nand U11381 ( n11348,n11344,n11345 );
   nand U11382 ( n11345,n11384,n11385 );
   nand U11383 ( n11385,n11186,n10538 );
   nand U11384 ( n11384,n11386,n11187 );
   and U11385 ( n11344,n11387,n11388 );
   nand U11386 ( n11388,n11386,n11186 );
   nand U11387 ( n11387,n11187,n10538 );
   or U11388 ( n11347,n11353,n11352 );
   and U11389 ( n11352,n11389,n11390 );
   nand U11390 ( n11390,n10541,n11186 );
   nand U11391 ( n11389,n11133,n11187 );
   nand U11392 ( n11353,n11391,n11392 );
   nand U11393 ( n11392,n11186,n11133 );
   nand U11394 ( n11391,n11187,n10541 );
   not U11395 ( n11346,n11343 );
   nand U11396 ( n11343,n11393,n11394 );
   nand U11397 ( n11394,n11395,n11396 );
   nand U11398 ( n11330,n11397,n11393 );
   nand U11399 ( n11393,n11398,n11399 );
   nand U11400 ( n11397,n11400,n11401 );
   or U11401 ( n11401,n11396,n11395 );
   and U11402 ( n11395,n11402,n11403 );
   nand U11403 ( n11403,n11404,n11186 );
   nand U11404 ( n11402,n11187,n10535 );
   nand U11405 ( n11396,n11405,n11406 );
   nand U11406 ( n11406,n11186,n10535 );
   nand U11407 ( n11405,n11404,n11187 );
   or U11408 ( n11400,n11399,n11398 );
   and U11409 ( n11398,n11407,n11408 );
   nand U11410 ( n11408,n11186,n10947 );
   nand U11411 ( n11407,n11187,n10532 );
   nand U11412 ( n11399,n11409,n11410 );
   nand U11413 ( n11410,n11186,n10532 );
   nand U11414 ( n11409,n11187,n10947 );
   or U11415 ( n11329,n11323,n11325 );
   and U11416 ( n11325,n11411,n11412 );
   nand U11417 ( n11412,n11413,n11186 );
   nand U11418 ( n11411,n11187,n10529 );
   nand U11419 ( n11323,n11414,n11415 );
   nand U11420 ( n11415,n11186,n10529 );
   nand U11421 ( n11414,n11413,n11187 );
   nand U11422 ( n11295,n11416,n11315,n11314 );
   and U11423 ( n11314,n11417,n11418 );
   nand U11424 ( n11418,n11186,n10520 );
   nand U11425 ( n11417,n11187,n11419 );
   nand U11426 ( n11315,n11420,n11421 );
   nand U11427 ( n11421,n11186,n11419 );
   nand U11428 ( n11420,n11187,n10520 );
   not U11429 ( n11416,n11313 );
   nand U11430 ( n11313,n11422,n11306 );
   nand U11431 ( n11306,n11303,n11304 );
   nand U11432 ( n11304,n11423,n11424 );
   nand U11433 ( n11424,n11186,n10514 );
   nand U11434 ( n11423,n11425,n11187 );
   and U11435 ( n11303,n11426,n11427 );
   nand U11436 ( n11427,n11425,n11186 );
   nand U11437 ( n11426,n11187,n10514 );
   or U11438 ( n11422,n11305,n11307 );
   and U11439 ( n11307,n11428,n11429 );
   nand U11440 ( n11429,n11186,n10517 );
   nand U11441 ( n11428,n11430,n11187 );
   nand U11442 ( n11305,n11431,n11432 );
   nand U11443 ( n11432,n11430,n11186 );
   nand U11444 ( n11431,n11187,n10517 );
   nand U11445 ( n11293,n11301,n11302 );
   nand U11446 ( n11302,n11433,n11434 );
   nand U11447 ( n11434,n10511,n11186 );
   nand U11448 ( n11433,n10861,n11187 );
   and U11449 ( n11301,n11435,n11436 );
   nand U11450 ( n11436,n11186,n10861 );
   nand U11451 ( n11435,n11187,n10511 );
   nand U11452 ( n11290,n11437,n11438 );
   nand U11453 ( n11438,n11186,n10852 );
   nand U11454 ( n11437,n11187,n10508 );
   not U11455 ( n11237,n11234 );
   nand U11456 ( n11234,n11439,n11233 );
   nand U11457 ( n11233,n11440,n11441 );
   nand U11458 ( n11439,n11232,n11230 );
   nand U11459 ( n11230,n11442,n11443 );
   nand U11460 ( n11443,n10790,n11186 );
   nand U11461 ( n11442,n11187,n10490 );
   and U11462 ( n11232,n11444,n11445 );
   nand U11463 ( n11445,n11186,n10490 );
   nand U11464 ( n11444,n10790,n11187 );
   or U11465 ( n11221,n11441,n11440 );
   and U11466 ( n11440,n11446,n11447 );
   nand U11467 ( n11447,n11186,n10487 );
   nand U11468 ( n11446,n11448,n11187 );
   nand U11469 ( n11441,n11449,n11450 );
   nand U11470 ( n11450,n11448,n11186 );
   nand U11471 ( n11449,n11187,n10487 );
   nand U11472 ( n11215,n11451,n11452 );
   nand U11473 ( n11214,n11453,n11454 );
   nand U11474 ( n11454,n11455,n11456 );
   nand U11475 ( n11456,n11220,n11229,n11228 );
   and U11476 ( n11228,n11457,n11458 );
   nand U11477 ( n11458,n11186,n10484 );
   nand U11478 ( n11457,n10770,n11187 );
   nand U11479 ( n11229,n11459,n11460 );
   nand U11480 ( n11460,n10770,n11186 );
   nand U11481 ( n11459,n11187,n10484 );
   nand U11482 ( n11220,n11461,n11462 );
   or U11483 ( n11455,n11462,n11461 );
   and U11484 ( n11461,n11463,n11464 );
   nand U11485 ( n11464,n11465,n11186 );
   nand U11486 ( n11463,n11187,n10481 );
   nand U11487 ( n11462,n11466,n11467 );
   nand U11488 ( n11467,n11186,n10481 );
   nand U11489 ( n11466,n11465,n11187 );
   not U11490 ( n11453,n11224 );
   nor U11491 ( n11224,n11219,n11218 );
   and U11492 ( n11218,n11468,n11469 );
   nand U11493 ( n11469,n11186,n10478 );
   nand U11494 ( n11468,n11470,n11187 );
   nand U11495 ( n11219,n11471,n11472 );
   nand U11496 ( n11472,n11470,n11186 );
   nand U11497 ( n11471,n11187,n10478 );
   or U11498 ( n11207,n11452,n11451 );
   and U11499 ( n11451,n11473,n11474 );
   nand U11500 ( n11474,n11186,n10475 );
   nand U11501 ( n11473,n11475,n11187 );
   nand U11502 ( n11452,n11476,n11477 );
   nand U11503 ( n11477,n11475,n11186 );
   nand U11504 ( n11476,n11187,n10475 );
   nand U11505 ( n11197,n11205,n11202,n11206 );
   and U11506 ( n11206,n11478,n11479 );
   nand U11507 ( n11479,n10705,n11186 );
   nand U11508 ( n11478,n11187,n10469 );
   nand U11509 ( n11202,n11480,n11481 );
   nand U11510 ( n11205,n11482,n11483 );
   nand U11511 ( n11483,n11186,n10469 );
   nand U11512 ( n11482,n10705,n11187 );
   or U11513 ( n11196,n11481,n11480 );
   and U11514 ( n11480,n11484,n11485 );
   nand U11515 ( n11485,n11186,n10466 );
   nand U11516 ( n11484,n10697,n11187 );
   nand U11517 ( n11481,n11486,n11487 );
   nand U11518 ( n11487,n10697,n11186 );
   nand U11519 ( n11486,n11187,n10466 );
   or U11520 ( n11171,n11191,n11190 );
   and U11521 ( n11190,n11488,n11489 );
   nand U11522 ( n11489,n11186,n10674 );
   nand U11523 ( n11488,n11187,n10457 );
   nand U11524 ( n11191,n11490,n11491 );
   nand U11525 ( n11491,n11186,n10457 );
   nand U11526 ( n11490,n11187,n10674 );
   nand U11527 ( n11494,n11161,n11492 );
   nand U11528 ( n11169,n11493,n11495 );
   nand U11529 ( n11495,n10662,n11496 );
   nand U11530 ( n11153,n11497,n11030,n11498 );
   xor U11531 ( n11497,n10662,n11499 );
   nand U11532 ( n11499,n11500,n11501,n11502,n11503 );
   nor U11533 ( n11503,n11504,n11505,n11506,n11507 );
   nand U11534 ( n11507,n11508,n11509,n11510,n11511 );
   nand U11535 ( n11506,n11512,n11513,n11514,n11515 );
   nand U11536 ( n11505,n11516,n11517,n11518,n11519 );
   nand U11537 ( n11504,n11520,n11521,n11522,n11523 );
   not U11538 ( n11522,n11524 );
   nor U11539 ( n11502,n11525,n11526,n11527,n11528 );
   nand U11540 ( n11526,n11529,n11530 );
   nand U11541 ( n11525,n11531,n11532,n11533,n11534 );
   nor U11542 ( n11501,n11535,n11536,n11537,n11538 );
   nor U11543 ( n11500,n11539,n11540,n11541,n11542 );
   xor U11544 ( n11542,n10457,n10674 );
   xor U11545 ( n11539,n10460,n10679 );
   nand U11546 ( n11545,n11546,p1_datao_reg_0_ );
   nand U11547 ( n11544,p2_ir_reg_0_,n11547 );
   or U11548 ( n11547,n11548,n11549 );
   nand U11549 ( n11543,n11550,n11551 );
   nand U11550 ( n11555,p2_ir_reg_1_,n11556 );
   nand U11551 ( n11556,n11557,n11558 );
   nand U11552 ( n11558,n11549,n11559 );
   nand U11553 ( n11554,n11549,p2_ir_reg_0_,n11560 );
   nand U11554 ( n11553,n11550,n11561 );
   nand U11555 ( n11552,n11546,p1_datao_reg_1_ );
   nand U11556 ( n11565,n11566,n11549 );
   not U11557 ( n11566,n11567 );
   nand U11558 ( n11564,n11550,n11568 );
   nand U11559 ( n11563,n11546,p1_datao_reg_2_ );
   nand U11560 ( n11562,n11548,p2_ir_reg_2_ );
   nand U11561 ( n11572,p2_ir_reg_3_,n11573 );
   nand U11562 ( n11573,n11557,n11574 );
   nand U11563 ( n11574,n11549,n11575 );
   nand U11564 ( n11571,n11549,n11576,n11577 );
   nand U11565 ( n11570,n11550,n11578 );
   nand U11566 ( n11569,n11546,p1_datao_reg_3_ );
   nand U11567 ( n11582,n11583,n11584,n11549 );
   nand U11568 ( n11581,n11585,n11550 );
   nand U11569 ( n11580,n11546,p1_datao_reg_4_ );
   nand U11570 ( n11579,n11548,p2_ir_reg_4_ );
   nand U11571 ( n11589,p2_ir_reg_5_,n11590 );
   nand U11572 ( n11590,n11557,n11591 );
   nand U11573 ( n11591,n11549,n11592 );
   nand U11574 ( n11588,n11549,n11584,n11593 );
   nand U11575 ( n11587,n11594,n11550 );
   nand U11576 ( n11586,n11546,p1_datao_reg_5_ );
   nand U11577 ( n11598,n11599,n11600,n11549 );
   nand U11578 ( n11597,n11550,n11601 );
   nand U11579 ( n11596,n11546,p1_datao_reg_6_ );
   nand U11580 ( n11595,n11548,p2_ir_reg_6_ );
   nand U11581 ( n11605,p2_ir_reg_7_,n11606 );
   nand U11582 ( n11606,n11557,n11607 );
   nand U11583 ( n11607,n11549,n11608 );
   nand U11584 ( n11604,n11549,n11600,n11609 );
   nand U11585 ( n11603,n11610,n11550 );
   nand U11586 ( n11602,n11546,p1_datao_reg_7_ );
   nand U11587 ( n11614,n11615,n11616,n11549 );
   nand U11588 ( n11613,n11617,n11550 );
   nand U11589 ( n11612,n11546,p1_datao_reg_8_ );
   nand U11590 ( n11611,n11548,p2_ir_reg_8_ );
   nand U11591 ( n11621,p2_ir_reg_9_,n11622 );
   nand U11592 ( n11622,n11557,n11623 );
   nand U11593 ( n11623,n11549,n11624 );
   nand U11594 ( n11620,n11549,n11616,n11625 );
   nand U11595 ( n11619,n11626,n11550 );
   nand U11596 ( n11618,n11546,p1_datao_reg_9_ );
   nand U11597 ( n11630,n11631,n11549 );
   not U11598 ( n11631,n11632 );
   nand U11599 ( n11629,n11550,n11633 );
   nand U11600 ( n11628,n11546,p1_datao_reg_10_ );
   nand U11601 ( n11627,n11548,p2_ir_reg_10_ );
   nand U11602 ( n11637,p2_ir_reg_11_,n11638 );
   nand U11603 ( n11638,n11557,n11639 );
   nand U11604 ( n11639,n11549,n11640 );
   nand U11605 ( n11636,n11549,n11641,n11642 );
   nand U11606 ( n11635,n11643,n11550 );
   nand U11607 ( n11634,n11546,p1_datao_reg_11_ );
   nand U11608 ( n11647,n11648,n11549 );
   not U11609 ( n11648,n11649 );
   nand U11610 ( n11646,n11650,n11550 );
   nand U11611 ( n11645,n11546,p1_datao_reg_12_ );
   nand U11612 ( n11644,n11548,p2_ir_reg_12_ );
   nand U11613 ( n11654,p2_ir_reg_13_,n11655 );
   nand U11614 ( n11655,n11557,n11656 );
   nand U11615 ( n11656,n11549,n11657 );
   nand U11616 ( n11653,n11549,n11658,n11659 );
   nand U11617 ( n11652,n11550,n11660 );
   nand U11618 ( n11651,n11546,p1_datao_reg_13_ );
   nand U11619 ( n11664,n11665,n11549 );
   not U11620 ( n11665,n11666 );
   nand U11621 ( n11663,n11550,n11667 );
   nand U11622 ( n11662,n11546,p1_datao_reg_14_ );
   nand U11623 ( n11661,n11548,p2_ir_reg_14_ );
   nand U11624 ( n11671,p2_ir_reg_15_,n11672 );
   nand U11625 ( n11672,n11557,n11673 );
   nand U11626 ( n11673,n11549,n11674 );
   nand U11627 ( n11670,n11549,n11675,n11676 );
   nand U11628 ( n11669,n11677,n11550 );
   nand U11629 ( n11668,n11546,p1_datao_reg_15_ );
   nand U11630 ( n11681,n11682,n11549 );
   not U11631 ( n11682,n11683 );
   nand U11632 ( n11680,n11684,n11550 );
   nand U11633 ( n11679,p1_datao_reg_16_,n11546 );
   nand U11634 ( n11678,n11548,p2_ir_reg_16_ );
   nand U11635 ( n11688,p2_ir_reg_17_,n11689 );
   nand U11636 ( n11689,n11557,n11690 );
   nand U11637 ( n11690,n11549,n11691 );
   nand U11638 ( n11687,n11549,n11692,n11693 );
   nand U11639 ( n11686,n11694,n11550 );
   nand U11640 ( n11685,p1_datao_reg_17_,n11546 );
   nand U11641 ( n11698,p2_ir_reg_18_,n11699 );
   nand U11642 ( n11699,n11557,n11700 );
   nand U11643 ( n11700,n11549,n11701 );
   nand U11644 ( n11697,n11549,n11702,n11703 );
   nand U11645 ( n11696,n11704,n11550 );
   nand U11646 ( n11695,p1_datao_reg_18_,n11546 );
   nand U11647 ( n11708,n11709,n11710,n11549 );
   nand U11648 ( n11707,n11711,n11550 );
   nand U11649 ( n11706,p1_datao_reg_19_,n11546 );
   nand U11650 ( n11705,n11548,p2_ir_reg_19_ );
   nand U11651 ( n11715,n11716,n11717,n11549 );
   nand U11652 ( n11714,n11718,n11550 );
   nand U11653 ( n11713,p1_datao_reg_20_,n11546 );
   nand U11654 ( n11712,n11548,p2_ir_reg_20_ );
   nand U11655 ( n11722,p2_ir_reg_21_,n11723 );
   nand U11656 ( n11723,n11557,n11724 );
   nand U11657 ( n11724,n11549,n11725 );
   nand U11658 ( n11721,n11549,n11717,n11726 );
   nand U11659 ( n11720,n11727,n11550 );
   nand U11660 ( n11719,p1_datao_reg_21_,n11546 );
   nand U11661 ( n11731,n11732,n11549 );
   not U11662 ( n11732,n11733 );
   nand U11663 ( n11730,n11734,n11550 );
   nand U11664 ( n11729,p1_datao_reg_22_,n11546 );
   nand U11665 ( n11728,n11548,p2_ir_reg_22_ );
   nand U11666 ( n11738,p2_ir_reg_23_,n11739 );
   nand U11667 ( n11739,n11557,n11740 );
   nand U11668 ( n11740,n11549,n11741 );
   nand U11669 ( n11737,n11549,n11742,n11743 );
   nand U11670 ( n11736,n11744,n11550 );
   nand U11671 ( n11735,p1_datao_reg_23_,n11546 );
   nand U11672 ( n11748,n11749,n11549 );
   not U11673 ( n11749,n11750 );
   nand U11674 ( n11747,n11751,n11550 );
   nand U11675 ( n11746,p1_datao_reg_24_,n11546 );
   nand U11676 ( n11745,n11548,p2_ir_reg_24_ );
   nand U11677 ( n11755,p2_ir_reg_25_,n11756 );
   nand U11678 ( n11756,n11557,n11757 );
   nand U11679 ( n11757,n11549,n11758 );
   nand U11680 ( n11754,n11549,n11759,n11760 );
   nand U11681 ( n11753,n11761,n11550 );
   nand U11682 ( n11752,p1_datao_reg_25_,n11546 );
   nand U11683 ( n11765,n11766,n11549 );
   not U11684 ( n11766,n11767 );
   nand U11685 ( n11764,n11768,n11550 );
   nand U11686 ( n11763,p1_datao_reg_26_,n11546 );
   nand U11687 ( n11762,n11548,p2_ir_reg_26_ );
   nand U11688 ( n11772,p2_ir_reg_27_,n11773 );
   nand U11689 ( n11773,n11557,n11774 );
   nand U11690 ( n11774,n11549,n11775 );
   nand U11691 ( n11771,n11549,n11776,n11777 );
   nand U11692 ( n11770,n11778,n11550 );
   nand U11693 ( n11769,p1_datao_reg_27_,n11546 );
   nand U11694 ( n11782,p2_ir_reg_28_,n11783 );
   nand U11695 ( n11783,n11557,n11784 );
   nand U11696 ( n11784,n11549,n11785 );
   nand U11697 ( n11781,n11549,n11786,n11787 );
   nand U11698 ( n11780,n11788,n11550 );
   nand U11699 ( n11779,p1_datao_reg_28_,n11546 );
   nand U11700 ( n11792,n11793,n11794,n11549 );
   nand U11701 ( n11791,n11550,n11795 );
   nand U11702 ( n11790,n11546,p1_datao_reg_29_ );
   nand U11703 ( n11789,n11548,p2_ir_reg_29_ );
   nand U11704 ( n11799,p2_ir_reg_30_,n11800 );
   nand U11705 ( n11800,n11557,n11801 );
   nand U11706 ( n11801,n11802,n11549 );
   nand U11707 ( n11798,n11549,n11794,n11803 );
   not U11708 ( n11794,n11802 );
   nand U11709 ( n11797,n11804,n11550 );
   nand U11710 ( n11796,n11546,p1_datao_reg_30_ );
   nand U11711 ( n11807,n11546,p1_datao_reg_31_ );
   nand U11712 ( n11806,n11549,n11803,n11802 );
   nor U11713 ( n11802,n11809,p2_ir_reg_29_ );
   not U11714 ( n11548,n11557 );
   nand U11715 ( n11557,p2_state_reg,n11810 );
   nand U11716 ( n11805,n11550,n11811 );
   nor U11717 ( n11829,n11830,n11831 );
   and U11718 ( n11828,n11016,n11832 );
   nor U11719 ( n11827,n11833,n11834 );
   nand U11720 ( n11825,n11835,n11017 );
   nand U11721 ( n11824,p2_reg2_reg_0_,n11836 );
   nand U11722 ( n11823,n11837,n11018 );
   nand U11723 ( n11018,n11838,n11839 );
   nand U11724 ( n11839,n11016,n11008 );
   or U11725 ( n11838,n11521,n10812 );
   nand U11726 ( n11521,n11840,n11841 );
   nand U11727 ( n11840,n11373,n11006 );
   nor U11728 ( n11849,n10983,n11831 );
   and U11729 ( n11848,n11850,n11007 );
   xor U11730 ( n11007,n11851,n11531 );
   nor U11731 ( n11847,n11006,n11852 );
   and U11732 ( n11846,n11009,n11853 );
   xor U11733 ( n11009,n11841,n11531 );
   nand U11734 ( n11531,n11854,n11855 );
   nand U11735 ( n11855,n11830,n11005 );
   nand U11736 ( n11844,p2_reg2_reg_1_,n11836 );
   nand U11737 ( n11842,n11835,n11379 );
   nor U11738 ( n11863,n10971,n11831 );
   nor U11739 ( n11862,n11864,n11865 );
   nor U11740 ( n11861,n11866,n11834 );
   nand U11741 ( n11859,n11835,n10995 );
   nand U11742 ( n11858,p2_reg2_reg_2_,n11836 );
   nand U11743 ( n11857,n11837,n10996 );
   nand U11744 ( n10996,n11867,n11868,n11869,n11870 );
   nand U11745 ( n11870,n11871,n11872,n11873 );
   nand U11746 ( n11871,n11874,n11875,n11876 );
   nand U11747 ( n11869,n10994,n11877 );
   not U11748 ( n10994,n11864 );
   nand U11749 ( n11864,n11878,n11872 );
   nand U11750 ( n11872,n11879,n11880 );
   not U11751 ( n11879,n11532 );
   nand U11752 ( n11878,n11881,n11875 );
   not U11753 ( n11881,n11882 );
   nand U11754 ( n11868,n11883,n11884,n10733 );
   or U11755 ( n11884,n11532,n11885 );
   nand U11756 ( n11532,n11886,n11887 );
   nand U11757 ( n11883,n11874,n11875,n11885 );
   nor U11758 ( n11885,n11888,n11889 );
   nand U11759 ( n11867,n10781,n10547 );
   nor U11760 ( n11897,n10958,n11831 );
   nor U11761 ( n11896,n10983,n11852 );
   and U11762 ( n11895,n10985,n11853 );
   xor U11763 ( n10985,n11541,n11898 );
   nand U11764 ( n11898,n11899,n11900 );
   nand U11765 ( n11900,n11888,n11886 );
   and U11766 ( n11894,n10986,n11901 );
   nand U11767 ( n10986,n11902,n11903 );
   nand U11768 ( n11902,n11904,n11874,n11541 );
   nand U11769 ( n11904,n11880,n11875 );
   nor U11770 ( n11892,n11905,n11906 );
   nor U11771 ( n11906,n11836,n10977 );
   nand U11772 ( n10977,n11873,n11907 );
   nand U11773 ( n11907,n11903,n11908 );
   nand U11774 ( n11908,n11541,n11132 );
   or U11775 ( n11903,n11541,n11132 );
   xor U11776 ( n11541,n11133,n10541 );
   nor U11777 ( n11905,n11837,n11909 );
   nand U11778 ( n11890,n11835,n11133 );
   nor U11779 ( n11918,n11919,n11831 );
   and U11780 ( n11917,n11850,n10972 );
   nand U11781 ( n10972,n11920,n11921 );
   nand U11782 ( n11921,n11922,n11533 );
   nand U11783 ( n11920,n11923,n11924 );
   nand U11784 ( n11923,n11925,n11926 );
   nor U11785 ( n11916,n10971,n11852 );
   nor U11786 ( n11915,n10973,n11927 );
   xor U11787 ( n10973,n11533,n11928 );
   nand U11788 ( n11533,n11929,n11930 );
   nand U11789 ( n11913,p2_reg2_reg_4_,n11836 );
   nand U11790 ( n11911,n11835,n11386 );
   nor U11791 ( n11939,n10935,n11831 );
   and U11792 ( n11938,n11850,n10961 );
   nand U11793 ( n10961,n11940,n11941 );
   nand U11794 ( n11941,n11942,n11534 );
   nand U11795 ( n11940,n11943,n11944 );
   nand U11796 ( n11943,n11945,n11946 );
   nor U11797 ( n11937,n10958,n11852 );
   and U11798 ( n11936,n11853,n10960,n10959 );
   nand U11799 ( n10959,n11947,n11930,n11948 );
   not U11800 ( n11948,n11534 );
   nand U11801 ( n10960,n11949,n11534 );
   nand U11802 ( n11534,n11950,n11951 );
   nand U11803 ( n11949,n11947,n11930 );
   nand U11804 ( n11947,n11952,n11929 );
   not U11805 ( n11952,n11928 );
   nand U11806 ( n11934,p2_reg2_reg_5_,n11836 );
   nand U11807 ( n11932,n11835,n11404 );
   nor U11808 ( n11960,n11961,n11831 );
   and U11809 ( n11959,n10946,n11832 );
   and U11810 ( n11958,n11962,n11856 );
   nand U11811 ( n11956,n11835,n10947 );
   nand U11812 ( n11955,p2_reg2_reg_6_,n11836 );
   nand U11813 ( n11954,n11837,n10948 );
   nand U11814 ( n10948,n11963,n11964,n11965 );
   nand U11815 ( n11965,n10781,n10535 );
   nand U11816 ( n11964,n11966,n10733 );
   xor U11817 ( n11966,n11508,n11967 );
   nand U11818 ( n11963,n11968,n10946 );
   nand U11819 ( n10946,n11969,n11970 );
   nand U11820 ( n11970,n11971,n11143,n11946,n11972 );
   nand U11821 ( n11971,n11944,n11945 );
   nand U11822 ( n11969,n11973,n11945,n11974 );
   not U11823 ( n11974,n11508 );
   nand U11824 ( n11508,n11975,n11976 );
   nand U11825 ( n11973,n11942,n11946 );
   not U11826 ( n11942,n11944 );
   nand U11827 ( n11944,n11926,n11977 );
   nand U11828 ( n11977,n11924,n11925 );
   nand U11829 ( n11968,n11978,n11979,n11980 );
   nor U11830 ( n11988,n10936,n11989 );
   and U11831 ( n11987,n11990,n11856 );
   nor U11832 ( n11986,n11836,n10929 );
   nand U11833 ( n10929,n10937,n11873 );
   nor U11834 ( n11985,n11837,n11991 );
   nor U11835 ( n11983,n11992,n11993 );
   and U11836 ( n11993,n11901,n10937 );
   and U11837 ( n10937,n11994,n11995 );
   nand U11838 ( n11995,n11538,n11996 );
   nand U11839 ( n11994,n11997,n11144 );
   and U11840 ( n11992,n11853,n10938,n10939 );
   nand U11841 ( n10939,n11998,n11975,n11999 );
   not U11842 ( n11999,n11538 );
   nand U11843 ( n11998,n12000,n11976 );
   nand U11844 ( n10938,n12001,n11976,n11538 );
   xor U11845 ( n11538,n11413,n10529 );
   nand U11846 ( n12001,n11975,n11967 );
   nand U11847 ( n11982,n12002,n10532 );
   nand U11848 ( n11981,n12003,n10526 );
   nor U11849 ( n12007,n12008,n12009,n12010 );
   nor U11850 ( n12010,n10901,n11831 );
   nor U11851 ( n12009,n12011,n11865 );
   nor U11852 ( n12008,n12012,n11834 );
   nand U11853 ( n12006,n11835,n10924 );
   nand U11854 ( n12005,p2_reg2_reg_8_,n11836 );
   nand U11855 ( n10925,n12013,n12014,n12015,n12016 );
   nor U11856 ( n12016,n12017,n12018,n12019,n12020 );
   nor U11857 ( n12020,n12021,n11979 );
   and U11858 ( n12021,n12022,n12023 );
   and U11859 ( n12019,n12024,n12025 );
   nor U11860 ( n12018,n12011,n11980 );
   not U11861 ( n12011,n10923 );
   nand U11862 ( n10923,n12022,n12026 );
   nand U11863 ( n12026,n12027,n12028,n11537 );
   nand U11864 ( n12027,n11996,n11144 );
   not U11865 ( n11996,n12029 );
   nor U11866 ( n12017,n11961,n10727 );
   nand U11867 ( n12015,n11873,n12030 );
   nand U11868 ( n12030,n12023,n12022 );
   or U11869 ( n12022,n11997,n12031,n11537 );
   not U11870 ( n11997,n12032 );
   nand U11871 ( n12023,n11537,n12033 );
   nand U11872 ( n12033,n12032,n11144 );
   nand U11873 ( n12032,n12029,n12028 );
   nand U11874 ( n12014,n12024,n12034 );
   nand U11875 ( n12013,n11051,n12024 );
   xor U11876 ( n12024,n12035,n11537 );
   xor U11877 ( n11537,n12036,n10914 );
   not U11878 ( n11051,n12037 );
   nor U11879 ( n12045,n10887,n11831 );
   and U11880 ( n12044,n11850,n10915 );
   xor U11881 ( n10915,n11509,n12046 );
   nor U11882 ( n12043,n10914,n11852 );
   nor U11883 ( n12042,n10916,n11927 );
   xor U11884 ( n10916,n12047,n11509 );
   nand U11885 ( n11509,n12048,n12049 );
   nand U11886 ( n12040,p2_reg2_reg_9_,n11836 );
   nand U11887 ( n12039,n11856,n12050 );
   nand U11888 ( n12038,n11835,n11340 );
   nor U11889 ( n12058,n10872,n11831 );
   and U11890 ( n12057,n11850,n10904 );
   nand U11891 ( n10904,n12059,n12060 );
   nand U11892 ( n12060,n12061,n11510 );
   nand U11893 ( n12059,n12062,n12063 );
   nand U11894 ( n12062,n12064,n12065 );
   nor U11895 ( n12056,n10901,n11852 );
   and U11896 ( n12055,n11853,n10903,n10902 );
   nand U11897 ( n10902,n11510,n12049,n12066 );
   nand U11898 ( n10903,n12067,n12048,n12068 );
   not U11899 ( n12068,n11510 );
   nand U11900 ( n11510,n12069,n12070 );
   nand U11901 ( n12067,n12071,n12049 );
   not U11902 ( n12071,n12047 );
   nand U11903 ( n12053,p2_reg2_reg_10_,n11836 );
   nand U11904 ( n12052,n11856,n12072 );
   nand U11905 ( n12051,n11835,n11419 );
   nor U11906 ( n12080,n10888,n11831 );
   nor U11907 ( n12079,n10887,n11852 );
   nor U11908 ( n12078,n10890,n11927 );
   xor U11909 ( n10890,n11524,n12081 );
   and U11910 ( n12077,n10891,n11901 );
   nor U11911 ( n12075,n12082,n12083 );
   nor U11912 ( n12083,n11836,n10881 );
   nand U11913 ( n10881,n11873,n10891 );
   nand U11914 ( n10891,n12084,n12085 );
   nand U11915 ( n12085,n12086,n11117,n11123 );
   nand U11916 ( n12086,n12064,n12063 );
   not U11917 ( n12063,n12061 );
   nand U11918 ( n12084,n12087,n12064,n11524 );
   nor U11919 ( n11524,n12088,n12089 );
   nand U11920 ( n12087,n12061,n12065 );
   nor U11921 ( n12061,n11137,n12090 );
   and U11922 ( n12090,n12091,n12046 );
   nor U11923 ( n12082,n11837,n12092 );
   nand U11924 ( n12074,n11856,n12093 );
   nand U11925 ( n12073,n11835,n11430 );
   nor U11926 ( n12101,n10874,n11989 );
   nor U11927 ( n12100,n12102,n11834 );
   nor U11928 ( n12099,n11836,n10866 );
   nand U11929 ( n10866,n11873,n10876 );
   nor U11930 ( n12098,n11837,n12103 );
   nor U11931 ( n12096,n12104,n12105 );
   nor U11932 ( n12105,n10873,n11831 );
   nor U11933 ( n12104,n10872,n11852 );
   nand U11934 ( n12095,n10876,n11901 );
   nand U11935 ( n11901,n11865,n12106 );
   nand U11936 ( n12106,n11837,n11877 );
   nand U11937 ( n10876,n12107,n12108 );
   nand U11938 ( n12108,n12109,n12110 );
   nand U11939 ( n12110,n12111,n12112 );
   nand U11940 ( n12107,n12111,n12112,n11511 );
   xor U11941 ( n10875,n12109,n12113 );
   not U11942 ( n12109,n11511 );
   nand U11943 ( n11511,n12114,n12115 );
   nor U11944 ( n12119,n12120,n12121,n12122 );
   nor U11945 ( n12122,n12123,n11831 );
   and U11946 ( n12121,n10860,n11832 );
   and U11947 ( n12120,n12124,n11856 );
   nand U11948 ( n12118,n11835,n10861 );
   nand U11949 ( n12117,p2_reg2_reg_13_,n11836 );
   nand U11950 ( n10862,n12125,n12126,n12127 );
   nand U11951 ( n12127,n10781,n10514 );
   nand U11952 ( n12126,n12128,n12129,n10733 );
   nand U11953 ( n12129,n12130,n12115,n11512 );
   nand U11954 ( n12130,n12113,n12114 );
   not U11955 ( n12113,n12131 );
   nand U11956 ( n12128,n12132,n12114,n12133 );
   nand U11957 ( n12132,n12131,n12115 );
   nor U11958 ( n12131,n12088,n12134 );
   nand U11959 ( n12125,n10860,n11008 );
   xor U11960 ( n10860,n12133,n12135 );
   not U11961 ( n12133,n11512 );
   nand U11962 ( n11512,n12136,n12137 );
   nor U11963 ( n12141,n12142,n12143,n12144 );
   nor U11964 ( n12144,n10835,n11831 );
   nor U11965 ( n12143,n10851,n11865 );
   and U11966 ( n12142,n12145,n11856 );
   nand U11967 ( n12140,n11835,n10852 );
   nand U11968 ( n12139,p2_reg2_reg_14_,n11836 );
   nand U11969 ( n10853,n12146,n12147 );
   nor U11970 ( n12147,n12148,n12149,n12150,n12151 );
   nor U11971 ( n12151,n11049,n12152 );
   nor U11972 ( n12150,n11978,n10851 );
   nor U11973 ( n12149,n11979,n10851 );
   nor U11974 ( n12148,n12153,n12152 );
   nor U11975 ( n12146,n12154,n12155,n12156,n12157 );
   nor U11976 ( n12157,n10873,n10727 );
   nor U11977 ( n12156,n12037,n12152 );
   nor U11978 ( n12155,n12158,n12152 );
   not U11979 ( n12152,n12159 );
   xor U11980 ( n12159,n11540,n12160 );
   nor U11981 ( n12154,n11980,n10851 );
   nand U11982 ( n10851,n12161,n12162 );
   nand U11983 ( n12162,n11540,n12163 );
   xor U11984 ( n11540,n12164,n12123 );
   nand U11985 ( n12161,n11111,n12165,n12166 );
   nor U11986 ( n12173,n10839,n11836 );
   and U11987 ( n10839,n12174,n12175 );
   nor U11988 ( n12175,n12176,n12177,n12178,n12179 );
   nor U11989 ( n12179,n11049,n12180 );
   nor U11990 ( n12178,n11978,n12181 );
   nor U11991 ( n12177,n11979,n12181 );
   nor U11992 ( n12176,n12153,n12180 );
   nor U11993 ( n12174,n12182,n12183,n12184,n12185 );
   nor U11994 ( n12185,n12123,n10727 );
   nor U11995 ( n12184,n12037,n12180 );
   nor U11996 ( n12183,n12158,n12180 );
   xor U11997 ( n12180,n11536,n12186 );
   nor U11998 ( n12182,n11980,n12181 );
   nor U11999 ( n12172,n11837,n12187 );
   nor U12000 ( n12171,n12188,n11989 );
   nand U12001 ( n12169,n11856,n12189 );
   nand U12002 ( n12168,n11832,n10843 );
   not U12003 ( n10843,n12181 );
   nand U12004 ( n12181,n12190,n12191 );
   nand U12005 ( n12191,n11536,n12192 );
   xor U12006 ( n11536,n12188,n10835 );
   nand U12007 ( n12190,n12193,n11110,n12194 );
   nand U12008 ( n12167,n12003,n10502 );
   nor U12009 ( n12202,n10834,n11989 );
   and U12010 ( n12201,n12203,n11856 );
   nor U12011 ( n12200,n11836,n10829 );
   nand U12012 ( n10829,n12204,n10733 );
   xor U12013 ( n12204,n12205,n12206 );
   nor U12014 ( n12199,n11837,n12207 );
   nand U12015 ( n12197,n12003,n10499 );
   nand U12016 ( n12196,n12002,n10505 );
   nand U12017 ( n12195,n11850,n10836 );
   nand U12018 ( n10836,n12208,n12209 );
   nand U12019 ( n12209,n12210,n11104,n12193,n11106 );
   nand U12020 ( n12210,n11110,n12194 );
   nand U12021 ( n12208,n12211,n11110,n12206 );
   not U12022 ( n12206,n11513 );
   nand U12023 ( n11513,n12212,n12213 );
   nand U12024 ( n12211,n12192,n12193 );
   not U12025 ( n12192,n12194 );
   nand U12026 ( n12194,n12214,n12165 );
   nand U12027 ( n12214,n12166,n11111 );
   nor U12028 ( n12222,n11146,n11831 );
   and U12029 ( n12221,n11850,n10825 );
   xor U12030 ( n10825,n12223,n11535 );
   nor U12031 ( n12220,n10822,n11852 );
   nor U12032 ( n12219,n11927,n10823,n10824 );
   and U12033 ( n10824,n12224,n12212,n11535 );
   nand U12034 ( n12224,n12225,n12213 );
   nor U12035 ( n10823,n12226,n11535 );
   xor U12036 ( n11535,n10499,n11270 );
   nand U12037 ( n12217,p2_reg2_reg_17_,n11836 );
   nand U12038 ( n12216,n11856,n12227 );
   nand U12039 ( n12215,n11835,n11270 );
   nor U12040 ( n12235,n12236,n11831 );
   and U12041 ( n12234,n11850,n10809 );
   xor U12042 ( n10809,n12237,n12238 );
   nand U12043 ( n11850,n11865,n12239 );
   nor U12044 ( n12233,n10808,n11852 );
   nor U12045 ( n12232,n10811,n11927 );
   xor U12046 ( n10811,n11514,n12240 );
   not U12047 ( n11514,n12238 );
   nor U12048 ( n12238,n12241,n12242 );
   nor U12049 ( n12242,n10496,n11147 );
   nand U12050 ( n12230,p2_reg2_reg_18_,n11836 );
   nand U12051 ( n12229,n11856,n12243 );
   nand U12052 ( n12228,n11835,n11147 );
   nor U12053 ( n12250,n10793,n11836 );
   and U12054 ( n10793,n12251,n12252,n12253,n12254 );
   nor U12055 ( n12254,n12255,n12256,n12257,n12258 );
   nor U12056 ( n12258,n11978,n12259 );
   nor U12057 ( n12257,n12037,n12260 );
   nor U12058 ( n12256,n12153,n12260 );
   nor U12059 ( n12255,n12158,n12260 );
   nor U12060 ( n12253,n12261,n12262 );
   nor U12061 ( n12262,n11146,n10727 );
   nor U12062 ( n12261,n11979,n12259 );
   or U12063 ( n12252,n12260,n11049 );
   xor U12064 ( n12260,n11523,n12263 );
   nand U12065 ( n12251,n10797,n12264 );
   and U12066 ( n12249,n11836,p2_reg2_reg_19_ );
   nor U12067 ( n12248,n12265,n11989 );
   nand U12068 ( n12246,n11856,n12266 );
   nand U12069 ( n12245,n11832,n10797 );
   not U12070 ( n10797,n12259 );
   xor U12071 ( n12259,n11523,n12267 );
   nand U12072 ( n11523,n12268,n12269 );
   nand U12073 ( n12244,n12003,n10490 );
   nor U12074 ( n12276,n10785,n11836 );
   and U12075 ( n10785,n12277,n12278,n12279,n12280 );
   nor U12076 ( n12280,n12281,n12282,n12283,n12284 );
   nor U12077 ( n12284,n12236,n10727 );
   nor U12078 ( n12283,n11980,n12285 );
   nor U12079 ( n12282,n12153,n12286,n12287 );
   nor U12080 ( n12281,n12158,n12286,n12287 );
   nor U12081 ( n12279,n12288,n12289 );
   nor U12082 ( n12289,n12037,n12286,n12287 );
   not U12083 ( n12287,n12290 );
   not U12084 ( n12286,n12291 );
   nor U12085 ( n12288,n11979,n12285 );
   nand U12086 ( n12278,n12290,n12291,n12025 );
   not U12087 ( n12025,n11049 );
   nand U12088 ( n12291,n11515,n12269,n12292 );
   nand U12089 ( n12292,n12268,n12263 );
   nand U12090 ( n12290,n12293,n12294,n12295 );
   nand U12091 ( n12293,n12296,n12269 );
   nand U12092 ( n12277,n10789,n11873 );
   and U12093 ( n12275,n11836,p2_reg2_reg_20_ );
   nor U12094 ( n12274,n12297,n11989 );
   nand U12095 ( n12272,n11856,n12298 );
   nand U12096 ( n12271,n11832,n10789 );
   not U12097 ( n10789,n12285 );
   xor U12098 ( n12285,n11515,n12299 );
   nand U12099 ( n11515,n12294,n12300 );
   nand U12100 ( n12270,n12003,n10487 );
   nor U12101 ( n12308,n10780,n11989 );
   and U12102 ( n12307,n12309,n11856 );
   and U12103 ( n12306,n10779,n11837 );
   nand U12104 ( n10779,n12310,n12311 );
   nand U12105 ( n12311,n12312,n12313,n10733 );
   nand U12106 ( n12313,n12314,n12315,n11516 );
   nand U12107 ( n12315,n12295,n12263 );
   not U12108 ( n12263,n12296 );
   nand U12109 ( n12312,n12316,n12317,n12318 );
   not U12110 ( n12318,n11516 );
   nand U12111 ( n12317,n12314,n12319 );
   nand U12112 ( n12316,n12296,n12314 );
   nor U12113 ( n12296,n12241,n12320 );
   nand U12114 ( n12310,n10782,n11008 );
   and U12115 ( n12305,n11836,p2_reg2_reg_21_ );
   nand U12116 ( n12303,n12003,n10484 );
   nand U12117 ( n12302,n12002,n10490 );
   nand U12118 ( n12301,n11832,n10782 );
   and U12119 ( n10782,n12321,n12322 );
   or U12120 ( n12322,n11516,n12323 );
   nand U12121 ( n11516,n12324,n12325 );
   nand U12122 ( n12321,n11087,n12326,n12323 );
   nor U12123 ( n12330,n12331,n12332,n12333 );
   nor U12124 ( n12333,n10745,n11831 );
   and U12125 ( n12332,n10769,n11832 );
   nand U12126 ( n10769,n12334,n12335 );
   or U12127 ( n12335,n12336,n12337 );
   nand U12128 ( n12334,n12337,n11529 );
   and U12129 ( n12331,n12338,n11856 );
   nand U12130 ( n12329,n11835,n10770 );
   nand U12131 ( n12328,p2_reg2_reg_22_,n11836 );
   nand U12132 ( n10771,n12339,n12340,n12341,n12342 );
   nor U12133 ( n12342,n12343,n12344,n12345,n12346 );
   nor U12134 ( n12346,n11979,n12347 );
   nor U12135 ( n12345,n12348,n12037 );
   nor U12136 ( n12344,n12348,n11049 );
   nor U12137 ( n12343,n12349,n10727 );
   nand U12138 ( n12341,n12350,n11873 );
   nand U12139 ( n12340,n12351,n12034 );
   nand U12140 ( n12034,n12153,n12158 );
   not U12141 ( n12351,n12348 );
   xor U12142 ( n12348,n11529,n12352 );
   nand U12143 ( n12339,n12350,n12264 );
   not U12144 ( n12350,n12347 );
   nand U12145 ( n12347,n12353,n12354 );
   nand U12146 ( n12354,n12336,n12355 );
   nor U12147 ( n12336,n11081,n12356 );
   or U12148 ( n12353,n12355,n11529 );
   xor U12149 ( n11529,n10484,n12357 );
   nor U12150 ( n12365,n10760,n11989 );
   and U12151 ( n12364,n12366,n11856 );
   nor U12152 ( n12363,n11836,n10753 );
   nand U12153 ( n10753,n11008,n10761 );
   and U12154 ( n12362,n11836,p2_reg2_reg_23_ );
   nor U12155 ( n12360,n12367,n12368 );
   nor U12156 ( n12368,n10759,n11852 );
   and U12157 ( n12367,n10762,n11853 );
   xor U12158 ( n10762,n11530,n12369 );
   nand U12159 ( n12359,n11832,n10761 );
   nand U12160 ( n10761,n12370,n12371,n12372 );
   and U12161 ( n12372,n12373,n12374 );
   nand U12162 ( n12374,n11081,n12375 );
   nand U12163 ( n12373,n12356,n12376 );
   nand U12164 ( n12371,n12376,n12355 );
   nor U12165 ( n12376,n11530,n11081 );
   not U12166 ( n11081,n12377 );
   xor U12167 ( n11530,n10481,n10760 );
   nand U12168 ( n12370,n12337,n12375 );
   and U12169 ( n12375,n11080,n11149 );
   not U12170 ( n12337,n12355 );
   nand U12171 ( n12355,n12378,n12326 );
   nand U12172 ( n12378,n12323,n11087 );
   nand U12173 ( n12358,n12003,n10478 );
   nor U12174 ( n12382,n12383,n12384,n12385,n12386 );
   and U12175 ( n12386,n11836,p2_reg2_reg_24_ );
   nor U12176 ( n12385,n10747,n11989 );
   and U12177 ( n12384,n12387,n11856 );
   nor U12178 ( n12383,n10746,n11831 );
   nor U12179 ( n12381,n12388,n12389 );
   nor U12180 ( n12389,n10749,n11865 );
   nor U12181 ( n12388,n10749,n12239 );
   xor U12182 ( n10749,n12390,n11517 );
   nand U12183 ( n12380,n11853,n10748 );
   xor U12184 ( n10748,n12391,n11517 );
   nand U12185 ( n11517,n12392,n12393 );
   nand U12186 ( n12379,n12002,n10481 );
   nor U12187 ( n12397,n12398,n12399,n12400,n12401 );
   and U12188 ( n12401,n11836,p2_reg2_reg_25_ );
   nor U12189 ( n12400,n10731,n11989 );
   and U12190 ( n12399,n12402,n11856 );
   nor U12191 ( n12398,n10728,n11831 );
   nor U12192 ( n12396,n12403,n12404 );
   nor U12193 ( n12404,n10734,n11865 );
   nor U12194 ( n12403,n10734,n12239 );
   nand U12195 ( n12239,n11837,n11008 );
   xor U12196 ( n10734,n11518,n12405 );
   nand U12197 ( n12395,n11853,n10732 );
   xor U12198 ( n10732,n11518,n12406 );
   nand U12199 ( n11518,n12407,n12408 );
   not U12200 ( n11853,n11927 );
   nand U12201 ( n11927,n11837,n10733 );
   nand U12202 ( n12394,n12002,n10478 );
   not U12203 ( n12002,n11852 );
   nand U12204 ( n11852,n11837,n10781 );
   nor U12205 ( n12412,n12413,n12414,n12415 );
   nor U12206 ( n12415,n12416,n11831 );
   nor U12207 ( n12414,n11865,n10713,n10712 );
   nor U12208 ( n10712,n12417,n12418 );
   nor U12209 ( n10713,n11519,n12419 );
   and U12210 ( n12413,n12420,n11856 );
   nand U12211 ( n12411,n11835,n10715 );
   nand U12212 ( n12410,p2_reg2_reg_26_,n11836 );
   nand U12213 ( n10716,n12421,n12422,n12423,n12424 );
   nand U12214 ( n12424,n12425,n12426,n11877 );
   nand U12215 ( n12423,n10733,n12427,n12428 );
   nand U12216 ( n12428,n12429,n12430,n12431 );
   nand U12217 ( n12427,n12432,n11519 );
   nand U12218 ( n12432,n12429,n12407 );
   nand U12219 ( n12429,n12408,n12406 );
   nand U12220 ( n12406,n12392,n12433 );
   nand U12221 ( n12433,n12393,n12391 );
   nand U12222 ( n12422,n12425,n12426,n11873 );
   not U12223 ( n11873,n11978 );
   nand U12224 ( n12426,n12434,n12418 );
   not U12225 ( n12434,n11519 );
   nand U12226 ( n11519,n12430,n12435 );
   nand U12227 ( n12425,n12436,n12419 );
   not U12228 ( n12436,n12417 );
   nand U12229 ( n12417,n12437,n11071 );
   nand U12230 ( n12421,n10781,n10475 );
   nor U12231 ( n12444,n10700,n11836 );
   and U12232 ( n10700,n12445,n12446 );
   nor U12233 ( n12446,n12447,n12448,n12449,n12450 );
   nor U12234 ( n12450,n11978,n12451,n12452 );
   nor U12235 ( n12452,n12453,n11520 );
   and U12236 ( n12453,n12454,n11071 );
   nor U12237 ( n12451,n12455,n12456 );
   nor U12238 ( n12449,n12037,n12457 );
   nor U12239 ( n12448,n12458,n11979 );
   nor U12240 ( n12447,n12458,n11980 );
   and U12241 ( n12458,n12459,n12460 );
   nand U12242 ( n12460,n12456,n11520 );
   and U12243 ( n12456,n12437,n12461 );
   nor U12244 ( n12445,n12462,n12463,n12464,n12465 );
   nor U12245 ( n12465,n10728,n10727 );
   nor U12246 ( n12464,n12158,n12457 );
   nor U12247 ( n12463,n11049,n12457 );
   nor U12248 ( n12462,n12153,n12457 );
   xor U12249 ( n12457,n11520,n12466 );
   nand U12250 ( n12466,n12430,n12467,n12468 );
   and U12251 ( n12443,n11836,p2_reg2_reg_27_ );
   nor U12252 ( n12442,n12469,n11989 );
   nand U12253 ( n12440,n11856,n12470 );
   nand U12254 ( n12439,n11832,n10704 );
   nand U12255 ( n10704,n12459,n12471 );
   nand U12256 ( n12471,n12461,n12437,n11520 );
   nand U12257 ( n12459,n12454,n11071,n12455 );
   not U12258 ( n12455,n11520 );
   nand U12259 ( n11520,n12472,n12473 );
   nand U12260 ( n12454,n12437,n12418 );
   nand U12261 ( n12438,n12003,n10466 );
   nor U12262 ( n12480,n10691,n11836 );
   and U12263 ( n10691,n12481,n12482,n12483,n12484 );
   nor U12264 ( n12484,n12485,n12486,n12487,n12488 );
   nor U12265 ( n12488,n12489,n11980 );
   nor U12266 ( n12487,n12489,n11978 );
   nor U12267 ( n12486,n12490,n12153 );
   nor U12268 ( n12485,n12490,n11049 );
   nor U12269 ( n12483,n12491,n12492 );
   nor U12270 ( n12492,n12416,n10727 );
   nor U12271 ( n12491,n11979,n12489 );
   xor U12272 ( n12489,n12493,n12494 );
   or U12273 ( n12482,n12037,n12490 );
   or U12274 ( n12481,n12158,n12490 );
   xor U12275 ( n12490,n12494,n12495 );
   and U12276 ( n12479,n11836,p2_reg2_reg_28_ );
   nor U12277 ( n12478,n12496,n11989 );
   nand U12278 ( n12476,n11856,n12497 );
   nand U12279 ( n12475,n11832,n10695 );
   xor U12280 ( n10695,n12494,n12498 );
   nand U12281 ( n12474,n12003,n10463 );
   not U12282 ( n12003,n11831 );
   nand U12283 ( n10729,n12499,n12500 );
   nor U12284 ( n12504,n12505,n12506 );
   nor U12285 ( n12506,n11064,n11989 );
   not U12286 ( n11989,n11835 );
   and U12287 ( n12505,n10687,n11832 );
   not U12288 ( n11832,n11865 );
   nand U12289 ( n11865,n12507,n12508,n11837 );
   nand U12290 ( n10687,n12509,n12510,n12511 );
   nand U12291 ( n12510,n11527,n11068,n12498 );
   nand U12292 ( n12509,n12512,n12513 );
   not U12293 ( n12512,n12498 );
   nand U12294 ( n12498,n11069,n12514 );
   or U12295 ( n12514,n12461,n11075 );
   not U12296 ( n11075,n12515 );
   nand U12297 ( n12461,n12419,n11071 );
   nand U12298 ( n12502,p2_reg2_reg_29_,n11836 );
   nand U12299 ( n10685,n12516,n12517,n12518,n12519 );
   nand U12300 ( n12519,n12520,n10460,n12499 );
   nand U12301 ( n10460,n12521,n12522,n12523,n12524 );
   nand U12302 ( n12523,p2_reg2_reg_30_,n12525 );
   nand U12303 ( n12522,p2_reg1_reg_30_,n12526 );
   nand U12304 ( n12521,p2_reg0_reg_30_,n12527 );
   or U12305 ( n12518,n12528,n10812 );
   xor U12306 ( n12528,n11527,n12529 );
   nand U12307 ( n12529,n12530,n12531 );
   nand U12308 ( n12531,n12532,n12533 );
   nand U12309 ( n12533,n10697,n12495 );
   or U12310 ( n12530,n12495,n10697 );
   nand U12311 ( n12495,n12534,n12535,n12536,n12473 );
   nand U12312 ( n12473,n10705,n10469 );
   nand U12313 ( n12536,n12537,n12472 );
   not U12314 ( n12537,n12467 );
   nand U12315 ( n12467,n12431,n12538 );
   nand U12316 ( n12538,n12408,n12393 );
   nand U12317 ( n12393,n11470,n10478 );
   nand U12318 ( n12408,n11475,n10475 );
   nand U12319 ( n12535,n12539,n12472 );
   not U12320 ( n12539,n12430 );
   nand U12321 ( n12430,n10715,n10472 );
   nand U12322 ( n12534,n12540,n12472 );
   nand U12323 ( n12472,n12416,n12469 );
   not U12324 ( n12540,n12468 );
   nand U12325 ( n12468,n12431,n12392,n12541 );
   not U12326 ( n12541,n12391 );
   nand U12327 ( n12391,n12542,n12543 );
   nand U12328 ( n12543,n12544,n10760 );
   or U12329 ( n12544,n12369,n10745 );
   nand U12330 ( n12542,n10745,n12369 );
   nand U12331 ( n12369,n12545,n12546 );
   nand U12332 ( n12546,n12547,n12357 );
   nand U12333 ( n12547,n10484,n12352 );
   or U12334 ( n12545,n12352,n10484 );
   nand U12335 ( n12352,n12548,n12324,n12549 );
   nand U12336 ( n12549,n12325,n12550 );
   nand U12337 ( n12550,n12314,n12551 );
   nand U12338 ( n12551,n12241,n12295 );
   nor U12339 ( n12241,n10807,n11146 );
   and U12340 ( n12314,n12294,n12552 );
   nand U12341 ( n12552,n12553,n12300 );
   not U12342 ( n12553,n12269 );
   nand U12343 ( n12269,n10798,n10493 );
   nand U12344 ( n12294,n10790,n10490 );
   nand U12345 ( n12324,n11448,n10487 );
   nand U12346 ( n12548,n12295,n12325,n12320 );
   and U12347 ( n12320,n12554,n12240 );
   nand U12348 ( n12240,n12555,n12556 );
   nand U12349 ( n12556,n12557,n10499 );
   or U12350 ( n12557,n12226,n11270 );
   nand U12351 ( n12555,n11270,n12226 );
   nand U12352 ( n12226,n12213,n12558 );
   nand U12353 ( n12558,n12205,n12212 );
   nand U12354 ( n12212,n10822,n10834 );
   not U12355 ( n12205,n12225 );
   nand U12356 ( n12225,n12559,n12560 );
   nand U12357 ( n12560,n12561,n12188 );
   or U12358 ( n12561,n12186,n10835 );
   nand U12359 ( n12559,n10835,n12186 );
   nand U12360 ( n12186,n12562,n12563 );
   nand U12361 ( n12563,n12164,n12564 );
   nand U12362 ( n12564,n10508,n12160 );
   or U12363 ( n12562,n12160,n10508 );
   nand U12364 ( n12160,n12565,n12136,n12566 );
   nand U12365 ( n12566,n12137,n12567 );
   nand U12366 ( n12567,n12568,n12115 );
   nand U12367 ( n12115,n11425,n10514 );
   nand U12368 ( n12568,n12088,n12114 );
   nor U12369 ( n12088,n10889,n10872 );
   nand U12370 ( n12136,n10861,n10511 );
   nand U12371 ( n12565,n12137,n12114,n12134 );
   nor U12372 ( n12134,n12089,n12081 );
   and U12373 ( n12081,n12070,n12569 );
   nand U12374 ( n12569,n12570,n12069 );
   nand U12375 ( n12069,n10887,n10900 );
   nand U12376 ( n12570,n12049,n12066 );
   nand U12377 ( n12066,n12048,n12047 );
   nand U12378 ( n12047,n12571,n12572 );
   nand U12379 ( n12572,n12573,n12035 );
   nand U12380 ( n12035,n12574,n12575,n12576 );
   or U12381 ( n12576,n11975,n11961 );
   nand U12382 ( n12575,n12577,n11976,n12000 );
   not U12383 ( n12000,n11967 );
   nand U12384 ( n11967,n12578,n11950 );
   nand U12385 ( n11950,n11919,n10957 );
   nand U12386 ( n12578,n12579,n11929,n11951 );
   nand U12387 ( n11951,n11404,n10535 );
   nand U12388 ( n11929,n11386,n10538 );
   nand U12389 ( n12579,n11928,n11930 );
   nand U12390 ( n11930,n10958,n10970 );
   nand U12391 ( n11928,n12580,n12581,n12582 );
   nand U12392 ( n12582,n12583,n10541 );
   nand U12393 ( n12581,n12584,n11886,n11888 );
   nor U12394 ( n11888,n11841,n12585 );
   nor U12395 ( n12585,n10547,n11379 );
   nand U12396 ( n12584,n10971,n10984 );
   nand U12397 ( n12580,n12586,n11133 );
   nand U12398 ( n12586,n11899,n10971 );
   not U12399 ( n11899,n12583 );
   nand U12400 ( n12583,n11887,n12587 );
   nand U12401 ( n12587,n11889,n11886 );
   nand U12402 ( n11886,n10983,n12588 );
   not U12403 ( n11889,n11854 );
   nand U12404 ( n11854,n11379,n10547 );
   nand U12405 ( n11887,n10995,n10544 );
   nand U12406 ( n11976,n10935,n12589 );
   nand U12407 ( n12577,n11961,n10936 );
   nand U12408 ( n12574,n11413,n12590 );
   nand U12409 ( n12590,n11961,n11975 );
   nand U12410 ( n11975,n10947,n10532 );
   nand U12411 ( n12573,n10914,n12036 );
   nand U12412 ( n12571,n10924,n10526 );
   nand U12413 ( n12048,n10901,n10913 );
   nand U12414 ( n12049,n11340,n10523 );
   nand U12415 ( n12070,n11419,n10520 );
   nor U12416 ( n12089,n10517,n11430 );
   nand U12417 ( n12114,n10888,n10874 );
   nand U12418 ( n12137,n10873,n11116 );
   nand U12419 ( n12213,n11265,n10502 );
   nand U12420 ( n12554,n11146,n10807 );
   nand U12421 ( n12325,n12349,n10780 );
   not U12422 ( n12295,n12319 );
   nand U12423 ( n12319,n12268,n12300 );
   nand U12424 ( n12300,n12591,n12297 );
   nand U12425 ( n12268,n12236,n12265 );
   nand U12426 ( n12392,n10726,n10747 );
   and U12427 ( n12431,n12435,n12407 );
   nand U12428 ( n12435,n10728,n12592 );
   nand U12429 ( n12517,n12593,n11008 );
   nand U12430 ( n11008,n10987,n11978 );
   not U12431 ( n10987,n11877 );
   nand U12432 ( n11877,n11979,n11980 );
   not U12433 ( n11980,n12264 );
   nor U12434 ( n12264,n11368,n12594 );
   nand U12435 ( n12593,n12595,n12596,n12511 );
   and U12436 ( n12511,n12597,n12598 );
   nand U12437 ( n12598,n12599,n11527 );
   or U12438 ( n12597,n11068,n11527 );
   nand U12439 ( n12596,n11527,n11068,n12600 );
   nand U12440 ( n11068,n12532,n10697 );
   nand U12441 ( n12595,n12513,n12493 );
   not U12442 ( n12493,n12600 );
   nand U12443 ( n12600,n11069,n12601 );
   nand U12444 ( n12601,n12515,n11071,n12419 );
   not U12445 ( n12419,n12418 );
   nand U12446 ( n12418,n11072,n12602 );
   nand U12447 ( n12602,n12405,n11088 );
   nand U12448 ( n11088,n10475,n10731 );
   nand U12449 ( n12405,n11150,n12603 );
   nand U12450 ( n12603,n12390,n11089 );
   nand U12451 ( n11089,n10747,n10478 );
   and U12452 ( n12390,n12604,n12605 );
   nand U12453 ( n12605,n11149,n12606 );
   nand U12454 ( n12606,n11080,n12607 );
   nand U12455 ( n12607,n11084,n12377 );
   not U12456 ( n11084,n12326 );
   nand U12457 ( n12326,n10780,n10487 );
   nor U12458 ( n11080,n12356,n12608 );
   nor U12459 ( n12608,n11465,n10745 );
   nor U12460 ( n12356,n10770,n10759 );
   nand U12461 ( n12604,n12323,n11087,n12377,n11149 );
   nand U12462 ( n11149,n11465,n10745 );
   not U12463 ( n11465,n10760 );
   nand U12464 ( n12377,n10770,n10759 );
   not U12465 ( n10770,n12357 );
   nand U12466 ( n11087,n12349,n11448 );
   not U12467 ( n11448,n10780 );
   nor U12468 ( n12323,n11094,n12609 );
   and U12469 ( n12609,n12299,n11086 );
   nand U12470 ( n11086,n10490,n12297 );
   nand U12471 ( n12299,n11096,n12610 );
   nand U12472 ( n12610,n11098,n12267 );
   nand U12473 ( n12267,n12611,n12612 );
   nand U12474 ( n12612,n11147,n12613 );
   or U12475 ( n12613,n12237,n11146 );
   nand U12476 ( n12611,n11146,n12237 );
   nand U12477 ( n12237,n11100,n12614 );
   nand U12478 ( n12614,n11103,n12223 );
   nand U12479 ( n12223,n12615,n11106 );
   nand U12480 ( n11106,n11265,n10822 );
   nand U12481 ( n12615,n12616,n11104,n11107 );
   and U12482 ( n11107,n12193,n12617 );
   nand U12483 ( n12617,n12618,n11110 );
   not U12484 ( n12618,n12165 );
   nand U12485 ( n12165,n12164,n10508 );
   nand U12486 ( n12193,n12188,n10505 );
   nand U12487 ( n11104,n10834,n10502 );
   nand U12488 ( n12616,n11111,n11110,n12166 );
   not U12489 ( n12166,n12163 );
   nand U12490 ( n12163,n12619,n12620 );
   nand U12491 ( n12620,n11138,n12135 );
   nand U12492 ( n12135,n12621,n11120 );
   nand U12493 ( n11120,n11425,n10888 );
   nand U12494 ( n12621,n12111,n12112,n11134 );
   nand U12495 ( n11134,n10514,n10874 );
   nand U12496 ( n12112,n12046,n11117,n11139 );
   not U12497 ( n11139,n11130 );
   nand U12498 ( n11130,n12064,n12091 );
   nand U12499 ( n12091,n11340,n10901 );
   nand U12500 ( n12046,n12622,n12623,n12624 );
   nand U12501 ( n12624,n12031,n12036 );
   not U12502 ( n12031,n11144 );
   nand U12503 ( n12623,n12625,n10526 );
   nand U12504 ( n12625,n10924,n11144 );
   nand U12505 ( n11144,n10936,n10529 );
   nand U12506 ( n12622,n11140,n12029 );
   nand U12507 ( n12029,n11145,n11143,n12626 );
   or U12508 ( n12626,n11127,n11922 );
   not U12509 ( n11922,n11924 );
   nand U12510 ( n11924,n12627,n12628 );
   nand U12511 ( n12628,n10984,n12629 );
   or U12512 ( n12629,n11132,n10541 );
   nand U12513 ( n12627,n11132,n10541 );
   nand U12514 ( n11132,n11882,n11875 );
   nand U12515 ( n11875,n12588,n10544 );
   nand U12516 ( n11882,n11876,n11874 );
   nand U12517 ( n11874,n10995,n10983 );
   not U12518 ( n11876,n11880 );
   nand U12519 ( n11880,n12630,n12631 );
   nand U12520 ( n12631,n12632,n11379 );
   nand U12521 ( n12632,n10547,n11851 );
   or U12522 ( n12630,n11851,n10547 );
   nand U12523 ( n11127,n11972,n11945,n11925 );
   nand U12524 ( n11925,n10958,n11386 );
   nand U12525 ( n11143,n12589,n10532 );
   not U12526 ( n12589,n10947 );
   nand U12527 ( n11145,n12633,n11972 );
   nand U12528 ( n11972,n10935,n10947 );
   nand U12529 ( n12633,n11946,n12634 );
   nand U12530 ( n12634,n12635,n11945 );
   nand U12531 ( n11945,n11404,n11919 );
   not U12532 ( n12635,n11926 );
   nand U12533 ( n11926,n10970,n10538 );
   nand U12534 ( n11946,n10957,n10535 );
   not U12535 ( n11140,n11129 );
   nand U12536 ( n11129,n12028,n12636 );
   nand U12537 ( n12636,n10914,n10924 );
   nand U12538 ( n12028,n11413,n11961 );
   nand U12539 ( n12111,n12637,n11117 );
   nand U12540 ( n11117,n11430,n10872 );
   nand U12541 ( n12637,n11123,n12638 );
   nand U12542 ( n12638,n11137,n12064 );
   nand U12543 ( n12064,n10887,n11419 );
   nor U12544 ( n11137,n11340,n10901 );
   not U12545 ( n11340,n10913 );
   and U12546 ( n11123,n12065,n12639 );
   nand U12547 ( n12639,n10889,n10517 );
   nand U12548 ( n12065,n10900,n10520 );
   nand U12549 ( n11138,n11116,n10511 );
   nand U12550 ( n12619,n10873,n10861 );
   nand U12551 ( n11110,n10844,n10835 );
   nand U12552 ( n11111,n12123,n10852 );
   nand U12553 ( n11103,n10821,n10499 );
   nand U12554 ( n11100,n10808,n11270 );
   not U12555 ( n11270,n10821 );
   nand U12556 ( n11098,n12265,n10493 );
   nand U12557 ( n11096,n10798,n12236 );
   not U12558 ( n10798,n12265 );
   nor U12559 ( n11094,n12297,n10490 );
   nand U12560 ( n11150,n10726,n11470 );
   not U12561 ( n11470,n10747 );
   nand U12562 ( n11071,n10715,n10728 );
   not U12563 ( n10715,n12592 );
   nand U12564 ( n11069,n12515,n12640 );
   nand U12565 ( n12640,n12641,n12437 );
   nand U12566 ( n12437,n12592,n10472 );
   nand U12567 ( n12641,n12469,n10469 );
   nand U12568 ( n12515,n12416,n10705 );
   not U12569 ( n10705,n12469 );
   nor U12570 ( n12513,n11527,n12599 );
   not U12571 ( n12599,n11065 );
   nand U12572 ( n11065,n12496,n10466 );
   xor U12573 ( n11527,n10463,n10688 );
   not U12574 ( n10688,n11064 );
   nand U12575 ( n11064,n12642,n12643,n12644 );
   nand U12576 ( n12643,n11812,n12645 );
   or U12577 ( n12642,n11812,n11795 );
   nand U12578 ( n12516,n10781,n10466 );
   not U12579 ( n10781,n10727 );
   nand U12580 ( n12648,n11835,n10679 );
   not U12581 ( n10679,n11059 );
   nand U12582 ( n11059,n12650,n12651,n12644 );
   or U12583 ( n12651,n11808,p1_datao_reg_30_ );
   or U12584 ( n12650,n11804,n11812 );
   nand U12585 ( n12647,p2_reg2_reg_30_,n11836 );
   and U12586 ( n12649,n12503,n12654 );
   or U12587 ( n12654,n10672,n11836 );
   nand U12588 ( n10672,n12520,n10457,n12499 );
   nand U12589 ( n10457,n12655,n12656,n12657,n12524 );
   nand U12590 ( n12657,p2_reg2_reg_31_,n12525 );
   nand U12591 ( n12656,p2_reg1_reg_31_,n12526 );
   nand U12592 ( n12655,p2_reg0_reg_31_,n12527 );
   nand U12593 ( n12520,n12644,n12658 );
   nand U12594 ( n12658,n12659,n12660 );
   nand U12595 ( n12503,n11856,n12661 );
   nand U12596 ( n11834,n12662,n11837 );
   nand U12597 ( n12653,n11835,n10674 );
   nand U12598 ( n10674,n12663,n12664 );
   nand U12599 ( n12664,n11811,n12665 );
   nand U12600 ( n12663,n12666,p1_datao_reg_31_ );
   nand U12601 ( n12652,p2_reg2_reg_31_,n11836 );
   nand U12602 ( n12668,n12669,n12670 );
   nand U12603 ( n12670,n12671,n12672,n10649 );
   nand U12604 ( n12672,n12673,n10665 );
   nand U12605 ( n12673,n10666,n12674 );
   nand U12606 ( n12674,n12675,n10661,n11165 );
   nand U12607 ( n12675,n12508,n11030 );
   nand U12608 ( n12671,n10653,n12676 );
   nand U12609 ( n12676,n10667,n10655 );
   nand U12610 ( n10667,n12677,n12678 );
   nand U12611 ( n12677,n12507,n11161 );
   nor U12612 ( n12682,n12683,n12684,n12685 );
   and U12613 ( n12685,p2_addr_reg_19_,n12686 );
   nor U12614 ( n12684,n10662,n12687 );
   nand U12615 ( n12681,n12688,n12689,n12690 );
   nand U12616 ( n12689,n12691,n12692,n12693 );
   not U12617 ( n12693,n12694 );
   nand U12618 ( n12691,p2_reg2_reg_18_,n12695 );
   nand U12619 ( n12688,n12696,n12695,n12694 );
   or U12620 ( n12695,n12697,n12698 );
   nand U12621 ( n12696,n12692,n12699 );
   nand U12622 ( n12692,n12698,n12697 );
   nand U12623 ( n12680,n12700,n12701 );
   xor U12624 ( n12700,n12702,n12703 );
   nand U12625 ( n12703,n12704,n12705 );
   nand U12626 ( n12705,n12706,n12707 );
   or U12627 ( n12707,n12708,n12709 );
   nand U12628 ( n12704,n12709,n12708 );
   nand U12629 ( n12702,n12710,n12711 );
   nand U12630 ( n12711,n12712,n11159 );
   nand U12631 ( n12710,n12694,n12713 );
   xor U12632 ( n12694,p2_reg2_reg_19_,n12508 );
   nand U12633 ( n12679,n12714,n12715,n12716 );
   nand U12634 ( n12715,n12717,n12718,n12719 );
   not U12635 ( n12719,n12712 );
   nand U12636 ( n12717,p2_reg1_reg_18_,n12720 );
   nand U12637 ( n12714,n12721,n12720,n12712 );
   xor U12638 ( n12712,p2_reg1_reg_19_,n12508 );
   or U12639 ( n12720,n12722,n12698 );
   nand U12640 ( n12721,n12718,n12723 );
   nand U12641 ( n12718,n12698,n12722 );
   nand U12642 ( n12728,n12687,n12729,n12730,n12731 );
   nand U12643 ( n12731,n12732,n12701 );
   nand U12644 ( n12730,n12716,n12733 );
   xor U12645 ( n12733,n12722,n12723 );
   nand U12646 ( n12729,n12690,n12734 );
   xor U12647 ( n12734,n12697,n12699 );
   not U12648 ( n12706,n12698 );
   nand U12649 ( n12726,n12735,n12698 );
   nand U12650 ( n12735,n12736,n12737,n12738 );
   nand U12651 ( n12738,n12739,n12690 );
   xor U12652 ( n12739,p2_reg2_reg_18_,n12697 );
   nand U12653 ( n12697,n12740,n12741 );
   nand U12654 ( n12741,p2_reg2_reg_17_,n12742 );
   or U12655 ( n12742,n12743,n12744 );
   nand U12656 ( n12740,n12743,n12744 );
   or U12657 ( n12737,n12745,n12732 );
   xor U12658 ( n12732,n12709,n12708 );
   nand U12659 ( n12708,n12746,n12747 );
   nand U12660 ( n12747,n12748,n12749 );
   or U12661 ( n12749,n12750,n12751 );
   nand U12662 ( n12746,n12751,n12750 );
   nand U12663 ( n12709,n12752,n12753 );
   nand U12664 ( n12753,n12713,n12699 );
   not U12665 ( n12699,p2_reg2_reg_18_ );
   nand U12666 ( n12752,n11159,n12723 );
   not U12667 ( n12723,p2_reg1_reg_18_ );
   nand U12668 ( n12736,n12754,n12716 );
   xor U12669 ( n12754,p2_reg1_reg_18_,n12722 );
   nand U12670 ( n12722,n12755,n12756 );
   nand U12671 ( n12756,p2_reg1_reg_17_,n12757 );
   or U12672 ( n12757,n12758,n12744 );
   nand U12673 ( n12755,n12758,n12744 );
   nand U12674 ( n12725,p2_addr_reg_18_,n12686 );
   nand U12675 ( n12724,p2_reg3_reg_18_,p2_u3151 );
   nand U12676 ( n12763,n12687,n12764,n12765,n12766 );
   nand U12677 ( n12766,n12767,n12701 );
   nand U12678 ( n12765,n12716,n12768 );
   xor U12679 ( n12768,n12758,n12769 );
   nand U12680 ( n12764,n12690,n12770 );
   xor U12681 ( n12770,n12743,n12771 );
   not U12682 ( n12748,n12744 );
   nand U12683 ( n12761,n12772,n12744 );
   nand U12684 ( n12772,n12773,n12774,n12775 );
   nand U12685 ( n12775,n12776,n12690 );
   xor U12686 ( n12776,p2_reg2_reg_17_,n12743 );
   nand U12687 ( n12743,n12777,n12778 );
   nand U12688 ( n12778,p2_reg2_reg_16_,n12779 );
   or U12689 ( n12779,n12780,n12781 );
   nand U12690 ( n12777,n12781,n12780 );
   or U12691 ( n12774,n12745,n12767 );
   xor U12692 ( n12767,n12751,n12750 );
   nand U12693 ( n12750,n12782,n12783 );
   nand U12694 ( n12782,n12784,n12785 );
   nand U12695 ( n12751,n12786,n12787 );
   nand U12696 ( n12787,n12713,n12771 );
   not U12697 ( n12771,p2_reg2_reg_17_ );
   nand U12698 ( n12786,n11159,n12769 );
   not U12699 ( n12769,p2_reg1_reg_17_ );
   nand U12700 ( n12773,n12788,n12716 );
   xor U12701 ( n12788,p2_reg1_reg_17_,n12758 );
   nand U12702 ( n12758,n12789,n12790 );
   nand U12703 ( n12790,p2_reg1_reg_16_,n12791 );
   or U12704 ( n12791,n12792,n12781 );
   nand U12705 ( n12789,n12781,n12792 );
   nand U12706 ( n12760,p2_addr_reg_17_,n12686 );
   nand U12707 ( n12759,p2_reg3_reg_17_,p2_u3151 );
   nor U12708 ( n12795,n12796,n12797,n12798 );
   nor U12709 ( n12798,n12799,n12781 );
   nor U12710 ( n12799,n12800,n12801,n12802 );
   nor U12711 ( n12802,n12803,n12804 );
   xor U12712 ( n12803,p2_reg2_reg_16_,n12780 );
   nor U12713 ( n12801,n12805,n12806 );
   xor U12714 ( n12805,p2_reg1_reg_16_,n12792 );
   nor U12715 ( n12797,n12807,n12808 );
   nor U12716 ( n12807,n12809,n12810 );
   nor U12717 ( n12810,n12804,n12811 );
   xor U12718 ( n12811,n12780,n12207 );
   nand U12719 ( n12780,n12812,n12813 );
   nand U12720 ( n12813,p2_reg2_reg_15_,n12814 );
   or U12721 ( n12814,n12815,n12816 );
   nand U12722 ( n12812,n12815,n12816 );
   nor U12723 ( n12809,n12806,n12817 );
   xor U12724 ( n12817,n12792,n12818 );
   nand U12725 ( n12792,n12819,n12820 );
   nand U12726 ( n12820,p2_reg1_reg_15_,n12821 );
   or U12727 ( n12821,n12822,n12816 );
   nand U12728 ( n12819,n12822,n12816 );
   nand U12729 ( n12794,n12701,n12823 );
   nand U12730 ( n12823,n12824,n12825 );
   nand U12731 ( n12825,n12785,n12783,n12784 );
   and U12732 ( n12784,n12826,n12827 );
   or U12733 ( n12827,n12828,n12808 );
   nand U12734 ( n12783,n12808,n12828 );
   not U12735 ( n12808,n12781 );
   nand U12736 ( n12785,n12829,n12830 );
   nand U12737 ( n12824,n12831,n12829,n12832 );
   xor U12738 ( n12832,n12781,n12828 );
   nand U12739 ( n12828,n12833,n12834 );
   nand U12740 ( n12834,n12713,n12207 );
   not U12741 ( n12207,p2_reg2_reg_16_ );
   nand U12742 ( n12833,n11159,n12818 );
   not U12743 ( n12818,p2_reg1_reg_16_ );
   nand U12744 ( n12831,n12835,n12826 );
   nand U12745 ( n12826,n12836,n12816 );
   nand U12746 ( n12793,p2_addr_reg_16_,n12686 );
   nor U12747 ( n12840,n12841,n12842 );
   nor U12748 ( n12842,n12843,n12844 );
   nor U12749 ( n12841,n12829,n12835,n12745 );
   nand U12750 ( n12829,n12845,n12846 );
   nand U12751 ( n12839,p2_reg3_reg_15_,p2_u3151 );
   nand U12752 ( n12838,n12847,n12816 );
   nand U12753 ( n12847,n12848,n12849,n12850 );
   nand U12754 ( n12850,n12851,n12690 );
   xor U12755 ( n12851,p2_reg2_reg_15_,n12815 );
   nand U12756 ( n12849,n12852,n12701 );
   xor U12757 ( n12852,n12835,n12836 );
   nand U12758 ( n12848,n12853,n12716 );
   xor U12759 ( n12853,p2_reg1_reg_15_,n12822 );
   nand U12760 ( n12837,n12845,n12854 );
   nand U12761 ( n12854,n12687,n12855,n12856,n12857 );
   nand U12762 ( n12857,n12836,n12701,n12835 );
   not U12763 ( n12835,n12830 );
   nand U12764 ( n12830,n12858,n12859 );
   nand U12765 ( n12859,n12860,n12861 );
   nand U12766 ( n12861,n12862,n12863 );
   nand U12767 ( n12858,n12864,n12865 );
   not U12768 ( n12836,n12846 );
   nand U12769 ( n12846,n12866,n12867 );
   nand U12770 ( n12867,n12713,n12187 );
   nand U12771 ( n12866,n11159,n12868 );
   nand U12772 ( n12856,n12716,n12869 );
   xor U12773 ( n12869,n12822,n12868 );
   not U12774 ( n12868,p2_reg1_reg_15_ );
   nand U12775 ( n12822,n12870,n12871 );
   nand U12776 ( n12871,p2_reg1_reg_14_,n12872 );
   or U12777 ( n12872,n12873,n12865 );
   nand U12778 ( n12870,n12865,n12873 );
   nand U12779 ( n12855,n12690,n12874 );
   xor U12780 ( n12874,n12815,n12187 );
   not U12781 ( n12187,p2_reg2_reg_15_ );
   nand U12782 ( n12815,n12875,n12876 );
   nand U12783 ( n12876,p2_reg2_reg_14_,n12877 );
   or U12784 ( n12877,n12878,n12865 );
   nand U12785 ( n12875,n12865,n12878 );
   not U12786 ( n12845,n12816 );
   nand U12787 ( n12882,n12865,n12883 );
   nand U12788 ( n12883,n12884,n12885,n12886 );
   nand U12789 ( n12886,n12887,n12690 );
   xor U12790 ( n12887,p2_reg2_reg_14_,n12878 );
   nand U12791 ( n12885,n12701,n12888 );
   xor U12792 ( n12888,n12863,n12860 );
   nand U12793 ( n12884,n12889,n12716 );
   xor U12794 ( n12889,p2_reg1_reg_14_,n12873 );
   nand U12795 ( n12881,n12862,n12890 );
   nand U12796 ( n12890,n12687,n12891,n12892,n12893 );
   nand U12797 ( n12893,n12894,n12701 );
   xor U12798 ( n12894,n12864,n12860 );
   and U12799 ( n12860,n12895,n12896 );
   nand U12800 ( n12896,n12897,n12898 );
   or U12801 ( n12898,n12899,n12900 );
   nand U12802 ( n12895,n12900,n12899 );
   not U12803 ( n12864,n12863 );
   nand U12804 ( n12863,n12901,n12902 );
   nand U12805 ( n12902,n12713,n12903 );
   nand U12806 ( n12901,n11159,n12904 );
   nand U12807 ( n12892,n12716,n12905 );
   xor U12808 ( n12905,n12873,n12904 );
   not U12809 ( n12904,p2_reg1_reg_14_ );
   nand U12810 ( n12873,n12906,n12907 );
   nand U12811 ( n12907,p2_reg1_reg_13_,n12908 );
   or U12812 ( n12908,n12909,n12910 );
   nand U12813 ( n12906,n12909,n12910 );
   nand U12814 ( n12891,n12690,n12911 );
   xor U12815 ( n12911,n12878,n12903 );
   not U12816 ( n12903,p2_reg2_reg_14_ );
   nand U12817 ( n12878,n12912,n12913 );
   nand U12818 ( n12913,p2_reg2_reg_13_,n12914 );
   or U12819 ( n12914,n12915,n12910 );
   nand U12820 ( n12912,n12915,n12910 );
   nand U12821 ( n12880,p2_addr_reg_14_,n12686 );
   nand U12822 ( n12879,p2_reg3_reg_14_,p2_u3151 );
   nand U12823 ( n12920,n12687,n12921,n12922,n12923 );
   nand U12824 ( n12923,n12924,n12701 );
   nand U12825 ( n12922,n12716,n12925 );
   xor U12826 ( n12925,n12909,n12926 );
   nand U12827 ( n12921,n12690,n12927 );
   xor U12828 ( n12927,n12915,n12928 );
   nand U12829 ( n12918,n12929,n12910 );
   nand U12830 ( n12929,n12930,n12931,n12932 );
   nand U12831 ( n12932,n12933,n12690 );
   xor U12832 ( n12933,p2_reg2_reg_13_,n12915 );
   nand U12833 ( n12915,n12934,n12935 );
   nand U12834 ( n12935,p2_reg2_reg_12_,n12936 );
   or U12835 ( n12936,n12937,n12938 );
   nand U12836 ( n12934,n12938,n12937 );
   or U12837 ( n12931,n12745,n12924 );
   xor U12838 ( n12924,n12900,n12899 );
   nand U12839 ( n12899,n12939,n12940 );
   nand U12840 ( n12940,n12941,n12942 );
   nand U12841 ( n12942,n12943,n12944 );
   or U12842 ( n12939,n12944,n12943 );
   nand U12843 ( n12900,n12945,n12946 );
   nand U12844 ( n12946,n12713,n12928 );
   not U12845 ( n12928,p2_reg2_reg_13_ );
   nand U12846 ( n12945,n11159,n12926 );
   not U12847 ( n12926,p2_reg1_reg_13_ );
   nand U12848 ( n12930,n12947,n12716 );
   xor U12849 ( n12947,p2_reg1_reg_13_,n12909 );
   nand U12850 ( n12909,n12948,n12949 );
   nand U12851 ( n12949,p2_reg1_reg_12_,n12950 );
   or U12852 ( n12950,n12951,n12938 );
   nand U12853 ( n12948,n12938,n12951 );
   nand U12854 ( n12917,p2_addr_reg_13_,n12686 );
   nand U12855 ( n12916,p2_reg3_reg_13_,p2_u3151 );
   nand U12856 ( n12955,n12938,n12956 );
   nand U12857 ( n12956,n12957,n12958,n12959 );
   nand U12858 ( n12959,n12960,n12690 );
   xor U12859 ( n12960,p2_reg2_reg_12_,n12937 );
   nand U12860 ( n12958,n12961,n12701 );
   xor U12861 ( n12961,n12944,n12962 );
   nand U12862 ( n12957,n12963,n12716 );
   xor U12863 ( n12963,p2_reg1_reg_12_,n12951 );
   nand U12864 ( n12954,n12941,n12964 );
   nand U12865 ( n12964,n12687,n12965,n12966,n12967 );
   nand U12866 ( n12967,n12701,n12968 );
   xor U12867 ( n12968,n12944,n12943 );
   not U12868 ( n12943,n12962 );
   nand U12869 ( n12962,n12969,n12970 );
   nand U12870 ( n12970,n12713,n12103 );
   nand U12871 ( n12969,n11159,n12971 );
   nand U12872 ( n12944,n12972,n12973 );
   nand U12873 ( n12973,n12974,n12975,n12976,n12977 );
   nand U12874 ( n12974,n12978,n12979 );
   nand U12875 ( n12972,n12980,n12977 );
   nand U12876 ( n12980,n12981,n12982 );
   nand U12877 ( n12982,n12975,n12983,n12984 );
   nand U12878 ( n12966,n12716,n12985 );
   xor U12879 ( n12985,n12951,n12971 );
   not U12880 ( n12971,p2_reg1_reg_12_ );
   nand U12881 ( n12951,n12986,n12987 );
   nand U12882 ( n12987,p2_reg1_reg_11_,n12988 );
   or U12883 ( n12988,n12989,n12990 );
   nand U12884 ( n12986,n12989,n12990 );
   nand U12885 ( n12965,n12690,n12991 );
   xor U12886 ( n12991,n12937,n12103 );
   not U12887 ( n12103,p2_reg2_reg_12_ );
   nand U12888 ( n12937,n12992,n12993 );
   nand U12889 ( n12993,p2_reg2_reg_11_,n12994 );
   or U12890 ( n12994,n12995,n12990 );
   nand U12891 ( n12992,n12995,n12990 );
   not U12892 ( n12941,n12938 );
   nand U12893 ( n12953,p2_addr_reg_12_,n12686 );
   nand U12894 ( n12952,p2_reg3_reg_12_,p2_u3151 );
   nor U12895 ( n12998,n12999,n13000,n13001 );
   nor U12896 ( n13001,n13002,n13003 );
   nor U12897 ( n13003,n13004,n13005 );
   nor U12898 ( n13005,n12804,n13006 );
   xor U12899 ( n13006,n12995,n12092 );
   nor U12900 ( n13004,n12806,n13007 );
   xor U12901 ( n13007,n12989,n13008 );
   nor U12902 ( n13000,n13009,n12990 );
   nor U12903 ( n13009,n12800,n13010,n13011 );
   nor U12904 ( n13011,n13012,n12804 );
   xor U12905 ( n13012,p2_reg2_reg_11_,n12995 );
   nand U12906 ( n12995,n13013,n13014 );
   nand U12907 ( n13014,p2_reg2_reg_10_,n13015 );
   or U12908 ( n13015,n13016,n13017 );
   nand U12909 ( n13013,n13017,n13016 );
   nor U12910 ( n13010,n13018,n12806 );
   xor U12911 ( n13018,p2_reg1_reg_11_,n12989 );
   nand U12912 ( n12989,n13019,n13020 );
   nand U12913 ( n13020,p2_reg1_reg_10_,n13021 );
   or U12914 ( n13021,n13022,n13017 );
   nand U12915 ( n13019,n13017,n13022 );
   nand U12916 ( n12997,n12701,n13023 );
   nand U12917 ( n13023,n13024,n13025 );
   nand U12918 ( n13025,n13026,n12977,n12981 );
   and U12919 ( n12981,n13027,n13028 );
   or U12920 ( n13028,n13029,n13002 );
   nand U12921 ( n12977,n13002,n13029 );
   not U12922 ( n13002,n12990 );
   nand U12923 ( n13026,n13030,n12975 );
   nand U12924 ( n13024,n13031,n12975,n13032 );
   xor U12925 ( n13032,n12990,n13029 );
   nand U12926 ( n13029,n13033,n13034 );
   nand U12927 ( n13034,n12713,n12092 );
   not U12928 ( n12092,p2_reg2_reg_11_ );
   nand U12929 ( n13033,n11159,n13008 );
   not U12930 ( n13008,p2_reg1_reg_11_ );
   nand U12931 ( n13031,n13027,n13035 );
   nand U12932 ( n13027,n13036,n13017 );
   nand U12933 ( n12996,p2_addr_reg_11_,n12686 );
   nor U12934 ( n13040,n13041,n13042 );
   nor U12935 ( n13042,n12843,n13043 );
   nor U12936 ( n13041,n12975,n12745,n13035 );
   nand U12937 ( n12975,n13044,n13045 );
   nand U12938 ( n13039,p2_reg3_reg_10_,p2_u3151 );
   nand U12939 ( n13038,n13017,n13046 );
   nand U12940 ( n13046,n13047,n13048,n13049 );
   nand U12941 ( n13049,n13050,n12690 );
   xor U12942 ( n13050,p2_reg2_reg_10_,n13016 );
   nand U12943 ( n13048,n12701,n13051 );
   xor U12944 ( n13051,n13030,n13045 );
   not U12945 ( n13030,n13035 );
   nand U12946 ( n13047,n13052,n12716 );
   xor U12947 ( n13052,p2_reg1_reg_10_,n13022 );
   nand U12948 ( n13037,n13044,n13053 );
   nand U12949 ( n13053,n12687,n13054,n13055,n13056 );
   nand U12950 ( n13056,n13036,n13035,n12701 );
   nand U12951 ( n13035,n13057,n13058 );
   nand U12952 ( n13058,n12978,n13059 );
   nand U12953 ( n13059,n12984,n12976 );
   or U12954 ( n13057,n12976,n12984 );
   not U12955 ( n13036,n13045 );
   nand U12956 ( n13045,n13060,n13061 );
   nand U12957 ( n13061,n12713,n13062 );
   nand U12958 ( n13060,n11159,n13063 );
   nand U12959 ( n13055,n12716,n13064 );
   xor U12960 ( n13064,n13022,n13063 );
   not U12961 ( n13063,p2_reg1_reg_10_ );
   nand U12962 ( n13022,n13065,n13066 );
   nand U12963 ( n13066,p2_reg1_reg_9_,n13067 );
   or U12964 ( n13067,n13068,n12983 );
   nand U12965 ( n13065,n13068,n12983 );
   nand U12966 ( n13054,n12690,n13069 );
   xor U12967 ( n13069,n13016,n13062 );
   not U12968 ( n13062,p2_reg2_reg_10_ );
   nand U12969 ( n13016,n13070,n13071 );
   nand U12970 ( n13071,p2_reg2_reg_9_,n13072 );
   or U12971 ( n13072,n13073,n12983 );
   nand U12972 ( n13070,n13073,n12983 );
   nand U12973 ( n13078,n12687,n13079,n13080,n13081 );
   nand U12974 ( n13081,n12701,n13082 );
   xor U12975 ( n13082,n12976,n12984 );
   not U12976 ( n12984,n12979 );
   nand U12977 ( n13080,n12716,n13083 );
   xor U12978 ( n13083,n13068,n13084 );
   nand U12979 ( n13079,n12690,n13085 );
   xor U12980 ( n13085,n13073,n13086 );
   not U12981 ( n12978,n12983 );
   nand U12982 ( n13076,n13087,n12983 );
   nand U12983 ( n13087,n13088,n13089,n13090 );
   nand U12984 ( n13090,n13091,n12690 );
   xor U12985 ( n13091,p2_reg2_reg_9_,n13073 );
   nand U12986 ( n13073,n13092,n13093 );
   nand U12987 ( n13093,p2_reg2_reg_8_,n13094 );
   or U12988 ( n13094,n13095,n13096 );
   nand U12989 ( n13092,n13096,n13095 );
   nand U12990 ( n13089,n13097,n12701 );
   xor U12991 ( n13097,n12976,n12979 );
   nand U12992 ( n12979,n13098,n13099 );
   nand U12993 ( n13099,n12713,n13086 );
   not U12994 ( n13086,p2_reg2_reg_9_ );
   nand U12995 ( n13098,n11159,n13084 );
   not U12996 ( n13084,p2_reg1_reg_9_ );
   nand U12997 ( n12976,n13100,n13101 );
   nand U12998 ( n13101,n13102,n13103 );
   nand U12999 ( n13102,n13104,n13105 );
   nand U13000 ( n13088,n13106,n12716 );
   xor U13001 ( n13106,p2_reg1_reg_9_,n13068 );
   nand U13002 ( n13068,n13107,n13108 );
   nand U13003 ( n13108,p2_reg1_reg_8_,n13109 );
   or U13004 ( n13109,n13110,n13096 );
   nand U13005 ( n13107,n13096,n13110 );
   nand U13006 ( n13075,p2_addr_reg_9_,n12686 );
   nand U13007 ( n13074,p2_reg3_reg_9_,p2_u3151 );
   nor U13008 ( n13114,n13115,n13116 );
   nor U13009 ( n13116,n12843,n13117 );
   nor U13010 ( n13115,n12745,n13118,n13119 );
   nor U13011 ( n13119,n13120,n13121,n13122 );
   and U13012 ( n13122,n13105,n13104 );
   nor U13013 ( n13118,n13123,n13103 );
   nor U13014 ( n13123,n13121,n13105 );
   nand U13015 ( n13113,p2_reg3_reg_8_,p2_u3151 );
   nand U13016 ( n13112,n13096,n13124 );
   nand U13017 ( n13124,n13125,n13126,n13127 );
   nand U13018 ( n13127,n13128,n12690 );
   xor U13019 ( n13128,p2_reg2_reg_8_,n13095 );
   nand U13020 ( n13126,n12701,n13100,n13120 );
   not U13021 ( n13120,n13103 );
   nand U13022 ( n13103,n13129,n13130 );
   nand U13023 ( n13130,n13131,n13132 );
   nand U13024 ( n13132,n13133,n13134 );
   not U13025 ( n13131,n13135 );
   not U13026 ( n13100,n13121 );
   nor U13027 ( n13121,n13105,n13104 );
   nand U13028 ( n13105,n13136,n13137 );
   nand U13029 ( n13137,n12713,n13138 );
   nand U13030 ( n13136,n11159,n13139 );
   nand U13031 ( n13125,n13140,n12716 );
   xor U13032 ( n13140,p2_reg1_reg_8_,n13110 );
   nand U13033 ( n13111,n13104,n13141 );
   nand U13034 ( n13141,n13142,n13143,n12687 );
   nand U13035 ( n13143,n12716,n13144 );
   xor U13036 ( n13144,n13110,n13139 );
   not U13037 ( n13139,p2_reg1_reg_8_ );
   nand U13038 ( n13110,n13145,n13146 );
   nand U13039 ( n13146,p2_reg1_reg_7_,n13147 );
   or U13040 ( n13147,n13148,n13149 );
   nand U13041 ( n13145,n13148,n13149 );
   nand U13042 ( n13142,n12690,n13150 );
   xor U13043 ( n13150,n13095,n13138 );
   not U13044 ( n13138,p2_reg2_reg_8_ );
   nand U13045 ( n13095,n13151,n13152 );
   nand U13046 ( n13152,p2_reg2_reg_7_,n13153 );
   or U13047 ( n13153,n13154,n13149 );
   nand U13048 ( n13151,n13154,n13149 );
   not U13049 ( n13104,n13096 );
   nor U13050 ( n13158,n13159,n13160 );
   nor U13051 ( n13160,n12843,n13161 );
   nor U13052 ( n13159,n13129,n13135,n12745 );
   or U13053 ( n13129,n13134,n13133 );
   nand U13054 ( n13157,p2_reg3_reg_7_,p2_u3151 );
   nand U13055 ( n13156,n13133,n13162 );
   nand U13056 ( n13162,n12687,n13163,n13164,n13165 );
   nand U13057 ( n13165,n13166,n12701 );
   xor U13058 ( n13166,n13134,n13135 );
   nand U13059 ( n13164,n12716,n13167 );
   xor U13060 ( n13167,n13148,n13168 );
   nand U13061 ( n13163,n12690,n13169 );
   xor U13062 ( n13169,n13154,n11991 );
   not U13063 ( n13133,n13149 );
   nand U13064 ( n13155,n13170,n13149 );
   nand U13065 ( n13170,n13171,n13172,n13173 );
   nand U13066 ( n13173,n13174,n12690 );
   xor U13067 ( n13174,p2_reg2_reg_7_,n13154 );
   nand U13068 ( n13154,n13175,n13176 );
   nand U13069 ( n13176,p2_reg2_reg_6_,n13177 );
   or U13070 ( n13177,n13178,n13179 );
   nand U13071 ( n13175,n13179,n13178 );
   nand U13072 ( n13172,n13134,n13135,n12701 );
   nand U13073 ( n13135,n13180,n13181 );
   not U13074 ( n13180,n13182 );
   nand U13075 ( n13134,n13183,n13184 );
   nand U13076 ( n13184,n12713,n11991 );
   not U13077 ( n11991,p2_reg2_reg_7_ );
   nand U13078 ( n13183,n11159,n13168 );
   not U13079 ( n13168,p2_reg1_reg_7_ );
   nand U13080 ( n13171,n13185,n12716 );
   xor U13081 ( n13185,p2_reg1_reg_7_,n13148 );
   nand U13082 ( n13148,n13186,n13187 );
   nand U13083 ( n13187,p2_reg1_reg_6_,n13188 );
   or U13084 ( n13188,n13189,n13179 );
   nand U13085 ( n13186,n13179,n13189 );
   nor U13086 ( n13193,n13194,n13195 );
   nor U13087 ( n13195,n12843,n13196 );
   nor U13088 ( n13194,n13197,n12745 );
   nor U13089 ( n13197,n13198,n13199 );
   nor U13090 ( n13199,n13182,n13181 );
   nand U13091 ( n13181,n13200,n13201,n13202 );
   nand U13092 ( n13202,n13203,n13204 );
   nand U13093 ( n13200,n13205,n13179 );
   nor U13094 ( n13198,n13206,n13207,n13208 );
   not U13095 ( n13208,n13203 );
   nor U13096 ( n13207,n13209,n13204 );
   not U13097 ( n13209,n13201 );
   nor U13098 ( n13206,n13210,n13182 );
   nor U13099 ( n13182,n13205,n13179 );
   and U13100 ( n13210,n13179,n13205 );
   nand U13101 ( n13205,n13211,n13212 );
   nand U13102 ( n13212,p2_reg1_reg_6_,n11159 );
   nand U13103 ( n13211,n12713,p2_reg2_reg_6_ );
   nand U13104 ( n13192,p2_reg3_reg_6_,p2_u3151 );
   nand U13105 ( n13191,n13179,n13213 );
   nand U13106 ( n13213,n13214,n13215 );
   nand U13107 ( n13215,n13216,n12716 );
   nand U13108 ( n13214,n13217,n12690 );
   nand U13109 ( n13190,n13218,n13219 );
   nand U13110 ( n13219,n13220,n13221,n12687 );
   or U13111 ( n13221,n12806,n13216 );
   xor U13112 ( n13216,p2_reg1_reg_6_,n13189 );
   nand U13113 ( n13189,n13222,n13223 );
   nand U13114 ( n13223,p2_reg1_reg_5_,n13224 );
   or U13115 ( n13224,n13225,n13226 );
   nand U13116 ( n13222,n13225,n13226 );
   or U13117 ( n13220,n12804,n13217 );
   xor U13118 ( n13217,p2_reg2_reg_6_,n13178 );
   nand U13119 ( n13178,n13227,n13228 );
   nand U13120 ( n13228,p2_reg2_reg_5_,n13229 );
   or U13121 ( n13229,n13230,n13226 );
   nand U13122 ( n13227,n13230,n13226 );
   nand U13123 ( n13235,n13201,n13203 );
   nand U13124 ( n13203,n13236,n13237 );
   nand U13125 ( n13201,n13238,n13226 );
   nand U13126 ( n13233,p2_addr_reg_5_,n12686 );
   nand U13127 ( n13232,p2_reg3_reg_5_,p2_u3151 );
   nor U13128 ( n13231,n13239,n13240 );
   nor U13129 ( n13240,n13236,n13241 );
   nor U13130 ( n13241,n13242,n13243,n13244 );
   nor U13131 ( n13244,n12806,n13245 );
   xor U13132 ( n13245,n13225,n13246 );
   nor U13133 ( n13243,n13204,n13238,n12745 );
   not U13134 ( n13238,n13237 );
   nor U13135 ( n13242,n12804,n13247 );
   xor U13136 ( n13247,n13230,n13248 );
   not U13137 ( n13236,n13226 );
   nor U13138 ( n13239,n13249,n13226 );
   nor U13139 ( n13249,n13250,n13251,n13252,n12800 );
   nor U13140 ( n13252,n13253,n12804 );
   xor U13141 ( n13253,p2_reg2_reg_5_,n13230 );
   nand U13142 ( n13230,n13254,n13255 );
   nand U13143 ( n13255,p2_reg2_reg_4_,n13256 );
   or U13144 ( n13256,n13257,n13258 );
   nand U13145 ( n13254,n13258,n13257 );
   nor U13146 ( n13251,n13259,n12806 );
   xor U13147 ( n13259,p2_reg1_reg_5_,n13225 );
   nand U13148 ( n13225,n13260,n13261 );
   nand U13149 ( n13261,p2_reg1_reg_4_,n13262 );
   or U13150 ( n13262,n13263,n13258 );
   nand U13151 ( n13260,n13258,n13263 );
   nor U13152 ( n13250,n13204,n12745,n13237 );
   nand U13153 ( n13237,n13264,n13265 );
   nand U13154 ( n13265,n12713,n13248 );
   not U13155 ( n13248,p2_reg2_reg_5_ );
   nand U13156 ( n13264,n11159,n13246 );
   not U13157 ( n13246,p2_reg1_reg_5_ );
   nand U13158 ( n13204,n13266,n13267 );
   nand U13159 ( n13266,n13268,n13269 );
   nor U13160 ( n13275,n13276,n13258 );
   nor U13161 ( n13276,n13277,n13278,n13279,n12800 );
   nor U13162 ( n13279,n13280,n12804 );
   xor U13163 ( n13280,p2_reg2_reg_4_,n13257 );
   nor U13164 ( n13278,n13281,n12806 );
   xor U13165 ( n13281,p2_reg1_reg_4_,n13263 );
   nor U13166 ( n13277,n13268,n12745,n13282 );
   nor U13167 ( n13274,n13283,n13284 );
   nor U13168 ( n13283,n13285,n13286,n13287 );
   nor U13169 ( n13287,n12806,n13288 );
   xor U13170 ( n13288,n13263,n13289 );
   nand U13171 ( n13263,n13290,n13291 );
   nand U13172 ( n13291,p2_reg1_reg_3_,n13292 );
   or U13173 ( n13292,n13293,n13294 );
   nand U13174 ( n13290,n13293,n13294 );
   nor U13175 ( n13286,n13268,n13295,n12745 );
   nor U13176 ( n13285,n12804,n13296 );
   xor U13177 ( n13296,n13257,n13297 );
   nand U13178 ( n13257,n13298,n13299 );
   nand U13179 ( n13299,p2_reg2_reg_3_,n13300 );
   or U13180 ( n13300,n13301,n13294 );
   nand U13181 ( n13298,n13301,n13294 );
   nand U13182 ( n13271,n13302,n13268,n12701 );
   nand U13183 ( n13268,n13303,n13304 );
   nand U13184 ( n13304,n13305,n13306 );
   nand U13185 ( n13302,n13269,n13267 );
   nand U13186 ( n13267,n13295,n13258 );
   not U13187 ( n13295,n13282 );
   nand U13188 ( n13269,n13284,n13282 );
   nand U13189 ( n13282,n13307,n13308 );
   nand U13190 ( n13308,n12713,n13297 );
   not U13191 ( n13297,p2_reg2_reg_4_ );
   nand U13192 ( n13307,n11159,n13289 );
   not U13193 ( n13289,p2_reg1_reg_4_ );
   not U13194 ( n13284,n13258 );
   nand U13195 ( n13270,p2_addr_reg_4_,n12686 );
   nor U13196 ( n13314,n13315,n13294 );
   nor U13197 ( n13315,n12800,n13316,n13317 );
   nor U13198 ( n13317,n13318,n12804 );
   xor U13199 ( n13318,p2_reg2_reg_3_,n13301 );
   nor U13200 ( n13316,n13319,n12806 );
   xor U13201 ( n13319,p2_reg1_reg_3_,n13293 );
   nor U13202 ( n13313,n13320,n13321 );
   nor U13203 ( n13321,n13322,n13323,n13324 );
   nor U13204 ( n13324,n12806,n13325 );
   xor U13205 ( n13325,n13293,n13326 );
   nand U13206 ( n13293,n13327,n13328 );
   nand U13207 ( n13328,p2_reg1_reg_2_,n13329 );
   or U13208 ( n13329,n13330,n13331 );
   nand U13209 ( n13327,n13331,n13330 );
   nor U13210 ( n13323,n13306,n13332,n12745 );
   nor U13211 ( n13322,n12804,n13333 );
   xor U13212 ( n13333,n13301,n11909 );
   nand U13213 ( n13301,n13334,n13335 );
   nand U13214 ( n13335,p2_reg2_reg_2_,n13336 );
   or U13215 ( n13336,n13337,n13331 );
   nand U13216 ( n13334,n13331,n13337 );
   nand U13217 ( n13310,n13338,n13339,n12701 );
   nand U13218 ( n13339,n13340,n13341 );
   or U13219 ( n13341,n13342,n13332 );
   nand U13220 ( n13338,n13305,n13303,n13306 );
   not U13221 ( n13306,n13340 );
   nor U13222 ( n13340,n13343,n13344 );
   and U13223 ( n13344,n13345,n13346 );
   nand U13224 ( n13346,n13347,n13348 );
   not U13225 ( n13303,n13332 );
   nor U13226 ( n13332,n13342,n13320 );
   nand U13227 ( n13305,n13320,n13342 );
   nand U13228 ( n13342,n13349,n13350 );
   nand U13229 ( n13350,n12713,n11909 );
   not U13230 ( n11909,p2_reg2_reg_3_ );
   nand U13231 ( n13349,n11159,n13326 );
   not U13232 ( n13326,p2_reg1_reg_3_ );
   nand U13233 ( n13309,p2_addr_reg_3_,n12686 );
   nor U13234 ( n13356,n13357,n13331 );
   nor U13235 ( n13357,n13358,n13359,n13360,n12800 );
   nor U13236 ( n13360,n13361,n12804 );
   xor U13237 ( n13361,p2_reg2_reg_2_,n13337 );
   nor U13238 ( n13359,n13362,n12806 );
   xor U13239 ( n13362,p2_reg1_reg_2_,n13330 );
   nor U13240 ( n13358,n12745,n13363 );
   xor U13241 ( n13363,n13348,n13345 );
   nor U13242 ( n13355,n13364,n13347 );
   nor U13243 ( n13364,n13365,n13366,n13367 );
   nor U13244 ( n13367,n12806,n13368 );
   xor U13245 ( n13368,n13330,n13369 );
   nand U13246 ( n13330,n13370,n13371 );
   nand U13247 ( n13371,p2_reg1_reg_1_,n13372 );
   nand U13248 ( n13372,n13373,n13374 );
   nand U13249 ( n13370,n13375,n13376 );
   nor U13250 ( n13366,n12745,n13345,n13377 );
   not U13251 ( n13377,n13348 );
   nor U13252 ( n13365,n12804,n13378 );
   xor U13253 ( n13378,n13337,n13379 );
   nand U13254 ( n13337,n13380,n13381 );
   nand U13255 ( n13381,p2_reg2_reg_1_,n13382 );
   nand U13256 ( n13382,n13373,n13383 );
   nand U13257 ( n13380,n13384,n13376 );
   nor U13258 ( n13354,p2_state_reg,n11866 );
   not U13259 ( n11866,p2_reg3_reg_2_ );
   nand U13260 ( n13352,n12701,n13345,n13343 );
   nor U13261 ( n13343,n13348,n13347 );
   not U13262 ( n13347,n13331 );
   nand U13263 ( n13348,n13385,n13386 );
   nand U13264 ( n13386,n12713,n13379 );
   not U13265 ( n13379,p2_reg2_reg_2_ );
   nand U13266 ( n13385,n11159,n13369 );
   not U13267 ( n13369,p2_reg1_reg_2_ );
   and U13268 ( n13345,n13387,n13388 );
   nand U13269 ( n13388,n13373,n13389 );
   nand U13270 ( n13389,n13390,n13391 );
   or U13271 ( n13387,n13391,n13390 );
   nand U13272 ( n13351,p2_addr_reg_2_,n12686 );
   nand U13273 ( n13396,n12687,n13397,n13398 );
   nor U13274 ( n13398,n13399,n13400,n13401,n13402 );
   nor U13275 ( n13402,n13403,n13404 );
   nor U13276 ( n13401,p2_reg1_reg_1_,n13375,n12806 );
   nor U13277 ( n13400,n13405,n13406 );
   nor U13278 ( n13399,p2_reg2_reg_1_,n13384,n12804 );
   nand U13279 ( n13397,n12701,n13407 );
   not U13280 ( n12687,n12800 );
   nand U13281 ( n13394,n13408,n13376 );
   nand U13282 ( n13408,n13409,n13410,n13411 );
   nor U13283 ( n13411,n13412,n13413,n13414 );
   nor U13284 ( n13414,n13403,n13375,n12806 );
   nor U13285 ( n13413,p2_reg1_reg_1_,n13404 );
   nor U13286 ( n13412,n12745,n13407 );
   xor U13287 ( n13407,n13390,n13391 );
   and U13288 ( n13390,n13415,n13416 );
   nand U13289 ( n13416,n12713,n13405 );
   not U13290 ( n13405,p2_reg2_reg_1_ );
   nand U13291 ( n13415,n11159,n13403 );
   not U13292 ( n13403,p2_reg1_reg_1_ );
   or U13293 ( n13410,n13406,p2_reg2_reg_1_ );
   nand U13294 ( n13409,n12690,n13383,p2_reg2_reg_1_ );
   nand U13295 ( n13393,p2_addr_reg_1_,n12686 );
   nand U13296 ( n13392,p2_reg3_reg_1_,p2_u3151 );
   nor U13297 ( n13418,n13419,n13420,n13421 );
   and U13298 ( n13421,n12686,p2_addr_reg_0_ );
   not U13299 ( n12686,n12843 );
   nor U13300 ( n13420,n13422,n11559 );
   nor U13301 ( n13422,n12800,n13423,n13424 );
   nor U13302 ( n13424,p2_reg2_reg_0_,n12804 );
   nor U13303 ( n13423,p2_reg1_reg_0_,n12806 );
   nand U13304 ( n12800,n13425,n13426 );
   or U13305 ( n13426,n11164,n10456 );
   nand U13306 ( n13425,n13427,n11164 );
   nor U13307 ( n13419,p2_state_reg,n11833 );
   not U13308 ( n11833,p2_reg3_reg_0_ );
   nand U13309 ( n13417,n12701,n13428 );
   nand U13310 ( n13428,n13429,n13430,n13391 );
   nand U13311 ( n13391,n13431,n13432,p2_ir_reg_0_ );
   nand U13312 ( n13432,p2_reg1_reg_0_,n11159 );
   nand U13313 ( n13431,n12713,p2_reg2_reg_0_ );
   nand U13314 ( n13430,n13375,n11159 );
   nand U13315 ( n13429,n13384,n12713 );
   nand U13316 ( n13406,n12690,n13384 );
   not U13317 ( n13384,n13383 );
   nand U13318 ( n13383,p2_reg2_reg_0_,n11559 );
   nand U13319 ( n13404,n12716,n13375 );
   not U13320 ( n13375,n13374 );
   nand U13321 ( n13374,p2_reg1_reg_0_,n11559 );
   nand U13322 ( n13427,n13434,n13435 );
   nand U13323 ( n13435,n12843,p2_state_reg,n11166 );
   nand U13324 ( n13434,n13436,n12843,n10650 );
   nand U13325 ( n12843,n13437,n13438,n13439 );
   nand U13326 ( n13438,n12644,n11496 );
   nand U13327 ( n13437,n13433,n11045 );
   nand U13328 ( n13436,n10812,n12667,n13440 );
   nor U13329 ( n13440,n12662,n12507,n11161 );
   not U13330 ( n12662,n12669 );
   not U13331 ( n10812,n10733 );
   nand U13332 ( n10733,n13441,n11049 );
   nand U13333 ( n11049,n11498,n11492,n10662 );
   and U13334 ( n13441,n12153,n12158,n12037 );
   nand U13335 ( n12037,n12508,n11492,n11498 );
   nand U13336 ( n12158,n13442,n11168 );
   nand U13337 ( n12153,n13442,n11498 );
   nor U13338 ( n13446,n13447,n13448,n13449 );
   nor U13339 ( n13449,n10822,n13450 );
   not U13340 ( n10822,n10502 );
   nor U13341 ( n13448,n12188,n13451 );
   and U13342 ( n13447,p2_u3151,p2_reg3_reg_15_ );
   nand U13343 ( n13445,n12189,n13452 );
   nand U13344 ( n13444,n13453,n13454 );
   xor U13345 ( n13454,n13455,n13456 );
   and U13346 ( n13455,n13457,n13458 );
   nand U13347 ( n13443,n13459,n10508 );
   nor U13348 ( n13463,n13464,n13465,n13466 );
   nor U13349 ( n13466,n10746,n13467 );
   nor U13350 ( n13465,n12592,n13451 );
   and U13351 ( n13464,p2_u3151,p2_reg3_reg_26_ );
   nand U13352 ( n13462,n13468,n10469 );
   nand U13353 ( n13461,n13469,n13470,n13453 );
   nand U13354 ( n13470,n13471,n13472 );
   nand U13355 ( n13471,n13473,n13474 );
   nand U13356 ( n13469,n13473,n13474,n13475 );
   not U13357 ( n13475,n13472 );
   nand U13358 ( n13472,n13476,n13477 );
   or U13359 ( n13474,n13478,n13479 );
   nand U13360 ( n13460,n12420,n13480 );
   nor U13361 ( n13484,n13485,n13486,n13487 );
   nor U13362 ( n13487,n11919,n13467 );
   nor U13363 ( n13486,n11961,n13450 );
   and U13364 ( n13485,p2_u3151,p2_reg3_reg_6_ );
   nand U13365 ( n13483,n11962,n13452 );
   nand U13366 ( n13482,n13453,n13488 );
   nand U13367 ( n13488,n13489,n13490,n13491 );
   nand U13368 ( n13491,n10935,n13492 );
   xor U13369 ( n13492,n13493,n13494 );
   nand U13370 ( n13490,n13494,n10532,n13493 );
   nand U13371 ( n13489,n13495,n13496 );
   nand U13372 ( n13481,n13497,n10947 );
   nor U13373 ( n13501,n13502,n13503,n13504 );
   nor U13374 ( n13504,n12236,n13450 );
   nor U13375 ( n13503,n10808,n13467 );
   nor U13376 ( n13502,p2_state_reg,n13505 );
   nand U13377 ( n13500,n13497,n11147 );
   not U13378 ( n11147,n10807 );
   nand U13379 ( n13499,n13453,n13506 );
   xor U13380 ( n13506,n13507,n13508 );
   xor U13381 ( n13507,n13509,n11146 );
   not U13382 ( n11146,n10496 );
   nand U13383 ( n13498,n12243,n13452 );
   nor U13384 ( n13513,n13514,n13515 );
   nor U13385 ( n13515,n11830,n13467 );
   nor U13386 ( n13514,n10971,n13450 );
   nand U13387 ( n13512,n13497,n10995 );
   nand U13388 ( n13511,n13453,n13516 );
   nand U13389 ( n13516,n13517,n13518,n13519 );
   nand U13390 ( n13519,n13520,n13521 );
   xor U13391 ( n13520,n10983,n13522 );
   nand U13392 ( n13518,n13523,n10544,n13524 );
   or U13393 ( n13517,n13525,n13524 );
   nand U13394 ( n13510,p2_reg3_reg_2_,n13526 );
   nor U13395 ( n13530,n12999,n13531,n13532 );
   nor U13396 ( n13532,n10888,n13450 );
   nor U13397 ( n13531,n10887,n13467 );
   not U13398 ( n10887,n10520 );
   nor U13399 ( n12999,p2_state_reg,n13533 );
   not U13400 ( n13533,p2_reg3_reg_11_ );
   nand U13401 ( n13529,n12093,n13452 );
   nand U13402 ( n13528,n13534,n13535,n13453 );
   nand U13403 ( n13535,n13536,n13537 );
   not U13404 ( n13537,n13538 );
   nand U13405 ( n13536,n13539,n13540 );
   nand U13406 ( n13534,n13541,n13538 );
   xor U13407 ( n13541,n13542,n10872 );
   nand U13408 ( n13527,n13497,n11430 );
   not U13409 ( n11430,n10889 );
   nor U13410 ( n13546,n13547,n13548,n13549 );
   nor U13411 ( n13549,n12349,n13467 );
   nor U13412 ( n13548,n12357,n13451 );
   nor U13413 ( n13547,p2_state_reg,n13550 );
   nand U13414 ( n13545,n13468,n10481 );
   nand U13415 ( n13544,n13453,n13551 );
   xor U13416 ( n13551,n13552,n13553 );
   xor U13417 ( n13552,n13554,n10759 );
   not U13418 ( n10759,n10484 );
   nand U13419 ( n13543,n12338,n13480 );
   nor U13420 ( n13558,n13559,n13560,n13561 );
   nor U13421 ( n13561,n12123,n13450 );
   not U13422 ( n12123,n10508 );
   nor U13423 ( n13560,n10888,n13467 );
   and U13424 ( n13559,p2_u3151,p2_reg3_reg_13_ );
   nand U13425 ( n13557,n13497,n10861 );
   nand U13426 ( n13556,n13562,n13563,n13453 );
   nand U13427 ( n13563,n13564,n13565,n13566 );
   nand U13428 ( n13566,n13567,n13568 );
   nand U13429 ( n13564,n13569,n13570 );
   nand U13430 ( n13562,n13571,n13567,n13572 );
   nand U13431 ( n13571,n13573,n13565 );
   nand U13432 ( n13555,n12124,n13452 );
   nor U13433 ( n13577,n13578,n13579,n13580 );
   nor U13434 ( n13580,n12349,n13450 );
   nor U13435 ( n13579,n12236,n13467 );
   nor U13436 ( n13578,p2_state_reg,n13581 );
   nand U13437 ( n13576,n13497,n10790 );
   nand U13438 ( n13575,n13582,n13453 );
   xor U13439 ( n13582,n13583,n13584 );
   xor U13440 ( n13583,n10490,n13585 );
   nand U13441 ( n13574,n12298,n13480 );
   nand U13442 ( n13588,n13453,n11016 );
   nand U13443 ( n11016,n11851,n13590 );
   nand U13444 ( n13590,n11373,n10550 );
   nand U13445 ( n11851,n11006,n11017 );
   nand U13446 ( n13587,n13497,n11017 );
   nand U13447 ( n13586,n13468,n10547 );
   nor U13448 ( n13594,n13595,n13596,n13597 );
   nor U13449 ( n13597,n10914,n13467 );
   nor U13450 ( n13596,n10913,n13451 );
   and U13451 ( n13595,p2_u3151,p2_reg3_reg_9_ );
   nand U13452 ( n13593,n12050,n13452 );
   nand U13453 ( n13592,n13598,n13453 );
   xor U13454 ( n13598,n13599,n13600 );
   xor U13455 ( n13600,n10523,n13601 );
   nand U13456 ( n13591,n13468,n10520 );
   nor U13457 ( n13605,n13273,n13606,n13607 );
   nor U13458 ( n13607,n10971,n13467 );
   nor U13459 ( n13606,n11919,n13450 );
   nor U13460 ( n13273,p2_state_reg,n13608 );
   nand U13461 ( n13604,n11931,n13452 );
   nand U13462 ( n13603,n13453,n13609 );
   xor U13463 ( n13609,n13610,n13611 );
   xor U13464 ( n13610,n13612,n10958 );
   nand U13465 ( n13602,n13497,n11386 );
   nor U13466 ( n13616,n13617,n13618,n13619 );
   nor U13467 ( n13619,n10746,n13450 );
   nor U13468 ( n13618,n10747,n13451 );
   nor U13469 ( n13617,p2_state_reg,n13620 );
   nand U13470 ( n13615,n13459,n10481 );
   nand U13471 ( n13614,n13621,n13453 );
   xor U13472 ( n13621,n13622,n13623 );
   and U13473 ( n13622,n13624,n13625 );
   nand U13474 ( n13613,n12387,n13480 );
   nor U13475 ( n13629,n13630,n13631,n13632 );
   and U13476 ( n13632,n13452,n12227 );
   nor U13477 ( n13631,n10821,n13451 );
   and U13478 ( n13630,p2_u3151,p2_reg3_reg_17_ );
   nand U13479 ( n13628,n13459,n10502 );
   nand U13480 ( n13627,n13633,n13634,n13453 );
   nand U13481 ( n13634,n13635,n13636 );
   nand U13482 ( n13636,n13637,n13638 );
   nand U13483 ( n13633,n13637,n13638,n13639 );
   nand U13484 ( n13626,n13468,n10496 );
   nor U13485 ( n13643,n13644,n13645,n13646 );
   nor U13486 ( n13646,n10958,n13467 );
   not U13487 ( n10958,n10538 );
   nor U13488 ( n13645,n10935,n13450 );
   and U13489 ( n13644,p2_u3151,p2_reg3_reg_5_ );
   nand U13490 ( n13642,n11953,n13452 );
   nand U13491 ( n13641,n13647,n13648,n13453 );
   nand U13492 ( n13648,n13649,n13650 );
   xor U13493 ( n13649,n11919,n13651 );
   nand U13494 ( n13647,n13652,n13653,n13654 );
   nand U13495 ( n13640,n13497,n11404 );
   nor U13496 ( n13658,n12796,n13659,n13660 );
   nor U13497 ( n13660,n10808,n13450 );
   nor U13498 ( n13659,n10834,n13451 );
   nor U13499 ( n12796,p2_state_reg,n13661 );
   nand U13500 ( n13657,n12203,n13452 );
   nand U13501 ( n13656,n13662,n13453 );
   xor U13502 ( n13662,n13663,n13664 );
   xor U13503 ( n13663,n10502,n13665 );
   nand U13504 ( n13655,n13459,n10505 );
   nor U13505 ( n13669,n13670,n13671,n13672 );
   nor U13506 ( n13672,n10728,n13450 );
   nor U13507 ( n13671,n10731,n13451 );
   and U13508 ( n13670,p2_u3151,p2_reg3_reg_25_ );
   nand U13509 ( n13668,n13459,n10478 );
   nand U13510 ( n13667,n13673,n13453 );
   xor U13511 ( n13673,n13674,n13478 );
   nand U13512 ( n13478,n13625,n13675 );
   nand U13513 ( n13675,n13624,n13623 );
   nor U13514 ( n13674,n13479,n13676 );
   not U13515 ( n13479,n13677 );
   nand U13516 ( n13666,n12402,n13480 );
   nor U13517 ( n13681,n13682,n13683,n13684 );
   nor U13518 ( n13684,n13685,n12102 );
   nor U13519 ( n13683,n10874,n13451 );
   nor U13520 ( n13682,p2_state_reg,n13686 );
   nand U13521 ( n13680,n13468,n10511 );
   nand U13522 ( n13679,n13687,n13688,n13453 );
   nand U13523 ( n13688,n13689,n13573 );
   not U13524 ( n13573,n13569 );
   xor U13525 ( n13689,n10888,n13690 );
   nand U13526 ( n13687,n13570,n13565,n13569 );
   nand U13527 ( n13569,n13539,n13691 );
   nand U13528 ( n13691,n13538,n13540 );
   nor U13529 ( n13538,n13692,n13693 );
   not U13530 ( n13539,n13694 );
   nand U13531 ( n13678,n13459,n10517 );
   nor U13532 ( n13698,n13699,n13700,n13701 );
   nor U13533 ( n13701,n10780,n13451 );
   nor U13534 ( n13700,n12591,n13467 );
   not U13535 ( n12591,n10490 );
   and U13536 ( n13699,p2_u3151,p2_reg3_reg_21_ );
   nand U13537 ( n13697,n13468,n10484 );
   nand U13538 ( n13696,n13702,n13703,n13453 );
   nand U13539 ( n13703,n13704,n13705 );
   nand U13540 ( n13705,n13706,n13707 );
   nand U13541 ( n13702,n13706,n13707,n13708 );
   nand U13542 ( n13695,n12309,n13480 );
   nor U13543 ( n13712,n13713,n13714 );
   nor U13544 ( n13714,n11006,n13467 );
   not U13545 ( n11006,n10550 );
   nor U13546 ( n13713,n10983,n13450 );
   nand U13547 ( n13711,n13497,n11379 );
   nand U13548 ( n13710,n13715,n13453 );
   xor U13549 ( n13715,n13716,n13717 );
   and U13550 ( n13716,n13718,n13719 );
   nand U13551 ( n13709,p2_reg3_reg_1_,n13526 );
   nand U13552 ( n13526,n13685,p2_state_reg );
   nor U13553 ( n13723,n13724,n13725,n13726 );
   nor U13554 ( n13726,n11961,n13467 );
   nor U13555 ( n13725,n13685,n12012 );
   not U13556 ( n12012,n13727 );
   and U13557 ( n13724,p2_u3151,p2_reg3_reg_8_ );
   nand U13558 ( n13722,n13497,n10924 );
   not U13559 ( n10924,n12036 );
   nand U13560 ( n13721,n13728,n13453 );
   xor U13561 ( n13728,n13729,n13730 );
   xor U13562 ( n13729,n13731,n10526 );
   nand U13563 ( n13720,n13468,n10523 );
   nor U13564 ( n13735,n13736,n13737,n13738 );
   nor U13565 ( n13738,n12416,n13467 );
   and U13566 ( n13737,n13480,n12497 );
   and U13567 ( n13736,p2_u3151,p2_reg3_reg_28_ );
   nand U13568 ( n13734,n13497,n10697 );
   not U13569 ( n10697,n12496 );
   nand U13570 ( n13733,n13739,n13740,n13453 );
   nand U13571 ( n13740,n13741,n13742 );
   nand U13572 ( n13742,n13743,n13744 );
   nand U13573 ( n13744,n13745,n13746 );
   not U13574 ( n13741,n13747 );
   nand U13575 ( n13739,n13747,n13748 );
   nand U13576 ( n13748,n13746,n13749 );
   nand U13577 ( n13749,n13750,n13743 );
   not U13578 ( n13750,n13745 );
   xor U13579 ( n13747,n12494,n13751 );
   not U13580 ( n12494,n11528 );
   xor U13581 ( n11528,n12532,n12496 );
   nand U13582 ( n12496,n13752,n13753,n12644 );
   nand U13583 ( n13753,n11812,n13754 );
   or U13584 ( n13752,n11788,n11812 );
   not U13585 ( n12532,n10466 );
   nand U13586 ( n13732,n13468,n10463 );
   nand U13587 ( n10463,n13755,n13756,n13757,n12524 );
   nand U13588 ( n12524,n13758,n12661 );
   nand U13589 ( n13757,p2_reg2_reg_29_,n12525 );
   nand U13590 ( n13756,p2_reg1_reg_29_,n12526 );
   nand U13591 ( n13755,p2_reg0_reg_29_,n12527 );
   nor U13592 ( n13762,n12683,n13763,n13764 );
   nor U13593 ( n13764,n12265,n13451 );
   and U13594 ( n13763,n13452,n12266 );
   nor U13595 ( n12683,p2_state_reg,n13765 );
   nand U13596 ( n13761,n13468,n10490 );
   nand U13597 ( n13760,n13453,n13766 );
   xor U13598 ( n13766,n13767,n13768 );
   xor U13599 ( n13768,n13769,n12236 );
   nand U13600 ( n13759,n13459,n10496 );
   nor U13601 ( n13773,n13774,n13312,n13775 );
   nor U13602 ( n13775,p2_reg3_reg_3_,n13685 );
   not U13603 ( n13685,n13452 );
   nor U13604 ( n13312,p2_state_reg,n11910 );
   nor U13605 ( n13774,n10983,n13467 );
   nand U13606 ( n13772,n13468,n10538 );
   nand U13607 ( n13771,n13776,n13777,n13453 );
   nand U13608 ( n13777,n13778,n13779 );
   nand U13609 ( n13779,n13780,n13781 );
   nand U13610 ( n13776,n13782,n13525,n13780,n13781 );
   nand U13611 ( n13782,n13524,n13783 );
   not U13612 ( n13524,n13522 );
   nand U13613 ( n13770,n13497,n11133 );
   nor U13614 ( n13787,n13788,n13789,n13790 );
   nor U13615 ( n13790,n10901,n13467 );
   nor U13616 ( n13789,n10900,n13451 );
   not U13617 ( n10900,n11419 );
   and U13618 ( n13788,p2_u3151,p2_reg3_reg_10_ );
   nand U13619 ( n13786,n12072,n13452 );
   nand U13620 ( n13785,n13453,n13791 );
   nand U13621 ( n13791,n13792,n13793 );
   nand U13622 ( n13793,n13794,n13795 );
   nand U13623 ( n13795,n13796,n13797 );
   nand U13624 ( n13792,n13693,n13796 );
   nor U13625 ( n13693,n13794,n13798 );
   nand U13626 ( n13784,n13468,n10517 );
   nor U13627 ( n13802,n13803,n13804,n13805 );
   nor U13628 ( n13805,n10726,n13450 );
   nor U13629 ( n13804,n10760,n13451 );
   and U13630 ( n13803,p2_u3151,p2_reg3_reg_23_ );
   nand U13631 ( n13801,n13459,n10484 );
   nand U13632 ( n13800,n13453,n13806 );
   xor U13633 ( n13806,n13807,n13808 );
   xor U13634 ( n13808,n10481,n13809 );
   not U13635 ( n13807,n13810 );
   nand U13636 ( n13799,n12366,n13480 );
   nor U13637 ( n13814,n13815,n13816,n13817 );
   nor U13638 ( n13817,n10835,n13450 );
   nor U13639 ( n13816,n12164,n13451 );
   nor U13640 ( n13815,p2_state_reg,n13818 );
   nand U13641 ( n13813,n12145,n13452 );
   nand U13642 ( n13812,n13819,n13453 );
   xor U13643 ( n13819,n13820,n13821 );
   nand U13644 ( n13821,n13822,n13823 );
   nor U13645 ( n13820,n13824,n13825 );
   not U13646 ( n13824,n13826 );
   nand U13647 ( n13811,n13459,n10511 );
   not U13648 ( n13459,n13467 );
   nor U13649 ( n13830,n13831,n13832,n13833 );
   nor U13650 ( n13833,n10728,n13467 );
   nor U13651 ( n13832,n12469,n13451 );
   nor U13652 ( n13831,p2_state_reg,n13834 );
   nand U13653 ( n13829,n13468,n10466 );
   nand U13654 ( n10466,n13835,n13836,n13837,n13838 );
   nand U13655 ( n13838,n13758,n12497 );
   or U13656 ( n12497,n12661,n13839 );
   and U13657 ( n13839,p2_reg3_reg_28_,n13840 );
   nand U13658 ( n13840,n13841,n13834 );
   not U13659 ( n13834,p2_reg3_reg_27_ );
   nor U13660 ( n12661,p2_reg3_reg_27_,p2_reg3_reg_28_,n13842 );
   nand U13661 ( n13837,p2_reg2_reg_28_,n12525 );
   nand U13662 ( n13836,p2_reg1_reg_28_,n12526 );
   nand U13663 ( n13835,p2_reg0_reg_28_,n12527 );
   not U13664 ( n13468,n13450 );
   nand U13665 ( n13828,n13843,n13453 );
   xor U13666 ( n13843,n13844,n13745 );
   nand U13667 ( n13745,n13845,n13476,n13846 );
   nand U13668 ( n13846,n13473,n13624,n13623,n13477 );
   nand U13669 ( n13623,n13847,n13848 );
   nand U13670 ( n13848,n13810,n13849 );
   nand U13671 ( n13849,n10745,n13809 );
   xor U13672 ( n13810,n13850,n10760 );
   nand U13673 ( n10760,n13851,n13852,n12644 );
   nand U13674 ( n13852,n11812,n13853 );
   or U13675 ( n13851,n11744,n11812 );
   or U13676 ( n13847,n13809,n10745 );
   not U13677 ( n10745,n10481 );
   nand U13678 ( n10481,n13854,n13855,n13856,n13857 );
   nand U13679 ( n13857,n13758,n12366 );
   nand U13680 ( n12366,n13858,n13859 );
   nand U13681 ( n13859,p2_reg3_reg_23_,n13860 );
   nand U13682 ( n13860,n13861,n13550 );
   nand U13683 ( n13856,p2_reg2_reg_23_,n12525 );
   nand U13684 ( n13855,p2_reg1_reg_23_,n12526 );
   nand U13685 ( n13854,p2_reg0_reg_23_,n12527 );
   nand U13686 ( n13809,n13862,n13863 );
   nand U13687 ( n13863,n13864,n13554 );
   nand U13688 ( n13554,n13865,n13707 );
   nand U13689 ( n13707,n12349,n13866 );
   xor U13690 ( n13866,n10780,n13751 );
   not U13691 ( n12349,n10487 );
   nand U13692 ( n13865,n13704,n13706 );
   nand U13693 ( n13706,n13867,n10487 );
   nand U13694 ( n10487,n13868,n13869,n13870,n13871 );
   nand U13695 ( n13871,n13758,n12309 );
   nand U13696 ( n12309,n13872,n13873 );
   nand U13697 ( n13873,p2_reg3_reg_21_,n13874 );
   or U13698 ( n13874,n13875,p2_reg3_reg_20_ );
   nand U13699 ( n13870,p2_reg2_reg_21_,n12525 );
   nand U13700 ( n13869,p2_reg1_reg_21_,n12526 );
   nand U13701 ( n13868,p2_reg0_reg_21_,n12527 );
   xor U13702 ( n13867,n13850,n10780 );
   nand U13703 ( n10780,n13876,n13877,n12644 );
   nand U13704 ( n13877,n11812,n13878 );
   or U13705 ( n13876,n11727,n11812 );
   not U13706 ( n13704,n13708 );
   nand U13707 ( n13708,n13879,n13880 );
   nand U13708 ( n13880,n13881,n10490 );
   nand U13709 ( n10490,n13882,n13883,n13884,n13885 );
   nand U13710 ( n13885,n13758,n12298 );
   xor U13711 ( n12298,n13581,n13875 );
   not U13712 ( n13581,p2_reg3_reg_20_ );
   nand U13713 ( n13884,p2_reg2_reg_20_,n12525 );
   nand U13714 ( n13883,p2_reg1_reg_20_,n12526 );
   nand U13715 ( n13882,p2_reg0_reg_20_,n12527 );
   or U13716 ( n13881,n13585,n13584 );
   nand U13717 ( n13879,n13584,n13585 );
   nand U13718 ( n13585,n13886,n13887 );
   nand U13719 ( n13887,n13769,n13888 );
   nand U13720 ( n13888,n12236,n13767 );
   and U13721 ( n13769,n13889,n13890 );
   nand U13722 ( n13890,n13891,n13509 );
   nand U13723 ( n13509,n13892,n13638 );
   nand U13724 ( n13638,n10808,n13893 );
   xor U13725 ( n13893,n10821,n13751 );
   not U13726 ( n10808,n10499 );
   nand U13727 ( n13892,n13635,n13637 );
   nand U13728 ( n13637,n13894,n10499 );
   nand U13729 ( n10499,n13895,n13896,n13897,n13898 );
   nand U13730 ( n13898,n13758,n12227 );
   nand U13731 ( n12227,n13899,n13900 );
   nand U13732 ( n13900,p2_reg3_reg_17_,n13901 );
   nand U13733 ( n13901,n13902,n13661 );
   not U13734 ( n13899,n13903 );
   nand U13735 ( n13897,p2_reg2_reg_17_,n12525 );
   nand U13736 ( n13896,p2_reg1_reg_17_,n12526 );
   nand U13737 ( n13895,p2_reg0_reg_17_,n12527 );
   xor U13738 ( n13894,n13850,n10821 );
   nand U13739 ( n10821,n13904,n13905,n13906 );
   nand U13740 ( n13906,n13907,n12744 );
   nand U13741 ( n12744,n13908,n13909,n11702 );
   nand U13742 ( n13909,n11693,n11810 );
   nand U13743 ( n13908,p2_ir_reg_17_,n11692,p2_ir_reg_31_ );
   nand U13744 ( n13905,n12665,n13910 );
   nand U13745 ( n13904,n12666,n13911 );
   not U13746 ( n13635,n13639 );
   nand U13747 ( n13639,n13912,n13913 );
   nand U13748 ( n13913,n13664,n13914 );
   or U13749 ( n13914,n13665,n10502 );
   xor U13750 ( n13664,n11265,n13751 );
   not U13751 ( n11265,n10834 );
   nand U13752 ( n10834,n13915,n13916,n13917 );
   nand U13753 ( n13917,n13907,n12781 );
   nand U13754 ( n12781,n13918,n13919 );
   or U13755 ( n13919,p2_ir_reg_16_,p2_ir_reg_31_ );
   nand U13756 ( n13918,p2_ir_reg_31_,n11683 );
   nand U13757 ( n11683,n11692,n13920 );
   nand U13758 ( n13920,p2_ir_reg_16_,n13921 );
   not U13759 ( n11692,n11691 );
   nand U13760 ( n13916,n12665,n13922 );
   nand U13761 ( n13915,n12666,n13923 );
   nand U13762 ( n13912,n13665,n10502 );
   nand U13763 ( n10502,n13924,n13925,n13926,n13927 );
   nand U13764 ( n13927,n13758,n12203 );
   xor U13765 ( n12203,n13661,n13928 );
   not U13766 ( n13661,p2_reg3_reg_16_ );
   nand U13767 ( n13926,p2_reg2_reg_16_,n12525 );
   nand U13768 ( n13925,p2_reg1_reg_16_,n12526 );
   nand U13769 ( n13924,p2_reg0_reg_16_,n12527 );
   nand U13770 ( n13665,n13457,n13929 );
   nand U13771 ( n13929,n13456,n13458 );
   nand U13772 ( n13458,n10835,n13930 );
   xor U13773 ( n13930,n13850,n10844 );
   not U13774 ( n10835,n10505 );
   nor U13775 ( n13456,n13931,n13825 );
   nor U13776 ( n13825,n13932,n10508 );
   and U13777 ( n13931,n13826,n13823,n13822 );
   and U13778 ( n13822,n13933,n13567,n13934 );
   nand U13779 ( n13934,n13935,n13568 );
   nand U13780 ( n13935,n13565,n13936 );
   nand U13781 ( n13936,n13694,n13572 );
   nor U13782 ( n13694,n13542,n10872 );
   nand U13783 ( n13565,n13690,n10514 );
   nand U13784 ( n13567,n13937,n10511 );
   xor U13785 ( n13937,n13850,n11116 );
   nand U13786 ( n13933,n13572,n13540,n13798 );
   not U13787 ( n13798,n13797 );
   nand U13788 ( n13797,n13938,n10520 );
   nand U13789 ( n13823,n13572,n13794,n13796,n13540 );
   nand U13790 ( n13540,n10872,n13542 );
   xor U13791 ( n13542,n10889,n13751 );
   nand U13792 ( n10889,n13939,n13940,n13941 );
   nand U13793 ( n13941,n13907,n12990 );
   nand U13794 ( n12990,n13942,n13943,n13944 );
   nand U13795 ( n13943,n11642,n11810 );
   nand U13796 ( n13942,p2_ir_reg_11_,n11641,p2_ir_reg_31_ );
   nand U13797 ( n13940,n12665,n13945 );
   not U13798 ( n13945,n11643 );
   nand U13799 ( n13939,n12666,n13946 );
   not U13800 ( n13946,p1_datao_reg_11_ );
   not U13801 ( n10872,n10517 );
   nand U13802 ( n10517,n13947,n13948,n13949,n13950 );
   nand U13803 ( n13950,n13758,n12093 );
   nand U13804 ( n12093,n13951,n13952 );
   nand U13805 ( n13952,p2_reg3_reg_11_,n13953 );
   nand U13806 ( n13949,p2_reg2_reg_11_,n12525 );
   nand U13807 ( n13948,p2_reg1_reg_11_,n12526 );
   nand U13808 ( n13947,p2_reg0_reg_11_,n12527 );
   not U13809 ( n13796,n13692 );
   nor U13810 ( n13692,n13938,n10520 );
   nand U13811 ( n10520,n13954,n13955,n13956,n13957 );
   nand U13812 ( n13957,n13758,n12072 );
   nand U13813 ( n12072,n13953,n13958 );
   nand U13814 ( n13958,p2_reg3_reg_10_,n13959 );
   nand U13815 ( n13956,p2_reg2_reg_10_,n12525 );
   nand U13816 ( n13955,p2_reg1_reg_10_,n12526 );
   nand U13817 ( n13954,p2_reg0_reg_10_,n12527 );
   xor U13818 ( n13938,n11419,n13751 );
   nand U13819 ( n11419,n13960,n13961,n13962 );
   nand U13820 ( n13962,n13044,n13907 );
   not U13821 ( n13044,n13017 );
   nand U13822 ( n13017,n13963,n13964 );
   or U13823 ( n13964,p2_ir_reg_10_,p2_ir_reg_31_ );
   nand U13824 ( n13963,p2_ir_reg_31_,n11632 );
   nand U13825 ( n11632,n11641,n13965 );
   nand U13826 ( n13965,p2_ir_reg_10_,n13966 );
   not U13827 ( n11641,n11640 );
   nand U13828 ( n13961,n12665,n11633 );
   nand U13829 ( n13960,p1_datao_reg_10_,n12666 );
   and U13830 ( n13794,n13967,n13968 );
   nand U13831 ( n13968,n13601,n13969 );
   or U13832 ( n13969,n13599,n10901 );
   and U13833 ( n13601,n13970,n13971 );
   nand U13834 ( n13971,n13972,n10526 );
   or U13835 ( n13972,n13731,n13730 );
   nand U13836 ( n13970,n13730,n13731 );
   nand U13837 ( n13731,n13973,n13974 );
   nand U13838 ( n13974,n13975,n13976 );
   nand U13839 ( n13976,n13652,n13977 );
   nand U13840 ( n13977,n13654,n13653 );
   not U13841 ( n13654,n13650 );
   nand U13842 ( n13973,n13978,n13979 );
   nand U13843 ( n13978,n13980,n13981 );
   xor U13844 ( n13730,n12036,n13850 );
   nand U13845 ( n12036,n13982,n13983,n13984 );
   nand U13846 ( n13984,n13907,n13096 );
   nand U13847 ( n13096,n13985,n13986 );
   or U13848 ( n13986,p2_ir_reg_31_,p2_ir_reg_8_ );
   nand U13849 ( n13985,p2_ir_reg_31_,n13987 );
   nand U13850 ( n13987,n11616,n11615 );
   nand U13851 ( n11615,p2_ir_reg_8_,n13988 );
   nand U13852 ( n13983,n12665,n13989 );
   not U13853 ( n13989,n11617 );
   nand U13854 ( n13982,n12666,n13990 );
   nand U13855 ( n13967,n10901,n13599 );
   xor U13856 ( n13599,n10913,n13751 );
   nand U13857 ( n10913,n13991,n13992,n13993 );
   nand U13858 ( n13993,n13907,n12983 );
   nand U13859 ( n12983,n13994,n13995,n13966 );
   nand U13860 ( n13995,n11810,n11625 );
   nand U13861 ( n13994,p2_ir_reg_31_,n11616,p2_ir_reg_9_ );
   not U13862 ( n11616,n11624 );
   nand U13863 ( n13992,n12665,n13996 );
   not U13864 ( n13996,n11626 );
   nand U13865 ( n13991,n12666,n13997 );
   not U13866 ( n10901,n10523 );
   nand U13867 ( n10523,n13998,n13999,n14000,n14001 );
   nand U13868 ( n14001,n13758,n12050 );
   nand U13869 ( n12050,n13959,n14002 );
   nand U13870 ( n14002,p2_reg3_reg_9_,n14003 );
   nand U13871 ( n14000,p2_reg2_reg_9_,n12525 );
   nand U13872 ( n13999,p2_reg1_reg_9_,n12526 );
   nand U13873 ( n13998,p2_reg0_reg_9_,n12527 );
   and U13874 ( n13572,n13570,n13568 );
   nand U13875 ( n13568,n14004,n10873 );
   not U13876 ( n10873,n10511 );
   nand U13877 ( n10511,n14005,n14006,n14007,n14008 );
   nand U13878 ( n14008,n13758,n12124 );
   nand U13879 ( n12124,n14009,n14010 );
   nand U13880 ( n14010,p2_reg3_reg_13_,n14011 );
   nand U13881 ( n14011,n14012,n13686 );
   not U13882 ( n13686,p2_reg3_reg_12_ );
   nand U13883 ( n14007,p2_reg2_reg_13_,n12525 );
   nand U13884 ( n14006,p2_reg1_reg_13_,n12526 );
   nand U13885 ( n14005,p2_reg0_reg_13_,n12527 );
   xor U13886 ( n14004,n11116,n13751 );
   not U13887 ( n11116,n10861 );
   nand U13888 ( n10861,n14013,n14014,n14015 );
   nand U13889 ( n14015,n12897,n13907 );
   not U13890 ( n12897,n12910 );
   nand U13891 ( n12910,n14016,n14017,n14018 );
   nand U13892 ( n14017,n11659,n11810 );
   nand U13893 ( n14016,p2_ir_reg_13_,n11658,p2_ir_reg_31_ );
   nand U13894 ( n14014,n12665,n11660 );
   nand U13895 ( n14013,p1_datao_reg_13_,n12666 );
   nand U13896 ( n13570,n10888,n14019 );
   not U13897 ( n14019,n13690 );
   xor U13898 ( n13690,n11425,n13751 );
   not U13899 ( n11425,n10874 );
   nand U13900 ( n10874,n14020,n14021,n14022 );
   nand U13901 ( n14022,n13907,n12938 );
   nand U13902 ( n12938,n14023,n14024 );
   or U13903 ( n14024,p2_ir_reg_12_,p2_ir_reg_31_ );
   nand U13904 ( n14023,p2_ir_reg_31_,n11649 );
   nand U13905 ( n11649,n11658,n14025 );
   nand U13906 ( n14025,p2_ir_reg_12_,n13944 );
   not U13907 ( n11658,n11657 );
   nand U13908 ( n14021,n12665,n14026 );
   not U13909 ( n14026,n11650 );
   nand U13910 ( n14020,n12666,n14027 );
   not U13911 ( n10888,n10514 );
   nand U13912 ( n10514,n14028,n14029,n14030,n14031 );
   nand U13913 ( n14031,n13758,n14032 );
   not U13914 ( n14032,n12102 );
   xor U13915 ( n12102,p2_reg3_reg_12_,n13951 );
   nand U13916 ( n14030,p2_reg2_reg_12_,n12525 );
   nand U13917 ( n14029,p2_reg1_reg_12_,n12526 );
   nand U13918 ( n14028,p2_reg0_reg_12_,n12527 );
   nand U13919 ( n13826,n13932,n10508 );
   nand U13920 ( n10508,n14033,n14034,n14035,n14036 );
   nand U13921 ( n14036,n13758,n12145 );
   xor U13922 ( n12145,n13818,n14009 );
   nand U13923 ( n14035,p2_reg2_reg_14_,n12525 );
   nand U13924 ( n14034,p2_reg1_reg_14_,n12526 );
   nand U13925 ( n14033,p2_reg0_reg_14_,n12527 );
   xor U13926 ( n13932,n12164,n13850 );
   not U13927 ( n12164,n10852 );
   nand U13928 ( n10852,n14037,n14038,n14039 );
   nand U13929 ( n14039,n12862,n13907 );
   not U13930 ( n12862,n12865 );
   nand U13931 ( n12865,n14040,n14041 );
   or U13932 ( n14041,p2_ir_reg_14_,p2_ir_reg_31_ );
   nand U13933 ( n14040,p2_ir_reg_31_,n11666 );
   nand U13934 ( n11666,n11675,n14042 );
   nand U13935 ( n14042,p2_ir_reg_14_,n14018 );
   nand U13936 ( n14038,n12665,n11667 );
   nand U13937 ( n14037,p1_datao_reg_14_,n12666 );
   nand U13938 ( n13457,n14043,n10505 );
   nand U13939 ( n10505,n14044,n14045,n14046,n14047 );
   nand U13940 ( n14047,n13758,n12189 );
   nand U13941 ( n12189,n13928,n14048 );
   nand U13942 ( n14048,p2_reg3_reg_15_,n14049 );
   nand U13943 ( n14049,n14050,n13818 );
   not U13944 ( n13818,p2_reg3_reg_14_ );
   nand U13945 ( n14046,p2_reg2_reg_15_,n12525 );
   nand U13946 ( n14045,p2_reg1_reg_15_,n12526 );
   nand U13947 ( n14044,p2_reg0_reg_15_,n12527 );
   xor U13948 ( n14043,n10844,n13751 );
   not U13949 ( n10844,n12188 );
   nand U13950 ( n12188,n14051,n14052,n14053 );
   nand U13951 ( n14053,n13907,n12816 );
   nand U13952 ( n12816,n14054,n14055,n13921 );
   nand U13953 ( n14055,n11676,n11810 );
   nand U13954 ( n14054,p2_ir_reg_15_,n11675,p2_ir_reg_31_ );
   not U13955 ( n11675,n11674 );
   nand U13956 ( n14052,n12665,n14056 );
   nand U13957 ( n14051,n12666,n14057 );
   not U13958 ( n14057,p1_datao_reg_15_ );
   nand U13959 ( n13891,n13508,n10496 );
   or U13960 ( n13889,n10496,n13508 );
   xor U13961 ( n13508,n13850,n10807 );
   nand U13962 ( n10807,n14058,n14059,n14060 );
   nand U13963 ( n14060,n13907,n12698 );
   nand U13964 ( n12698,n14061,n14062,n14063 );
   nand U13965 ( n14062,n11703,n11810 );
   nand U13966 ( n14061,p2_ir_reg_18_,n11702,p2_ir_reg_31_ );
   nand U13967 ( n14059,n12665,n14064 );
   not U13968 ( n14064,n11704 );
   nand U13969 ( n14058,n12666,n14065 );
   nand U13970 ( n10496,n14066,n14067,n14068,n14069 );
   nand U13971 ( n14069,n13758,n12243 );
   xor U13972 ( n12243,p2_reg3_reg_18_,n13903 );
   nand U13973 ( n14068,p2_reg2_reg_18_,n12525 );
   nand U13974 ( n14067,p2_reg1_reg_18_,n12526 );
   nand U13975 ( n14066,p2_reg0_reg_18_,n12527 );
   or U13976 ( n13886,n13767,n12236 );
   not U13977 ( n12236,n10493 );
   nand U13978 ( n10493,n14070,n14071,n14072,n14073 );
   nand U13979 ( n14073,n13758,n12266 );
   nand U13980 ( n12266,n13875,n14074 );
   nand U13981 ( n14074,p2_reg3_reg_19_,n14075 );
   nand U13982 ( n14075,n13903,n13505 );
   nand U13983 ( n14072,p2_reg2_reg_19_,n12525 );
   nand U13984 ( n14071,p2_reg1_reg_19_,n12526 );
   nand U13985 ( n14070,p2_reg0_reg_19_,n12527 );
   xor U13986 ( n13767,n13751,n12265 );
   nand U13987 ( n12265,n14076,n14077,n14078 );
   nand U13988 ( n14078,n13907,n10662 );
   nand U13989 ( n14077,n12665,n14079 );
   not U13990 ( n14079,n11711 );
   nand U13991 ( n14076,n12666,n14080 );
   xor U13992 ( n13584,n13751,n10790 );
   not U13993 ( n10790,n12297 );
   nand U13994 ( n12297,n14081,n14082,n12644 );
   nand U13995 ( n14082,n11812,n14083 );
   or U13996 ( n14081,n11718,n11812 );
   nand U13997 ( n13864,n13553,n10484 );
   or U13998 ( n13862,n10484,n13553 );
   xor U13999 ( n13553,n13850,n12357 );
   nand U14000 ( n12357,n14084,n14085,n12644 );
   nand U14001 ( n14085,n11812,n14086 );
   or U14002 ( n14084,n11734,n11812 );
   nand U14003 ( n10484,n14087,n14088,n14089,n14090 );
   nand U14004 ( n14090,n13758,n12338 );
   xor U14005 ( n12338,n13550,n13872 );
   not U14006 ( n13550,p2_reg3_reg_22_ );
   nand U14007 ( n14089,p2_reg2_reg_22_,n12525 );
   nand U14008 ( n14088,p2_reg1_reg_22_,n12526 );
   nand U14009 ( n14087,p2_reg0_reg_22_,n12527 );
   nand U14010 ( n13624,n10726,n14091 );
   xor U14011 ( n14091,n10747,n13751 );
   not U14012 ( n10726,n10478 );
   or U14013 ( n13476,n14092,n10728 );
   nand U14014 ( n13845,n14093,n13477,n13473 );
   not U14015 ( n13473,n13676 );
   nand U14016 ( n13676,n14094,n14095 );
   or U14017 ( n14095,n11072,n13850 );
   nand U14018 ( n11072,n11475,n10746 );
   not U14019 ( n11475,n10731 );
   or U14020 ( n14094,n12407,n13751 );
   nand U14021 ( n12407,n10746,n10731 );
   not U14022 ( n10746,n10475 );
   nand U14023 ( n13477,n10728,n14092 );
   xor U14024 ( n14092,n13751,n12592 );
   nand U14025 ( n12592,n14096,n14097,n12644 );
   nand U14026 ( n14097,n11812,n14098 );
   or U14027 ( n14096,n11768,n11812 );
   not U14028 ( n10728,n10472 );
   nand U14029 ( n10472,n14099,n14100,n14101,n14102 );
   nand U14030 ( n14102,n13758,n12420 );
   nand U14031 ( n12420,n13842,n14103 );
   nand U14032 ( n14103,p2_reg3_reg_26_,n14104 );
   not U14033 ( n13842,n13841 );
   nand U14034 ( n14101,p2_reg2_reg_26_,n12525 );
   nand U14035 ( n14100,p2_reg1_reg_26_,n12526 );
   nand U14036 ( n14099,p2_reg0_reg_26_,n12527 );
   nand U14037 ( n14093,n13625,n13677 );
   nand U14038 ( n13677,n14105,n10475 );
   nand U14039 ( n10475,n14106,n14107,n14108,n14109 );
   nand U14040 ( n14109,n13758,n12402 );
   nand U14041 ( n12402,n14104,n14110 );
   nand U14042 ( n14110,p2_reg3_reg_25_,n14111 );
   nand U14043 ( n14111,n14112,n13620 );
   nand U14044 ( n14108,p2_reg2_reg_25_,n12525 );
   nand U14045 ( n14107,p2_reg1_reg_25_,n12526 );
   nand U14046 ( n14106,p2_reg0_reg_25_,n12527 );
   xor U14047 ( n14105,n13850,n10731 );
   nand U14048 ( n10731,n14113,n14114,n12644 );
   nand U14049 ( n14114,n11812,n14115 );
   or U14050 ( n14113,n11761,n11812 );
   nand U14051 ( n13625,n14116,n10478 );
   nand U14052 ( n10478,n14117,n14118,n14119,n14120 );
   nand U14053 ( n14120,n13758,n12387 );
   xor U14054 ( n12387,n13620,n13858 );
   not U14055 ( n13620,p2_reg3_reg_24_ );
   nand U14056 ( n14119,p2_reg2_reg_24_,n12525 );
   nand U14057 ( n14118,p2_reg1_reg_24_,n12526 );
   nand U14058 ( n14117,p2_reg0_reg_24_,n12527 );
   xor U14059 ( n14116,n13850,n10747 );
   nand U14060 ( n10747,n14121,n14122,n12644 );
   nand U14061 ( n14122,n11812,n14123 );
   or U14062 ( n14121,n11751,n11812 );
   and U14063 ( n13844,n13746,n13743 );
   nand U14064 ( n13743,n14124,n10469 );
   xor U14065 ( n14124,n13850,n12469 );
   nand U14066 ( n13746,n12416,n14125 );
   xor U14067 ( n14125,n12469,n13751 );
   nand U14068 ( n12469,n14126,n14127,n12644 );
   nand U14069 ( n14127,n11812,n14128 );
   or U14070 ( n14126,n11778,n11812 );
   not U14071 ( n12416,n10469 );
   nand U14072 ( n10469,n14129,n14130,n14131,n14132 );
   nand U14073 ( n14132,n13758,n12470 );
   nand U14074 ( n14131,p2_reg2_reg_27_,n12525 );
   nand U14075 ( n14130,p2_reg1_reg_27_,n12526 );
   nand U14076 ( n14129,p2_reg0_reg_27_,n12527 );
   nand U14077 ( n13827,n12470,n13480 );
   nand U14078 ( n13480,n14133,n14134,n14135 );
   nand U14079 ( n14135,n14136,p2_state_reg );
   xor U14080 ( n12470,p2_reg3_reg_27_,n13841 );
   nor U14081 ( n13841,n14104,p2_reg3_reg_26_ );
   or U14082 ( n14104,p2_reg3_reg_24_,p2_reg3_reg_25_,n13858 );
   not U14083 ( n13858,n14112 );
   nor U14084 ( n14112,p2_reg3_reg_22_,p2_reg3_reg_23_,n13872 );
   not U14085 ( n13872,n13861 );
   nor U14086 ( n13861,p2_reg3_reg_20_,p2_reg3_reg_21_,n13875 );
   nand U14087 ( n13875,n13505,n13765,n13903 );
   nor U14088 ( n13903,p2_reg3_reg_16_,p2_reg3_reg_17_,n13928 );
   not U14089 ( n13928,n13902 );
   nor U14090 ( n13902,p2_reg3_reg_14_,p2_reg3_reg_15_,n14009 );
   not U14091 ( n14009,n14050 );
   nor U14092 ( n14050,p2_reg3_reg_12_,p2_reg3_reg_13_,n13951 );
   not U14093 ( n13951,n14012 );
   nor U14094 ( n14012,n13953,p2_reg3_reg_11_ );
   or U14095 ( n13953,n13959,p2_reg3_reg_10_ );
   or U14096 ( n13959,n14003,p2_reg3_reg_9_ );
   not U14097 ( n13765,p2_reg3_reg_19_ );
   not U14098 ( n13505,p2_reg3_reg_18_ );
   nor U14099 ( n14140,n14141,n14142,n14143 );
   nor U14100 ( n14143,n10935,n13467 );
   nor U14101 ( n14142,n10914,n13450 );
   not U14102 ( n12500,n12646 );
   nor U14103 ( n12659,n11164,n11159 );
   not U14104 ( n10914,n10526 );
   nand U14105 ( n10526,n14144,n14145,n14146,n14147 );
   nand U14106 ( n14147,n13758,n13727 );
   nand U14107 ( n13727,n14003,n14148 );
   nand U14108 ( n14148,p2_reg3_reg_8_,n14149 );
   or U14109 ( n14003,n14149,p2_reg3_reg_8_ );
   nand U14110 ( n14146,p2_reg2_reg_8_,n12525 );
   nand U14111 ( n14145,p2_reg1_reg_8_,n12526 );
   nand U14112 ( n14144,p2_reg0_reg_8_,n12527 );
   and U14113 ( n14141,p2_u3151,p2_reg3_reg_7_ );
   nand U14114 ( n14139,n11990,n13452 );
   nand U14115 ( n13452,n14133,n14134,n14150 );
   nand U14116 ( n14150,n14136,n10650 );
   nor U14117 ( n14136,n12667,n11025 );
   nand U14118 ( n14134,n14151,p2_state_reg );
   nand U14119 ( n14151,n14152,n14153,n14154,n14155 );
   and U14120 ( n14155,n11045,n11160,n11493 );
   nand U14121 ( n11493,n12499,n12508 );
   nand U14122 ( n14154,n12499,n11498 );
   not U14123 ( n12499,n11496 );
   nand U14124 ( n14153,n11024,n14156 );
   nand U14125 ( n14152,n14157,n14158 );
   nand U14126 ( n14133,n11031,n14156 );
   and U14127 ( n11031,n12507,n11161,n10650 );
   not U14128 ( n12507,n11163 );
   nand U14129 ( n14138,n14159,n14160,n13453 );
   nand U14130 ( n14161,n14162,n14163 );
   nand U14131 ( n14163,n11026,n11024 );
   nor U14132 ( n11024,n10659,n11168 );
   not U14133 ( n11026,n14156 );
   nand U14134 ( n14156,n10655,n10665,n10649 );
   nand U14135 ( n14162,n11025,n14157 );
   nand U14136 ( n14157,n14164,n12678,n11368,n11978 );
   nand U14137 ( n11978,n10663,n11161 );
   not U14138 ( n10663,n10661 );
   nand U14139 ( n10661,n11168,n11030 );
   nand U14140 ( n11368,n10660,n11492 );
   nand U14141 ( n12678,n14165,n11030 );
   not U14142 ( n14165,n11979 );
   nand U14143 ( n11979,n11161,n11498 );
   nor U14144 ( n11161,n10660,n12508 );
   or U14145 ( n14164,n10659,n11498 );
   nand U14146 ( n10659,n13442,n11030 );
   nor U14147 ( n13442,n10660,n10662 );
   not U14148 ( n11025,n14158 );
   nand U14149 ( n14160,n14166,n13981,n14167 );
   nand U14150 ( n14167,n13980,n13979 );
   nand U14151 ( n14166,n13496,n14168 );
   not U14152 ( n13496,n13493 );
   nand U14153 ( n14159,n14169,n13980,n13975 );
   and U14154 ( n13975,n13979,n14168 );
   nand U14155 ( n14168,n13494,n10935 );
   nand U14156 ( n13979,n11961,n14170 );
   xor U14157 ( n14170,n13850,n11413 );
   not U14158 ( n11961,n10529 );
   nand U14159 ( n13980,n14171,n10529 );
   nand U14160 ( n10529,n14172,n14173,n14174,n14175 );
   nand U14161 ( n14175,n13758,n11990 );
   nand U14162 ( n11990,n14149,n14176 );
   nand U14163 ( n14176,p2_reg3_reg_7_,n14177 );
   or U14164 ( n14149,n14177,p2_reg3_reg_7_ );
   nand U14165 ( n14174,p2_reg2_reg_7_,n12525 );
   nand U14166 ( n14173,p2_reg1_reg_7_,n12526 );
   nand U14167 ( n14172,p2_reg0_reg_7_,n12527 );
   xor U14168 ( n14171,n11413,n13751 );
   nand U14169 ( n14169,n13493,n13981 );
   not U14170 ( n13981,n13495 );
   nor U14171 ( n13495,n13494,n10935 );
   not U14172 ( n10935,n10532 );
   nand U14173 ( n10532,n14178,n14179,n14180,n14181 );
   nand U14174 ( n14181,p2_reg2_reg_6_,n12525 );
   nand U14175 ( n14180,p2_reg1_reg_6_,n12526 );
   nand U14176 ( n14179,p2_reg0_reg_6_,n12527 );
   nand U14177 ( n14178,n13758,n11962 );
   nand U14178 ( n11962,n14177,n14182 );
   nand U14179 ( n14182,p2_reg3_reg_6_,n14183 );
   or U14180 ( n14177,n14183,p2_reg3_reg_6_ );
   xor U14181 ( n13494,n10947,n13850 );
   nand U14182 ( n10947,n14184,n14185,n14186 );
   nand U14183 ( n14186,n13218,n13907 );
   not U14184 ( n13218,n13179 );
   nand U14185 ( n13179,n14187,n14188 );
   or U14186 ( n14188,p2_ir_reg_31_,p2_ir_reg_6_ );
   nand U14187 ( n14187,p2_ir_reg_31_,n14189 );
   nand U14188 ( n14189,n11600,n11599 );
   nand U14189 ( n11599,p2_ir_reg_6_,n14190 );
   nand U14190 ( n14185,n12665,n11601 );
   nand U14191 ( n14184,p1_datao_reg_6_,n12666 );
   nand U14192 ( n13493,n13653,n14191 );
   nand U14193 ( n14191,n13652,n13650 );
   nand U14194 ( n13650,n14192,n14193 );
   nand U14195 ( n14193,n14194,n13612 );
   nand U14196 ( n13612,n14195,n13781 );
   nand U14197 ( n13781,n14196,n10971 );
   not U14198 ( n10971,n10541 );
   xor U14199 ( n14196,n10984,n13751 );
   nand U14200 ( n14195,n13778,n13780 );
   nand U14201 ( n13780,n14197,n10541 );
   nand U14202 ( n10541,n14198,n14199,n14200,n14201 );
   nand U14203 ( n14201,p2_reg2_reg_3_,n12525 );
   nand U14204 ( n14200,p2_reg1_reg_3_,n12526 );
   nand U14205 ( n14199,p2_reg0_reg_3_,n12527 );
   nand U14206 ( n14198,n13758,n11910 );
   xor U14207 ( n14197,n13850,n10984 );
   not U14208 ( n10984,n11133 );
   nand U14209 ( n11133,n14202,n14203,n14204 );
   nand U14210 ( n14204,n13320,n13907 );
   not U14211 ( n13320,n13294 );
   nand U14212 ( n13294,n14205,n14206,n14207 );
   nand U14213 ( n14206,n11810,n11577 );
   nand U14214 ( n14205,p2_ir_reg_31_,n11576,p2_ir_reg_3_ );
   nand U14215 ( n14203,n12665,n11578 );
   nand U14216 ( n14202,p1_datao_reg_3_,n12666 );
   and U14217 ( n13778,n13783,n14208 );
   nand U14218 ( n14208,n13525,n13522 );
   nand U14219 ( n13522,n13718,n14209 );
   nand U14220 ( n14209,n13717,n13719 );
   nand U14221 ( n13719,n14210,n11830 );
   not U14222 ( n11830,n10547 );
   xor U14223 ( n14210,n11005,n13751 );
   nand U14224 ( n13717,n11841,n14211 );
   nand U14225 ( n14211,n11373,n13751 );
   not U14226 ( n11373,n11017 );
   nand U14227 ( n11841,n11017,n10550 );
   nand U14228 ( n10550,n14212,n14213,n14214,n14215 );
   nand U14229 ( n14215,p2_reg2_reg_0_,n12525 );
   nand U14230 ( n14214,p2_reg1_reg_0_,n12526 );
   nand U14231 ( n14213,p2_reg0_reg_0_,n12527 );
   nand U14232 ( n14212,p2_reg3_reg_0_,n13758 );
   nand U14233 ( n11017,n14216,n14217,n14218 );
   nand U14234 ( n14218,p2_ir_reg_0_,n13907 );
   nand U14235 ( n14217,n11551,n12665 );
   nand U14236 ( n14216,n12666,p1_datao_reg_0_ );
   nand U14237 ( n13718,n14219,n10547 );
   nand U14238 ( n10547,n14220,n14221,n14222,n14223 );
   nand U14239 ( n14223,p2_reg2_reg_1_,n12525 );
   nand U14240 ( n14222,p2_reg1_reg_1_,n12526 );
   nand U14241 ( n14221,p2_reg0_reg_1_,n12527 );
   nand U14242 ( n14220,p2_reg3_reg_1_,n13758 );
   xor U14243 ( n14219,n13850,n11005 );
   not U14244 ( n11005,n11379 );
   nand U14245 ( n11379,n14224,n14225,n14226 );
   nand U14246 ( n14226,n13373,n13907 );
   not U14247 ( n13373,n13376 );
   nand U14248 ( n13376,n14227,n14228,n14229 );
   nand U14249 ( n14228,n11560,n11810 );
   nand U14250 ( n14227,p2_ir_reg_1_,p2_ir_reg_0_,p2_ir_reg_31_ );
   nand U14251 ( n14225,n11561,n12665 );
   nand U14252 ( n14224,p1_datao_reg_1_,n12666 );
   nand U14253 ( n13525,n10983,n13523 );
   not U14254 ( n13523,n13521 );
   not U14255 ( n10983,n10544 );
   nand U14256 ( n13783,n13521,n10544 );
   nand U14257 ( n10544,n14230,n14231,n14232,n14233 );
   nand U14258 ( n14233,p2_reg2_reg_2_,n12525 );
   nand U14259 ( n14232,p2_reg1_reg_2_,n12526 );
   nand U14260 ( n14231,p2_reg0_reg_2_,n12527 );
   nand U14261 ( n14230,p2_reg3_reg_2_,n13758 );
   xor U14262 ( n13521,n10995,n13751 );
   not U14263 ( n10995,n12588 );
   nand U14264 ( n12588,n14234,n14235,n14236 );
   nand U14265 ( n14236,n13907,n13331 );
   nand U14266 ( n13331,n14237,n14238 );
   or U14267 ( n14238,p2_ir_reg_2_,p2_ir_reg_31_ );
   nand U14268 ( n14237,p2_ir_reg_31_,n11567 );
   nand U14269 ( n11567,n11576,n14239 );
   nand U14270 ( n14239,p2_ir_reg_2_,n14229 );
   not U14271 ( n11576,n11575 );
   nand U14272 ( n14235,n14240,n12665 );
   not U14273 ( n14240,n11568 );
   nand U14274 ( n14234,n12666,n14241 );
   not U14275 ( n14241,p1_datao_reg_2_ );
   nand U14276 ( n14194,n13611,n10538 );
   or U14277 ( n14192,n10538,n13611 );
   xor U14278 ( n13611,n11386,n13751 );
   not U14279 ( n11386,n10970 );
   nand U14280 ( n10970,n14242,n14243,n14244 );
   nand U14281 ( n14244,n13907,n13258 );
   nand U14282 ( n13258,n14245,n14246 );
   or U14283 ( n14246,p2_ir_reg_31_,p2_ir_reg_4_ );
   nand U14284 ( n14245,p2_ir_reg_31_,n14247 );
   nand U14285 ( n14247,n11584,n11583 );
   nand U14286 ( n11583,p2_ir_reg_4_,n14207 );
   nand U14287 ( n14243,n12665,n14248 );
   not U14288 ( n14248,n11585 );
   nand U14289 ( n14242,n12666,n14249 );
   not U14290 ( n14249,p1_datao_reg_4_ );
   nand U14291 ( n10538,n14250,n14251,n14252,n14253 );
   nand U14292 ( n14253,n11931,n13758 );
   xor U14293 ( n11931,p2_reg3_reg_3_,n13608 );
   nand U14294 ( n14252,p2_reg2_reg_4_,n12525 );
   nand U14295 ( n14251,p2_reg1_reg_4_,n12526 );
   nand U14296 ( n14250,p2_reg0_reg_4_,n12527 );
   nand U14297 ( n13652,n13651,n10535 );
   nand U14298 ( n13653,n11919,n14254 );
   not U14299 ( n14254,n13651 );
   xor U14300 ( n13651,n11404,n13751 );
   nand U14301 ( n14255,n11498,n11030,n10653 );
   nand U14302 ( n11163,n11168,n11492 );
   nand U14303 ( n12594,n11168,n10662 );
   not U14304 ( n10662,n12508 );
   not U14305 ( n11404,n10957 );
   nand U14306 ( n10957,n14256,n14257,n14258 );
   nand U14307 ( n14258,n13907,n13226 );
   nand U14308 ( n13226,n14259,n14260,n14190 );
   nand U14309 ( n14260,n11810,n11593 );
   nand U14310 ( n14259,p2_ir_reg_31_,n11584,p2_ir_reg_5_ );
   not U14311 ( n11584,n11592 );
   nand U14312 ( n14257,n12665,n14261 );
   not U14313 ( n14261,n11594 );
   nand U14314 ( n14256,n12666,n14262 );
   not U14315 ( n11919,n10535 );
   nand U14316 ( n10535,n14263,n14264,n14265,n14266 );
   nand U14317 ( n14266,n13758,n11953 );
   nand U14318 ( n11953,n14183,n14267 );
   nand U14319 ( n14267,p2_reg3_reg_5_,n14268 );
   or U14320 ( n14183,n14268,p2_reg3_reg_5_ );
   nand U14321 ( n14268,n13608,n11910 );
   not U14322 ( n11910,p2_reg3_reg_3_ );
   not U14323 ( n13608,p2_reg3_reg_4_ );
   nand U14324 ( n14265,p2_reg2_reg_5_,n12525 );
   nand U14325 ( n14264,p2_reg1_reg_5_,n12526 );
   not U14326 ( n14271,n14269 );
   nand U14327 ( n14263,p2_reg0_reg_5_,n12527 );
   nand U14328 ( n14269,n14272,n14273 );
   nand U14329 ( n14273,p2_ir_reg_29_,n11810 );
   nand U14330 ( n14272,p2_ir_reg_31_,n11793 );
   nand U14331 ( n11793,p2_ir_reg_29_,n11809 );
   xor U14332 ( n14270,n11810,n11803 );
   not U14333 ( n11803,p2_ir_reg_30_ );
   nand U14334 ( n14137,n13497,n11413 );
   not U14335 ( n11413,n10936 );
   nand U14336 ( n10936,n14274,n14275,n14276 );
   nand U14337 ( n14276,n13907,n13149 );
   nand U14338 ( n13149,n14277,n14278,n13988 );
   nand U14339 ( n14278,n11810,n11609 );
   nand U14340 ( n14277,p2_ir_reg_31_,n11600,p2_ir_reg_7_ );
   not U14341 ( n11600,n11608 );
   nand U14342 ( n14275,n12665,n14279 );
   not U14343 ( n14279,n11610 );
   nand U14344 ( n14274,n12666,n14280 );
   not U14345 ( n14280,p1_datao_reg_7_ );
   not U14346 ( n13497,n13451 );
   nand U14347 ( n14281,n12669,n14282 );
   or U14348 ( n14282,n12667,n14158 );
   nand U14349 ( n14158,n10653,n10666,n10649 );
   and U14350 ( n10649,n14283,n14284,n14285,n14286 );
   nor U14351 ( n14286,n14287,n14288,n14289,n14290 );
   not U14352 ( n11814,p2_d_reg_6_ );
   not U14353 ( n11816,p2_d_reg_13_ );
   not U14354 ( n11818,p2_d_reg_17_ );
   nor U14355 ( n14291,p2_d_reg_22_,p2_d_reg_24_,p2_d_reg_23_ );
   nor U14356 ( n14285,n14292,n14293,n14294,n14295 );
   not U14357 ( n11820,p2_d_reg_19_ );
   not U14358 ( n11817,p2_d_reg_16_ );
   nor U14359 ( n14296,p2_d_reg_7_,p2_d_reg_9_,p2_d_reg_8_ );
   not U14360 ( n11815,p2_d_reg_10_ );
   nor U14361 ( n14284,n14297,n14298,n14299,n14300 );
   not U14362 ( n11822,p2_d_reg_29_ );
   not U14363 ( n11813,p2_d_reg_2_ );
   not U14364 ( n11821,p2_d_reg_27_ );
   not U14365 ( n11819,p2_d_reg_18_ );
   nor U14366 ( n14283,n14301,n14302,n14303,n14304 );
   nor U14367 ( n14305,p2_d_reg_5_,p2_d_reg_4_,p2_d_reg_3_,p2_d_reg_30_ );
   nor U14368 ( n14306,p2_d_reg_20_,p2_d_reg_26_,p2_d_reg_25_ );
   nor U14369 ( n14307,p2_d_reg_15_,p2_d_reg_14_,p2_d_reg_12_,p2_d_reg_11_ );
   nor U14370 ( n14308,p2_d_reg_21_,p2_d_reg_31_,p2_d_reg_28_ );
   not U14371 ( n10666,n10655 );
   nand U14372 ( n10655,n11036,n14309 );
   nand U14373 ( n11036,n14310,n14311 );
   not U14374 ( n10653,n10665 );
   nand U14375 ( n10665,n11039,n14312 );
   and U14376 ( n14313,n14314,n14311 );
   xor U14377 ( n14314,n14315,n12660 );
   not U14378 ( n12660,p2_b_reg );
   nand U14379 ( n11039,n14315,n14310 );
   nand U14380 ( n12667,n10675,n14316 );
   nand U14381 ( n14316,n11168,n12508 );
   not U14382 ( n10675,n10730 );
   nand U14383 ( n12669,n10686,n11030 );
   not U14384 ( n10686,n10714 );
   nand U14385 ( n10714,n12508,n10660,n11168 );
   not U14386 ( n11168,n11498 );
   nand U14387 ( n11498,n14317,n14318 );
   nand U14388 ( n14318,p2_ir_reg_20_,n11810 );
   nand U14389 ( n14317,n11716,n11717,p2_ir_reg_31_ );
   nand U14390 ( n11716,p2_ir_reg_20_,n11710 );
   nand U14391 ( n12508,n14319,n14320 );
   nand U14392 ( n14320,p2_ir_reg_19_,n11810 );
   nand U14393 ( n14319,n11709,n11710,p2_ir_reg_31_ );
   nand U14394 ( n11709,p2_ir_reg_19_,n14063 );
   nor U14395 ( n10650,n13433,p2_u3151,n11166 );
   nand U14396 ( n14321,n11496,n11160,n12644 );
   not U14397 ( n11160,n13433 );
   nor U14398 ( n13433,n14310,n14315,n14311 );
   nand U14399 ( n14311,n14322,n14323,n14324 );
   nand U14400 ( n14323,n11760,n11810 );
   nand U14401 ( n14322,p2_ir_reg_25_,n11759,p2_ir_reg_31_ );
   nand U14402 ( n14315,n14325,n14326 );
   or U14403 ( n14326,p2_ir_reg_24_,p2_ir_reg_31_ );
   nand U14404 ( n14325,p2_ir_reg_31_,n11750 );
   nand U14405 ( n11750,n11759,n14327 );
   nand U14406 ( n14327,p2_ir_reg_24_,n14328 );
   not U14407 ( n11759,n11758 );
   nand U14408 ( n14310,n14329,n14330 );
   or U14409 ( n14330,p2_ir_reg_26_,p2_ir_reg_31_ );
   nand U14410 ( n14329,p2_ir_reg_31_,n11767 );
   nand U14411 ( n11767,n11776,n14331 );
   nand U14412 ( n14331,p2_ir_reg_26_,n14324 );
   nand U14413 ( n11496,n11165,n11492 );
   not U14414 ( n11492,n11030 );
   nand U14415 ( n11030,n14332,n14333,n14334 );
   nand U14416 ( n14333,n11726,n11810 );
   nand U14417 ( n14332,p2_ir_reg_21_,n11717,p2_ir_reg_31_ );
   not U14418 ( n11717,n11725 );
   not U14419 ( n11165,n10660 );
   nand U14420 ( n10660,n14335,n14336 );
   or U14421 ( n14336,p2_ir_reg_22_,p2_ir_reg_31_ );
   nand U14422 ( n14335,p2_ir_reg_31_,n11733 );
   nand U14423 ( n11733,n11742,n14337 );
   nand U14424 ( n14337,p2_ir_reg_22_,n14334 );
   and U14425 ( n13439,n14338,p2_state_reg );
   nand U14426 ( n14338,n11166,n12644 );
   nand U14427 ( n12644,n11159,n11164 );
   nand U14428 ( n11164,n14339,n14340,n11809 );
   nand U14429 ( n11809,n11785,n11787 );
   not U14430 ( n11785,n11786 );
   nand U14431 ( n14340,n11787,n11810 );
   not U14432 ( n11787,p2_ir_reg_28_ );
   nand U14433 ( n14339,p2_ir_reg_28_,n11786,p2_ir_reg_31_ );
   nand U14434 ( n11786,n11775,n11777 );
   nand U14435 ( n14342,n11777,n11810 );
   not U14436 ( n11777,p2_ir_reg_27_ );
   nand U14437 ( n14341,p2_ir_reg_27_,n11776,p2_ir_reg_31_ );
   not U14438 ( n11776,n11775 );
   nor U14439 ( n11775,n14324,p2_ir_reg_26_ );
   nand U14440 ( n14324,n11758,n11760 );
   not U14441 ( n11760,p2_ir_reg_25_ );
   nor U14442 ( n11758,n14328,p2_ir_reg_24_ );
   not U14443 ( n11166,n11045 );
   nand U14444 ( n11045,n14343,n14344,n14328 );
   nand U14445 ( n14328,n11741,n11743 );
   nand U14446 ( n14344,n11743,n11810 );
   not U14447 ( n11810,p2_ir_reg_31_ );
   not U14448 ( n11743,p2_ir_reg_23_ );
   nand U14449 ( n14343,p2_ir_reg_23_,n11742,p2_ir_reg_31_ );
   not U14450 ( n11742,n11741 );
   nor U14451 ( n11741,n14334,p2_ir_reg_22_ );
   nand U14452 ( n14334,n11725,n11726 );
   not U14453 ( n11726,p2_ir_reg_21_ );
   nor U14454 ( n11725,n11710,p2_ir_reg_20_ );
   or U14455 ( n11710,n14063,p2_ir_reg_19_ );
   nand U14456 ( n14063,n11701,n11703 );
   not U14457 ( n11703,p2_ir_reg_18_ );
   not U14458 ( n11701,n11702 );
   nand U14459 ( n11702,n11691,n11693 );
   not U14460 ( n11693,p2_ir_reg_17_ );
   nor U14461 ( n11691,n13921,p2_ir_reg_16_ );
   nand U14462 ( n13921,n11674,n11676 );
   not U14463 ( n11676,p2_ir_reg_15_ );
   nor U14464 ( n11674,n14018,p2_ir_reg_14_ );
   nand U14465 ( n14018,n11657,n11659 );
   not U14466 ( n11659,p2_ir_reg_13_ );
   nor U14467 ( n11657,n13944,p2_ir_reg_12_ );
   nand U14468 ( n13944,n11640,n11642 );
   not U14469 ( n11642,p2_ir_reg_11_ );
   nor U14470 ( n11640,n13966,p2_ir_reg_10_ );
   nand U14471 ( n13966,n11624,n11625 );
   not U14472 ( n11625,p2_ir_reg_9_ );
   nor U14473 ( n11624,n13988,p2_ir_reg_8_ );
   nand U14474 ( n13988,n11608,n11609 );
   not U14475 ( n11609,p2_ir_reg_7_ );
   nor U14476 ( n11608,n14190,p2_ir_reg_6_ );
   nand U14477 ( n14190,n11592,n11593 );
   not U14478 ( n11593,p2_ir_reg_5_ );
   nor U14479 ( n11592,n14207,p2_ir_reg_4_ );
   nand U14480 ( n14207,n11575,n11577 );
   not U14481 ( n11577,p2_ir_reg_3_ );
   nor U14482 ( n11575,n14229,p2_ir_reg_2_ );
   nand U14483 ( n14229,n11559,n11560 );
   not U14484 ( n11560,p2_ir_reg_1_ );
   not U14485 ( n11559,p2_ir_reg_0_ );
   nand U14486 ( n14346,p1_datao_reg_31_,n14347 );
   nand U14487 ( n14345,p1_u3973,n14348 );
   nand U14488 ( n14350,p1_datao_reg_30_,n14347 );
   nand U14489 ( n14349,p1_u3973,n14351 );
   nand U14490 ( n14353,p1_datao_reg_29_,n14347 );
   nand U14491 ( n14352,p1_u3973,n14354 );
   nand U14492 ( n14356,p1_datao_reg_28_,n14347 );
   nand U14493 ( n14355,p1_u3973,n14357 );
   nand U14494 ( n14359,p1_datao_reg_27_,n14347 );
   nand U14495 ( n14358,p1_u3973,n14360 );
   nand U14496 ( n14362,p1_datao_reg_26_,n14347 );
   nand U14497 ( n14361,p1_u3973,n14363 );
   nand U14498 ( n14365,p1_datao_reg_25_,n14347 );
   nand U14499 ( n14364,p1_u3973,n14366 );
   nand U14500 ( n14368,p1_datao_reg_24_,n14347 );
   nand U14501 ( n14367,p1_u3973,n14369 );
   nand U14502 ( n14371,p1_datao_reg_23_,n14347 );
   nand U14503 ( n14370,p1_u3973,n14372 );
   nand U14504 ( n14374,p1_datao_reg_22_,n14347 );
   nand U14505 ( n14373,p1_u3973,n14375 );
   nand U14506 ( n14377,p1_datao_reg_21_,n14347 );
   nand U14507 ( n14376,p1_u3973,n14378 );
   nand U14508 ( n14380,p1_datao_reg_20_,n14347 );
   nand U14509 ( n14379,p1_u3973,n14381 );
   nand U14510 ( n14383,p1_datao_reg_19_,n14347 );
   nand U14511 ( n14382,p1_u3973,n14384 );
   nand U14512 ( n14386,p1_datao_reg_18_,n14347 );
   nand U14513 ( n14385,p1_u3973,n14387 );
   nand U14514 ( n14389,p1_datao_reg_17_,n14347 );
   nand U14515 ( n14388,p1_u3973,n14390 );
   nand U14516 ( n14392,p1_datao_reg_16_,n14347 );
   nand U14517 ( n14391,p1_u3973,n14393 );
   nand U14518 ( n14395,p1_datao_reg_15_,n14347 );
   nand U14519 ( n14394,p1_u3973,n14396 );
   nand U14520 ( n14398,p1_datao_reg_14_,n14347 );
   nand U14521 ( n14397,p1_u3973,n14399 );
   nand U14522 ( n14401,p1_datao_reg_13_,n14347 );
   nand U14523 ( n14400,p1_u3973,n14402 );
   nand U14524 ( n14404,p1_datao_reg_12_,n14347 );
   nand U14525 ( n14403,p1_u3973,n14405 );
   nand U14526 ( n14407,p1_datao_reg_11_,n14347 );
   nand U14527 ( n14406,p1_u3973,n14408 );
   nand U14528 ( n14410,p1_datao_reg_10_,n14347 );
   nand U14529 ( n14409,p1_u3973,n14411 );
   nand U14530 ( n14413,p1_datao_reg_9_,n14347 );
   nand U14531 ( n14412,p1_u3973,n14414 );
   nand U14532 ( n14416,p1_datao_reg_8_,n14347 );
   nand U14533 ( n14415,p1_u3973,n14417 );
   nand U14534 ( n14419,p1_datao_reg_7_,n14347 );
   nand U14535 ( n14418,p1_u3973,n14420 );
   nand U14536 ( n14422,p1_datao_reg_6_,n14347 );
   nand U14537 ( n14421,p1_u3973,n14423 );
   nand U14538 ( n14425,p1_datao_reg_5_,n14347 );
   nand U14539 ( n14424,p1_u3973,n14426 );
   nand U14540 ( n14428,p1_datao_reg_4_,n14347 );
   nand U14541 ( n14427,p1_u3973,n14429 );
   nand U14542 ( n14431,p1_datao_reg_3_,n14347 );
   nand U14543 ( n14430,p1_u3973,n14432 );
   nand U14544 ( n14434,p1_datao_reg_2_,n14347 );
   nand U14545 ( n14433,p1_u3973,n14435 );
   nand U14546 ( n14437,p1_datao_reg_1_,n14347 );
   nand U14547 ( n14436,p1_u3973,n14438 );
   nand U14548 ( n14440,p1_datao_reg_0_,n14347 );
   nand U14549 ( n14439,p1_u3973,n14441 );
   nand U14550 ( n14442,p1_reg1_reg_31_,n14446 );
   nand U14551 ( n14448,p1_reg1_reg_30_,n14446 );
   nand U14552 ( n14447,n14444,n14449 );
   nand U14553 ( n14451,p1_reg1_reg_29_,n14446 );
   nand U14554 ( n14450,n14444,n14452 );
   nand U14555 ( n14454,p1_reg1_reg_28_,n14446 );
   nand U14556 ( n14453,n14444,n14455 );
   nand U14557 ( n14457,p1_reg1_reg_27_,n14446 );
   nand U14558 ( n14456,n14444,n14458 );
   nand U14559 ( n14460,p1_reg1_reg_26_,n14446 );
   nand U14560 ( n14459,n14444,n14461 );
   nand U14561 ( n14463,p1_reg1_reg_25_,n14446 );
   nand U14562 ( n14462,n14444,n14464 );
   nand U14563 ( n14466,p1_reg1_reg_24_,n14446 );
   nand U14564 ( n14465,n14444,n14467 );
   nand U14565 ( n14469,p1_reg1_reg_23_,n14446 );
   nand U14566 ( n14468,n14444,n14470 );
   nand U14567 ( n14472,p1_reg1_reg_22_,n14446 );
   nand U14568 ( n14471,n14444,n14473 );
   nand U14569 ( n14475,p1_reg1_reg_21_,n14446 );
   nand U14570 ( n14474,n14444,n14476 );
   nand U14571 ( n14478,p1_reg1_reg_20_,n14446 );
   nand U14572 ( n14477,n14444,n14479 );
   nand U14573 ( n14481,p1_reg1_reg_19_,n14446 );
   nand U14574 ( n14480,n14444,n14482 );
   nand U14575 ( n14484,p1_reg1_reg_18_,n14446 );
   nand U14576 ( n14483,n14444,n14485 );
   nand U14577 ( n14487,p1_reg1_reg_17_,n14446 );
   nand U14578 ( n14486,n14444,n14488 );
   nand U14579 ( n14490,p1_reg1_reg_16_,n14446 );
   nand U14580 ( n14489,n14444,n14491 );
   nand U14581 ( n14493,p1_reg1_reg_15_,n14446 );
   nand U14582 ( n14492,n14444,n14494 );
   nand U14583 ( n14496,p1_reg1_reg_14_,n14446 );
   nand U14584 ( n14495,n14444,n14497 );
   nand U14585 ( n14499,p1_reg1_reg_13_,n14446 );
   nand U14586 ( n14498,n14444,n14500 );
   nand U14587 ( n14502,p1_reg1_reg_12_,n14446 );
   nand U14588 ( n14501,n14444,n14503 );
   nand U14589 ( n14505,p1_reg1_reg_11_,n14446 );
   nand U14590 ( n14504,n14444,n14506 );
   nand U14591 ( n14508,p1_reg1_reg_10_,n14446 );
   nand U14592 ( n14507,n14444,n14509 );
   nand U14593 ( n14511,p1_reg1_reg_9_,n14446 );
   nand U14594 ( n14510,n14444,n14512 );
   nand U14595 ( n14514,p1_reg1_reg_8_,n14446 );
   nand U14596 ( n14513,n14444,n14515 );
   nand U14597 ( n14517,p1_reg1_reg_7_,n14446 );
   nand U14598 ( n14516,n14444,n14518 );
   nand U14599 ( n14520,p1_reg1_reg_6_,n14446 );
   nand U14600 ( n14519,n14444,n14521 );
   nand U14601 ( n14523,p1_reg1_reg_5_,n14446 );
   nand U14602 ( n14522,n14444,n14524 );
   nand U14603 ( n14526,p1_reg1_reg_4_,n14446 );
   nand U14604 ( n14525,n14444,n14527 );
   nand U14605 ( n14529,p1_reg1_reg_3_,n14446 );
   nand U14606 ( n14528,n14444,n14530 );
   nand U14607 ( n14532,p1_reg1_reg_2_,n14446 );
   nand U14608 ( n14531,n14444,n14533 );
   nand U14609 ( n14535,p1_reg1_reg_1_,n14446 );
   nand U14610 ( n14534,n14444,n14536 );
   nand U14611 ( n14538,p1_reg1_reg_0_,n14446 );
   nand U14612 ( n14537,n14444,n14539 );
   nand U14613 ( n14445,n14546,n14547,n14548 );
   nand U14614 ( n14548,n14549,n14550 );
   nand U14615 ( n14546,n14551,n14552 );
   nand U14616 ( n14543,p1_reg0_reg_31_,n14553 );
   nand U14617 ( n14449,n14556,n14547,n14557 );
   nand U14618 ( n14557,n14558,n14550 );
   not U14619 ( n14547,n14559 );
   nand U14620 ( n14556,n14560,n14561,n14551 );
   nand U14621 ( n14554,p1_reg0_reg_30_,n14553 );
   nand U14622 ( n14452,n14564,n14565,n14566,n14567 );
   or U14623 ( n14567,n14568,n14569 );
   nand U14624 ( n14566,n14551,n14570 );
   nand U14625 ( n14565,n14571,n14550 );
   not U14626 ( n14564,n14572 );
   nand U14627 ( n14562,p1_reg0_reg_29_,n14553 );
   nand U14628 ( n14455,n14575,n14576,n14577,n14578 );
   nand U14629 ( n14578,n14579,n14354 );
   nor U14630 ( n14577,n14580,n14581 );
   nor U14631 ( n14581,n14568,n14582 );
   and U14632 ( n14580,n14551,n14583 );
   nand U14633 ( n14576,n14584,n14550 );
   nand U14634 ( n14573,p1_reg0_reg_28_,n14553 );
   nand U14635 ( n14458,n14587,n14588,n14589 );
   nor U14636 ( n14589,n14590,n14591,n14592 );
   nor U14637 ( n14592,n14568,n14593 );
   and U14638 ( n14591,n14594,n14551 );
   nor U14639 ( n14590,n14595,n14596 );
   nand U14640 ( n14588,n14597,n14550 );
   nand U14641 ( n14585,p1_reg0_reg_27_,n14553 );
   nand U14642 ( n14461,n14600,n14601,n14602 );
   nor U14643 ( n14602,n14603,n14604,n14605 );
   nor U14644 ( n14605,n14568,n14606 );
   nor U14645 ( n14604,n14607,n14608 );
   nor U14646 ( n14603,n14609,n14596 );
   nand U14647 ( n14601,n14610,n14550 );
   nand U14648 ( n14598,p1_reg0_reg_26_,n14553 );
   nand U14649 ( n14464,n14613,n14614,n14615,n14616 );
   nor U14650 ( n14616,n14617,n14618,n14619 );
   nor U14651 ( n14619,n14620,n14596 );
   nor U14652 ( n14618,n14621,n14622 );
   nor U14653 ( n14617,n14623,n14624 );
   nand U14654 ( n14615,n14625,n14626 );
   not U14655 ( n14625,n14627 );
   nand U14656 ( n14614,n14551,n14628 );
   nand U14657 ( n14613,n14629,n14630 );
   nand U14658 ( n14611,p1_reg0_reg_25_,n14553 );
   nand U14659 ( n14467,n14633,n14634,n14635,n14636 );
   nor U14660 ( n14636,n14637,n14638,n14639 );
   nor U14661 ( n14639,n14640,n14596 );
   nor U14662 ( n14638,n14641,n14622 );
   nor U14663 ( n14637,n14623,n14642 );
   nand U14664 ( n14635,n14643,n14551 );
   nand U14665 ( n14634,n14644,n14630 );
   nand U14666 ( n14633,n14645,n14626 );
   not U14667 ( n14645,n14646 );
   nand U14668 ( n14631,p1_reg0_reg_24_,n14553 );
   nand U14669 ( n14470,n14649,n14650,n14651,n14652 );
   nand U14670 ( n14652,n14579,n14369 );
   nor U14671 ( n14651,n14653,n14654 );
   nor U14672 ( n14654,n14655,n14568 );
   and U14673 ( n14653,n14656,n14551 );
   nand U14674 ( n14650,n14657,n14550 );
   nand U14675 ( n14647,p1_reg0_reg_23_,n14553 );
   nand U14676 ( n14473,n14660,n14661,n14662,n14663 );
   nor U14677 ( n14663,n14664,n14665,n14666 );
   nor U14678 ( n14666,n14641,n14596 );
   nor U14679 ( n14665,n14667,n14622 );
   nor U14680 ( n14664,n14623,n14668 );
   or U14681 ( n14662,n14669,n14607 );
   nand U14682 ( n14660,n14670,n14630 );
   nand U14683 ( n14658,p1_reg0_reg_22_,n14553 );
   nand U14684 ( n14476,n14673,n14674,n14675,n14676 );
   nor U14685 ( n14676,n14677,n14678 );
   nor U14686 ( n14677,n14623,n14679 );
   nand U14687 ( n14675,n14579,n14375 );
   nand U14688 ( n14674,n14551,n14680 );
   nand U14689 ( n14673,n14681,n14682 );
   nand U14690 ( n14671,p1_reg0_reg_21_,n14553 );
   nand U14691 ( n14479,n14685,n14686,n14687 );
   nor U14692 ( n14687,n14688,n14689,n14690 );
   nor U14693 ( n14690,n14568,n14691 );
   nor U14694 ( n14689,n14607,n14692 );
   nor U14695 ( n14688,n14667,n14596 );
   nand U14696 ( n14686,n14693,n14550 );
   nand U14697 ( n14683,p1_reg0_reg_20_,n14553 );
   nand U14698 ( n14482,n14696,n14697,n14698,n14699 );
   nor U14699 ( n14699,n14700,n14701,n14702 );
   nor U14700 ( n14702,n14703,n14596 );
   nor U14701 ( n14701,n14704,n14622 );
   nor U14702 ( n14700,n14623,n14705 );
   nand U14703 ( n14698,n14706,n14626 );
   nand U14704 ( n14697,n14551,n14707 );
   nand U14705 ( n14696,n14708,n14630 );
   nand U14706 ( n14694,p1_reg0_reg_19_,n14553 );
   nand U14707 ( n14485,n14711,n14712,n14713,n14714 );
   nor U14708 ( n14714,n14715,n14716,n14717 );
   nor U14709 ( n14717,n14718,n14596 );
   nor U14710 ( n14716,n14719,n14622 );
   nor U14711 ( n14715,n14623,n14720 );
   nand U14712 ( n14713,n14721,n14551 );
   nand U14713 ( n14712,n14722,n14630 );
   nand U14714 ( n14711,n14723,n14626 );
   nand U14715 ( n14709,p1_reg0_reg_18_,n14553 );
   nand U14716 ( n14488,n14726,n14727,n14728 );
   nor U14717 ( n14728,n14729,n14730,n14731 );
   nor U14718 ( n14731,n14568,n14732 );
   and U14719 ( n14730,n14733,n14551 );
   nor U14720 ( n14729,n14704,n14596 );
   nand U14721 ( n14727,n14734,n14550 );
   nand U14722 ( n14724,p1_reg0_reg_17_,n14553 );
   nand U14723 ( n14491,n14737,n14738,n14739,n14740 );
   nand U14724 ( n14740,n14579,n14390 );
   nor U14725 ( n14739,n14741,n14742 );
   nor U14726 ( n14742,n14743,n14568 );
   nor U14727 ( n14741,n14607,n14744 );
   nand U14728 ( n14738,n14745,n14550 );
   nand U14729 ( n14735,p1_reg0_reg_16_,n14553 );
   nand U14730 ( n14494,n14748,n14749,n14750,n14751 );
   nor U14731 ( n14751,n14752,n14753,n14754 );
   nor U14732 ( n14754,n14755,n14596 );
   nor U14733 ( n14753,n14756,n14622 );
   nor U14734 ( n14752,n14623,n14757 );
   nand U14735 ( n14750,n14758,n14630 );
   nand U14736 ( n14748,n14551,n14759 );
   nand U14737 ( n14746,p1_reg0_reg_15_,n14553 );
   nand U14738 ( n14497,n14762,n14763,n14764,n14765 );
   nor U14739 ( n14765,n14766,n14767,n14768 );
   nor U14740 ( n14768,n14623,n14769 );
   nor U14741 ( n14767,n14770,n14596 );
   nand U14742 ( n14764,n14771,n14402 );
   nand U14743 ( n14763,n14772,n14630 );
   or U14744 ( n14762,n14773,n14607 );
   nand U14745 ( n14760,p1_reg0_reg_14_,n14553 );
   nand U14746 ( n14500,n14776,n14777,n14778 );
   nor U14747 ( n14778,n14779,n14780,n14781 );
   nor U14748 ( n14781,n14568,n14782 );
   and U14749 ( n14780,n14783,n14551 );
   nor U14750 ( n14779,n14756,n14596 );
   nand U14751 ( n14777,n14784,n14550 );
   nand U14752 ( n14774,p1_reg0_reg_13_,n14553 );
   nand U14753 ( n14503,n14787,n14788,n14789,n14790 );
   nor U14754 ( n14790,n14791,n14792,n14793 );
   nor U14755 ( n14793,n14794,n14596 );
   nor U14756 ( n14792,n14795,n14622 );
   nor U14757 ( n14791,n14623,n14796 );
   or U14758 ( n14789,n14797,n14607 );
   nand U14759 ( n14788,n14798,n14630 );
   nand U14760 ( n14787,n14799,n14626 );
   not U14761 ( n14799,n14800 );
   nand U14762 ( n14785,p1_reg0_reg_12_,n14553 );
   nand U14763 ( n14506,n14803,n14804,n14805 );
   nor U14764 ( n14805,n14806,n14807,n14808 );
   nor U14765 ( n14808,n14568,n14809 );
   and U14766 ( n14807,n14810,n14551 );
   nor U14767 ( n14806,n14811,n14596 );
   nand U14768 ( n14804,n14812,n14550 );
   nand U14769 ( n14801,p1_reg0_reg_11_,n14553 );
   nand U14770 ( n14509,n14815,n14816,n14817 );
   nor U14771 ( n14817,n14818,n14819,n14820 );
   nor U14772 ( n14820,n14568,n14821 );
   nor U14773 ( n14819,n14607,n14822 );
   nor U14774 ( n14818,n14795,n14596 );
   nand U14775 ( n14816,n14823,n14550 );
   nand U14776 ( n14813,p1_reg0_reg_10_,n14553 );
   nand U14777 ( n14512,n14826,n14827,n14828,n14829 );
   nor U14778 ( n14829,n14830,n14831,n14832 );
   nor U14779 ( n14832,n14833,n14596 );
   nor U14780 ( n14831,n14834,n14622 );
   nor U14781 ( n14830,n14623,n14835 );
   nand U14782 ( n14828,n14836,n14626 );
   nand U14783 ( n14827,n14551,n14837 );
   nand U14784 ( n14826,n14838,n14630 );
   nand U14785 ( n14824,p1_reg0_reg_9_,n14553 );
   nand U14786 ( n14515,n14841,n14842,n14843 );
   nor U14787 ( n14843,n14844,n14845,n14846 );
   nor U14788 ( n14846,n14568,n14847 );
   nor U14789 ( n14845,n14607,n14848 );
   nor U14790 ( n14844,n14849,n14596 );
   nand U14791 ( n14842,n14850,n14550 );
   nand U14792 ( n14839,p1_reg0_reg_8_,n14553 );
   nand U14793 ( n14518,n14853,n14854,n14855 );
   nor U14794 ( n14855,n14856,n14857,n14858 );
   nor U14795 ( n14858,n14568,n14859 );
   and U14796 ( n14857,n14860,n14551 );
   nor U14797 ( n14856,n14834,n14596 );
   nand U14798 ( n14854,n14861,n14550 );
   nand U14799 ( n14851,p1_reg0_reg_7_,n14553 );
   nand U14800 ( n14521,n14864,n14865,n14866 );
   nor U14801 ( n14866,n14867,n14868,n14869 );
   nor U14802 ( n14869,n14568,n14870 );
   nor U14803 ( n14868,n14607,n14871 );
   nor U14804 ( n14867,n14872,n14596 );
   nand U14805 ( n14865,n14873,n14550 );
   nand U14806 ( n14862,p1_reg0_reg_6_,n14553 );
   nand U14807 ( n14524,n14876,n14877,n14878,n14879 );
   nor U14808 ( n14879,n14880,n14881,n14882 );
   nor U14809 ( n14882,n14883,n14596 );
   nor U14810 ( n14881,n14884,n14622 );
   nor U14811 ( n14880,n14623,n14885 );
   nand U14812 ( n14878,n14886,n14626 );
   not U14813 ( n14886,n14887 );
   nand U14814 ( n14877,n14551,n14888 );
   nand U14815 ( n14876,n14889,n14630 );
   nand U14816 ( n14874,p1_reg0_reg_5_,n14553 );
   nand U14817 ( n14527,n14892,n14893,n14894,n14895 );
   nor U14818 ( n14895,n14896,n14897,n14898 );
   nor U14819 ( n14898,n14899,n14596 );
   nor U14820 ( n14897,n14900,n14622 );
   nor U14821 ( n14896,n14623,n14901 );
   or U14822 ( n14894,n14902,n14607 );
   nand U14823 ( n14893,n14903,n14630 );
   not U14824 ( n14903,n14904 );
   nand U14825 ( n14892,n14905,n14626 );
   nand U14826 ( n14890,p1_reg0_reg_4_,n14553 );
   nand U14827 ( n14530,n14908,n14909,n14910,n14911 );
   nor U14828 ( n14911,n14912,n14913,n14914 );
   nor U14829 ( n14914,n14623,n14915 );
   nor U14830 ( n14913,n14884,n14596 );
   nand U14831 ( n14910,n14771,n14435 );
   nand U14832 ( n14909,n14551,n14916 );
   nand U14833 ( n14908,n14917,n14630 );
   nand U14834 ( n14906,p1_reg0_reg_3_,n14553 );
   nand U14835 ( n14533,n14920,n14921,n14922,n14923 );
   nor U14836 ( n14923,n14924,n14925,n14926 );
   nor U14837 ( n14926,n14900,n14596 );
   nor U14838 ( n14925,n14927,n14622 );
   nor U14839 ( n14924,n14623,n14928 );
   or U14840 ( n14922,n14929,n14607 );
   nand U14841 ( n14920,n14930,n14630 );
   not U14842 ( n14930,n14931 );
   nand U14843 ( n14918,p1_reg0_reg_2_,n14553 );
   nand U14844 ( n14536,n14934,n14935,n14936,n14937 );
   nor U14845 ( n14937,n14938,n14939,n14940 );
   nor U14846 ( n14940,n14941,n14596 );
   nor U14847 ( n14939,n14942,n14622 );
   nor U14848 ( n14938,n14623,n14943 );
   nand U14849 ( n14936,n14944,n14626 );
   not U14850 ( n14944,n14945 );
   nand U14851 ( n14935,n14551,n14946 );
   nand U14852 ( n14934,n14947,n14630 );
   nand U14853 ( n14630,n14948,n14568 );
   nand U14854 ( n14932,p1_reg0_reg_1_,n14553 );
   nand U14855 ( n14539,n14951,n14952,n14953,n14954 );
   nand U14856 ( n14954,n14955,n14956 );
   nand U14857 ( n14955,n14623,n14607 );
   nand U14858 ( n14953,n14579,n14438 );
   nand U14859 ( n14952,n14957,n14682 );
   not U14860 ( n14951,n14958 );
   nand U14861 ( n14949,p1_reg0_reg_0_,n14553 );
   and U14862 ( n14542,n14960,n14961,n14962 );
   nand U14863 ( n14960,n14963,n14964,n14965 );
   nand U14864 ( n14964,n14966,n14967 );
   nand U14865 ( n14963,n14968,n14969 );
   nand U14866 ( n14969,n14967,n14970 );
   nand U14867 ( n14971,n14974,n14975 );
   nand U14868 ( n14976,n14974,n14978 );
   nor U14869 ( n14982,n14983,n14984,n14985 );
   nor U14870 ( n14985,n14569,n14986 );
   xor U14871 ( n14569,n14987,n14988 );
   and U14872 ( n14984,n14989,n14990 );
   and U14873 ( n14983,n14570,n14991 );
   xor U14874 ( n14570,n14992,n14993 );
   nand U14875 ( n14981,n14994,n14571 );
   nand U14876 ( n14980,p1_reg2_reg_29_,n14995 );
   nand U14877 ( n14572,n14997,n14998,n14999,n15000 );
   nor U14878 ( n15000,n15001,n15002 );
   nor U14879 ( n15002,n14595,n14622 );
   nor U14880 ( n15001,n15003,n15004 );
   nand U14881 ( n14999,n15005,n15006 );
   nand U14882 ( n15006,n15007,n15008,n15009 );
   or U14883 ( n15009,n15010,n14987 );
   nand U14884 ( n15008,n15010,n14987,n15011 );
   or U14885 ( n15007,n15011,n14987 );
   nand U14886 ( n15005,n15012,n15013 );
   nand U14887 ( n14998,n15014,n15015 );
   xor U14888 ( n15015,n15016,n14987 );
   nand U14889 ( n15016,n15011,n15010 );
   nand U14890 ( n15010,n15017,n15018 );
   nand U14891 ( n14997,n15019,n15020 );
   xor U14892 ( n15019,n15021,n14988 );
   nand U14893 ( n14988,n15022,n15023 );
   nand U14894 ( n15023,n14595,n15024 );
   nand U14895 ( n15024,n14584,n15025 );
   or U14896 ( n15022,n15025,n14584 );
   nand U14897 ( n15028,n15029,n11551 );
   nand U14898 ( n15027,p1_ir_reg_0_,n15030 );
   nand U14899 ( n15026,n15033,p2_datao_reg_0_ );
   nand U14900 ( n15037,n15032,n15038 );
   nand U14901 ( n15036,n15033,p2_datao_reg_1_ );
   nand U14902 ( n15035,n15031,p1_ir_reg_1_ );
   nand U14903 ( n15034,n15029,n11561 );
   nand U14904 ( n15042,n15043,n15044,n15032 );
   nand U14905 ( n15041,n15033,p2_datao_reg_2_ );
   nand U14906 ( n15040,n15031,p1_ir_reg_2_ );
   nand U14907 ( n15039,n15029,n11568 );
   nand U14908 ( n15048,n15049,n15032 );
   nand U14909 ( n15047,n15033,p2_datao_reg_3_ );
   nand U14910 ( n15046,n15031,p1_ir_reg_3_ );
   nand U14911 ( n15045,n15029,n11578 );
   nand U14912 ( n15053,n15054,n15055,n15032 );
   nand U14913 ( n15052,n15033,p2_datao_reg_4_ );
   nand U14914 ( n15051,n15031,p1_ir_reg_4_ );
   nand U14915 ( n15050,n15029,n11585 );
   nand U14916 ( n15059,p1_ir_reg_5_,n15060 );
   nand U14917 ( n15060,n15061,n15062 );
   nand U14918 ( n15062,n15032,n15063 );
   nand U14919 ( n15058,n15032,n15055,n15064 );
   nand U14920 ( n15057,n15033,p2_datao_reg_5_ );
   nand U14921 ( n15056,n15029,n11594 );
   nand U14922 ( n15068,n15069,n15070,n15032 );
   nand U14923 ( n15067,n15033,p2_datao_reg_6_ );
   nand U14924 ( n15066,n15031,p1_ir_reg_6_ );
   nand U14925 ( n15065,n15029,n11601 );
   nand U14926 ( n15074,p1_ir_reg_7_,n15075 );
   nand U14927 ( n15075,n15061,n15076 );
   nand U14928 ( n15076,n15032,n15077 );
   nand U14929 ( n15073,n15032,n15070,n15078 );
   nand U14930 ( n15072,n15033,p2_datao_reg_7_ );
   nand U14931 ( n15071,n15029,n11610 );
   nand U14932 ( n15082,n15083,n15084,n15032 );
   nand U14933 ( n15081,n15033,p2_datao_reg_8_ );
   nand U14934 ( n15080,n15031,p1_ir_reg_8_ );
   nand U14935 ( n15079,n15029,n11617 );
   nand U14936 ( n15088,n15089,n15032 );
   nand U14937 ( n15087,n15033,p2_datao_reg_9_ );
   nand U14938 ( n15086,n15031,p1_ir_reg_9_ );
   nand U14939 ( n15085,n15029,n11626 );
   nand U14940 ( n15093,n15094,n15032 );
   not U14941 ( n15094,n15095 );
   nand U14942 ( n15092,n15033,p2_datao_reg_10_ );
   nand U14943 ( n15091,n15031,p1_ir_reg_10_ );
   nand U14944 ( n15090,n15029,n11633 );
   nand U14945 ( n15099,n15100,n15032 );
   nand U14946 ( n15098,n15033,p2_datao_reg_11_ );
   nand U14947 ( n15097,n15031,p1_ir_reg_11_ );
   nand U14948 ( n15096,n15029,n11643 );
   nand U14949 ( n15104,n15105,n15106,n15032 );
   nand U14950 ( n15103,n15033,p2_datao_reg_12_ );
   nand U14951 ( n15102,n15031,p1_ir_reg_12_ );
   nand U14952 ( n15101,n15029,n11650 );
   nand U14953 ( n15110,p1_ir_reg_13_,n15111 );
   nand U14954 ( n15111,n15061,n15112 );
   nand U14955 ( n15112,n15032,n15113 );
   nand U14956 ( n15109,n15032,n15106,n15114 );
   nand U14957 ( n15108,n15033,p2_datao_reg_13_ );
   nand U14958 ( n15107,n15029,n11660 );
   nand U14959 ( n15118,n15119,n15032 );
   not U14960 ( n15119,n15120 );
   nand U14961 ( n15117,n15033,p2_datao_reg_14_ );
   nand U14962 ( n15116,n15031,p1_ir_reg_14_ );
   nand U14963 ( n15115,n15029,n11667 );
   nand U14964 ( n15124,p1_ir_reg_15_,n15125 );
   nand U14965 ( n15125,n15061,n15126 );
   nand U14966 ( n15126,n15032,n15127 );
   nand U14967 ( n15123,n15032,n15128,n15129 );
   nand U14968 ( n15122,n15033,p2_datao_reg_15_ );
   nand U14969 ( n15121,n15029,n11677 );
   nand U14970 ( n15133,n15134,n15135,n15032 );
   nand U14971 ( n15132,n15033,p2_datao_reg_16_ );
   nand U14972 ( n15131,n15031,p1_ir_reg_16_ );
   nand U14973 ( n15130,n15029,n11684 );
   nand U14974 ( n15139,p1_ir_reg_17_,n15140 );
   nand U14975 ( n15140,n15061,n15141 );
   nand U14976 ( n15141,n15032,n15142 );
   nand U14977 ( n15138,n15032,n15135,n15143 );
   nand U14978 ( n15137,n15033,p2_datao_reg_17_ );
   nand U14979 ( n15136,n15029,n11694 );
   nand U14980 ( n15147,p1_ir_reg_18_,n15148 );
   nand U14981 ( n15148,n15061,n15149 );
   nand U14982 ( n15149,n15032,n15150 );
   nand U14983 ( n15146,n15032,n15151,n15152 );
   nand U14984 ( n15145,n15033,p2_datao_reg_18_ );
   nand U14985 ( n15144,n15029,n11704 );
   nand U14986 ( n15156,n15157,n15158,n15032 );
   nand U14987 ( n15155,n15033,p2_datao_reg_19_ );
   nand U14988 ( n15154,n15031,p1_ir_reg_19_ );
   nand U14989 ( n15153,n15029,n11711 );
   nand U14990 ( n15162,n15163,n15164,n15032 );
   nand U14991 ( n15161,n15033,p2_datao_reg_20_ );
   nand U14992 ( n15160,n15031,p1_ir_reg_20_ );
   nand U14993 ( n15159,n15029,n11718 );
   nand U14994 ( n15168,p1_ir_reg_21_,n15169 );
   nand U14995 ( n15169,n15061,n15170 );
   nand U14996 ( n15170,n15032,n15171 );
   nand U14997 ( n15167,n15032,n15164,n15172 );
   nand U14998 ( n15166,n15033,p2_datao_reg_21_ );
   nand U14999 ( n15165,n15029,n11727 );
   nand U15000 ( n15176,n15177,n15178,n15032 );
   nand U15001 ( n15175,n15033,p2_datao_reg_22_ );
   nand U15002 ( n15174,n15031,p1_ir_reg_22_ );
   nand U15003 ( n15173,n15029,n11734 );
   nand U15004 ( n15182,p1_ir_reg_23_,n15183 );
   nand U15005 ( n15183,n15061,n15184 );
   nand U15006 ( n15184,n15032,n15185 );
   nand U15007 ( n15181,n15032,n15178,n15186 );
   nand U15008 ( n15180,n15033,p2_datao_reg_23_ );
   nand U15009 ( n15179,n15029,n11744 );
   nand U15010 ( n15190,n15191,n15192,n15032 );
   nand U15011 ( n15189,n15033,p2_datao_reg_24_ );
   nand U15012 ( n15188,n15031,p1_ir_reg_24_ );
   nand U15013 ( n15187,n15029,n11751 );
   nand U15014 ( n15196,p1_ir_reg_25_,n15197 );
   nand U15015 ( n15197,n15061,n15198 );
   nand U15016 ( n15198,n15032,n15199 );
   nand U15017 ( n15195,n15032,n15192,n15200 );
   nand U15018 ( n15194,n15033,p2_datao_reg_25_ );
   nand U15019 ( n15193,n15029,n11761 );
   nand U15020 ( n15204,n15205,n15206,n15032 );
   nand U15021 ( n15203,n15033,p2_datao_reg_26_ );
   nand U15022 ( n15202,n15031,p1_ir_reg_26_ );
   nand U15023 ( n15201,n15029,n11768 );
   nand U15024 ( n15210,p1_ir_reg_27_,n15211 );
   nand U15025 ( n15211,n15061,n15212 );
   nand U15026 ( n15212,n15032,n15213 );
   nand U15027 ( n15209,n15032,n15206,n15214 );
   nand U15028 ( n15208,n15033,p2_datao_reg_27_ );
   nand U15029 ( n15207,n15029,n11778 );
   nand U15030 ( n15218,n15219,n15220,n15032 );
   nand U15031 ( n15217,n15033,p2_datao_reg_28_ );
   nand U15032 ( n15216,n15031,p1_ir_reg_28_ );
   nand U15033 ( n15215,n15029,n11788 );
   nand U15034 ( n15224,p1_ir_reg_29_,n15225 );
   nand U15035 ( n15225,n15061,n15226 );
   nand U15036 ( n15226,n15227,n15032 );
   nand U15037 ( n15223,n15032,n15220,n15228 );
   nand U15038 ( n15222,n15033,p2_datao_reg_29_ );
   nand U15039 ( n15221,n15029,n11795 );
   nand U15040 ( n15232,p1_ir_reg_30_,n15233 );
   nand U15041 ( n15233,n15061,n15234 );
   nand U15042 ( n15234,n15235,n15032 );
   nand U15043 ( n15231,n15032,n15236,n15237 );
   nand U15044 ( n15230,n15033,p2_datao_reg_30_ );
   nand U15045 ( n15229,n15029,n11804 );
   nand U15046 ( n15240,n15029,n11811 );
   nand U15047 ( n15239,n15032,n15237,n15235 );
   not U15048 ( n15235,n15236 );
   nand U15049 ( n15236,n15227,n15228 );
   nand U15050 ( n15061,p1_state_reg,n15241 );
   nand U15051 ( n15238,n15033,p2_datao_reg_31_ );
   nand U15052 ( n14973,n14541,n15252 );
   nor U15053 ( n15259,n14927,n15260 );
   nor U15054 ( n15258,n15261,n15262 );
   nor U15055 ( n15262,n14991,n14994 );
   nor U15056 ( n15257,n15263,n14986 );
   nand U15057 ( n15255,n14990,p1_reg3_reg_0_ );
   nand U15058 ( n15254,p1_reg2_reg_0_,n14995 );
   nand U15059 ( n15253,n14996,n14958 );
   nand U15060 ( n14958,n15264,n15265 );
   nand U15061 ( n15265,n15266,n14626 );
   nand U15062 ( n15266,n15267,n15268 );
   nand U15063 ( n15264,n14957,n15020 );
   not U15064 ( n14957,n15263 );
   and U15065 ( n15276,n15277,n14947 );
   xor U15066 ( n14947,n15278,n15279 );
   nor U15067 ( n15275,n14942,n15280 );
   and U15068 ( n15274,n14946,n14991 );
   xor U15069 ( n14946,n14956,n15281 );
   nor U15070 ( n15273,n14945,n15282 );
   nand U15071 ( n14945,n15283,n15284 );
   nand U15072 ( n15284,n15267,n15279 );
   nand U15073 ( n15279,n15285,n15286 );
   nand U15074 ( n15283,n15287,n15288 );
   nor U15075 ( n15271,n15289,n15290 );
   nor U15076 ( n15290,n14996,n15291 );
   nor U15077 ( n15289,n14943,n15292 );
   nand U15078 ( n15270,n15293,n14435 );
   nand U15079 ( n15269,n14990,p1_reg3_reg_1_ );
   nor U15080 ( n15301,n14900,n15260 );
   nand U15081 ( n14929,n15303,n15304 );
   nand U15082 ( n15304,n15305,n15306 );
   nand U15083 ( n15305,n14943,n15261 );
   nor U15084 ( n15299,n15307,n14931 );
   nand U15085 ( n14931,n15308,n15309 );
   nand U15086 ( n15309,n15310,n15311 );
   nand U15087 ( n15308,n15312,n15313,n15314 );
   nor U15088 ( n15298,n14927,n15280 );
   nor U15089 ( n15296,n15315,n15316 );
   nor U15090 ( n15316,n14995,n14921 );
   nand U15091 ( n14921,n15317,n15318,n15319 );
   nand U15092 ( n15319,n15013,n15320,n15012 );
   nand U15093 ( n15318,n15321,n15313 );
   nand U15094 ( n15317,n15310,n15322 );
   nor U15095 ( n15315,n14996,n15323 );
   nand U15096 ( n15295,n14990,p1_reg3_reg_2_ );
   nand U15097 ( n15294,n14994,n15306 );
   nor U15098 ( n15331,n14884,n15260 );
   and U15099 ( n15330,n15277,n14917 );
   xor U15100 ( n14917,n15332,n15333 );
   nand U15101 ( n15333,n15334,n15335 );
   nand U15102 ( n15335,n15336,n14435 );
   nand U15103 ( n15336,n15314,n14928 );
   not U15104 ( n15314,n15311 );
   nand U15105 ( n15334,n15311,n15306 );
   nand U15106 ( n15311,n15286,n15337 );
   nor U15107 ( n15329,n14941,n15280 );
   and U15108 ( n15328,n14916,n14991 );
   xor U15109 ( n14916,n15303,n15338 );
   nor U15110 ( n15326,n15339,n15340 );
   and U15111 ( n15340,n14912,n14996 );
   nand U15112 ( n14912,n15341,n15342 );
   nand U15113 ( n15342,n15343,n15344 );
   nand U15114 ( n15343,n15012,n15320 );
   not U15115 ( n15012,n15345 );
   nand U15116 ( n15341,n15346,n15344 );
   nand U15117 ( n15344,n15347,n15348 );
   or U15118 ( n15348,n15332,n15349 );
   nand U15119 ( n15347,n15332,n15349 );
   and U15120 ( n15339,n14995,p1_reg2_reg_3_ );
   nand U15121 ( n15325,n14990,n15350 );
   nand U15122 ( n15324,n14994,n15338 );
   nor U15123 ( n15358,n15307,n14904 );
   xor U15124 ( n14904,n15359,n15360 );
   not U15125 ( n15307,n15277 );
   nor U15126 ( n15357,n14900,n15280 );
   nor U15127 ( n15356,n15361,n15362 );
   nor U15128 ( n15355,n15363,n15282 );
   not U15129 ( n15363,n14905 );
   nand U15130 ( n14905,n15364,n15365 );
   nand U15131 ( n15365,n15366,n15359 );
   not U15132 ( n15366,n15367 );
   nand U15133 ( n15364,n15368,n15367 );
   nand U15134 ( n15368,n15369,n15370 );
   nor U15135 ( n15353,n15371,n15372 );
   nor U15136 ( n15372,n14899,n15260 );
   nand U15137 ( n14902,n15373,n15374 );
   nand U15138 ( n15374,n15375,n15376 );
   nand U15139 ( n15375,n15377,n14915 );
   nand U15140 ( n15352,n14994,n15376 );
   nand U15141 ( n15351,p1_reg2_reg_4_,n14995 );
   and U15142 ( n15385,n15277,n14889 );
   xor U15143 ( n14889,n15386,n15387 );
   nor U15144 ( n15386,n15388,n15389 );
   not U15145 ( n15389,n15390 );
   nor U15146 ( n15388,n15391,n15360 );
   nor U15147 ( n15384,n14884,n15280 );
   and U15148 ( n15383,n14888,n14991 );
   xor U15149 ( n14888,n15392,n15373 );
   nor U15150 ( n15382,n14887,n15282 );
   nand U15151 ( n14887,n15393,n15394 );
   nand U15152 ( n15394,n15395,n15396,n15397 );
   nand U15153 ( n15393,n15387,n15398 );
   nor U15154 ( n15380,n15399,n15400 );
   nor U15155 ( n15400,n14996,n15401 );
   nor U15156 ( n15399,n14885,n15292 );
   nand U15157 ( n15379,n15293,n14423 );
   nand U15158 ( n15378,n14990,n15402 );
   nor U15159 ( n15410,n15411,n15292 );
   nor U15160 ( n15409,n15412,n15362 );
   nor U15161 ( n15408,n14864,n14995 );
   and U15162 ( n14864,n15413,n15414 );
   nor U15163 ( n15414,n15415,n15416,n15417,n15418 );
   nor U15164 ( n15418,n15419,n15013 );
   nor U15165 ( n15417,n15420,n14870 );
   nor U15166 ( n15416,n15419,n15320 );
   nor U15167 ( n15415,n15419,n15421 );
   nor U15168 ( n15413,n15422,n15423,n15424,n15425 );
   nor U15169 ( n15425,n14899,n14622 );
   nor U15170 ( n15424,n15426,n14870 );
   nor U15171 ( n15423,n15419,n15427 );
   nor U15172 ( n15419,n15428,n15429 );
   nor U15173 ( n15429,n15430,n15431 );
   nand U15174 ( n15431,n15432,n15433 );
   nand U15175 ( n15433,n15398,n15396 );
   not U15176 ( n15398,n15397 );
   not U15177 ( n15432,n15434 );
   nor U15178 ( n15428,n15435,n15436 );
   nor U15179 ( n15422,n15437,n14870 );
   nor U15180 ( n15407,n14996,n15438 );
   nand U15181 ( n15405,n15293,n14420 );
   or U15182 ( n15404,n15302,n14871 );
   nand U15183 ( n14871,n15439,n15440 );
   nand U15184 ( n15440,n15441,n14873 );
   nand U15185 ( n15441,n15442,n14885 );
   or U15186 ( n15403,n14986,n14870 );
   xor U15187 ( n14870,n15434,n15443 );
   nor U15188 ( n15451,n15452,n15292 );
   and U15189 ( n15450,n15453,n14990 );
   nor U15190 ( n15449,n14853,n14995 );
   and U15191 ( n14853,n15454,n15455,n15456,n15457 );
   nor U15192 ( n15457,n15458,n15459,n15460,n15461 );
   nor U15193 ( n15461,n15426,n14859 );
   nor U15194 ( n15460,n15420,n14859 );
   nor U15195 ( n15459,n15437,n14859 );
   nor U15196 ( n15458,n15013,n15462 );
   nor U15197 ( n15456,n15463,n15464 );
   nor U15198 ( n15464,n14883,n14622 );
   nand U15199 ( n15455,n15465,n15466 );
   nand U15200 ( n15454,n15465,n15014 );
   not U15201 ( n15465,n15462 );
   nand U15202 ( n15462,n15467,n15468 );
   nand U15203 ( n15468,n15469,n15470 );
   nand U15204 ( n15467,n15471,n15472 );
   nor U15205 ( n15448,n14996,n15473 );
   nand U15206 ( n15446,n15293,n14417 );
   nand U15207 ( n15445,n14991,n14860 );
   xor U15208 ( n14860,n15439,n14861 );
   or U15209 ( n15444,n14986,n14859 );
   nand U15210 ( n14859,n15474,n15475 );
   nand U15211 ( n15475,n15476,n15477,n15478 );
   nand U15212 ( n15474,n15479,n15480,n15471 );
   nand U15213 ( n15479,n15481,n15477 );
   not U15214 ( n15481,n15443 );
   nor U15215 ( n15489,n15490,n15292 );
   nor U15216 ( n15488,n15491,n15362 );
   nor U15217 ( n15487,n14841,n14995 );
   and U15218 ( n14841,n15492,n15493,n15494,n15495 );
   nor U15219 ( n15495,n15496,n15497,n15498,n15499 );
   nor U15220 ( n15499,n15500,n15320 );
   xor U15221 ( n15500,n15501,n15502 );
   nor U15222 ( n15498,n15503,n15013 );
   nor U15223 ( n15503,n15504,n15505 );
   nor U15224 ( n15504,n15506,n15507 );
   nor U15225 ( n15506,n15508,n15469 );
   nor U15226 ( n15497,n15437,n14847 );
   not U15227 ( n14847,n15509 );
   nor U15228 ( n15496,n14872,n14622 );
   nand U15229 ( n15494,n15509,n15510 );
   nand U15230 ( n15493,n15345,n15511 );
   nand U15231 ( n15511,n15512,n15513 );
   not U15232 ( n15513,n15505 );
   nor U15233 ( n15505,n15501,n15502 );
   nand U15234 ( n15512,n15502,n15501 );
   nand U15235 ( n15492,n15509,n15514 );
   nor U15236 ( n15486,n14996,n15515 );
   nand U15237 ( n15484,n15293,n14414 );
   or U15238 ( n15483,n15302,n14848 );
   nand U15239 ( n14848,n15516,n15517 );
   nand U15240 ( n15517,n15518,n14850 );
   nand U15241 ( n15518,n15519,n15452 );
   nand U15242 ( n15482,n15520,n15509 );
   xor U15243 ( n15509,n15502,n15521 );
   and U15244 ( n15529,n15277,n14838 );
   xor U15245 ( n14838,n15530,n15531 );
   nor U15246 ( n15528,n14834,n15280 );
   and U15247 ( n15527,n14837,n14991 );
   xor U15248 ( n14837,n15532,n15516 );
   nor U15249 ( n15526,n15533,n15282 );
   not U15250 ( n15533,n14836 );
   nand U15251 ( n14836,n15534,n15535 );
   nand U15252 ( n15535,n15536,n15530 );
   not U15253 ( n15536,n15537 );
   nand U15254 ( n15534,n15538,n15537 );
   nand U15255 ( n15538,n15539,n15540 );
   nor U15256 ( n15524,n15541,n15542 );
   nor U15257 ( n15542,n14996,n15543 );
   nor U15258 ( n15541,n14835,n15292 );
   nand U15259 ( n15523,n15293,n14411 );
   nand U15260 ( n15522,n14990,n15544 );
   nor U15261 ( n15552,n15553,n15292 );
   nor U15262 ( n15551,n15554,n15362 );
   nor U15263 ( n15550,n14815,n14995 );
   and U15264 ( n14815,n15555,n15556,n15557,n15558 );
   nor U15265 ( n15558,n15559,n15560,n15561,n15562 );
   nor U15266 ( n15562,n15427,n15563 );
   nor U15267 ( n15561,n15426,n14821 );
   nor U15268 ( n15560,n15420,n14821 );
   nor U15269 ( n15559,n15437,n14821 );
   nand U15270 ( n15557,n15564,n15466 );
   nand U15271 ( n15556,n15564,n15565 );
   nand U15272 ( n15565,n15013,n15320 );
   not U15273 ( n15564,n15563 );
   nand U15274 ( n15563,n15566,n15567 );
   nand U15275 ( n15567,n15568,n15569,n15570 );
   nand U15276 ( n15566,n15571,n15572 );
   nand U15277 ( n15555,n14771,n14414 );
   nor U15278 ( n15549,n14996,n15573 );
   nand U15279 ( n15547,n15293,n14408 );
   or U15280 ( n15546,n15302,n14822 );
   nand U15281 ( n14822,n15574,n15575 );
   nand U15282 ( n15575,n15576,n14823 );
   or U15283 ( n15545,n14986,n14821 );
   nand U15284 ( n14821,n15577,n15578 );
   nand U15285 ( n15578,n15579,n15580,n15581 );
   nand U15286 ( n15577,n15582,n15583,n15571 );
   nand U15287 ( n15582,n15531,n15580 );
   not U15288 ( n15531,n15584 );
   nor U15289 ( n15592,n15593,n15292 );
   nor U15290 ( n15591,n15594,n15362 );
   nor U15291 ( n15590,n14803,n14995 );
   and U15292 ( n14803,n15595,n15596 );
   nor U15293 ( n15596,n15597,n15598,n15599,n15600 );
   nor U15294 ( n15600,n15601,n15013 );
   nor U15295 ( n15599,n15437,n14809 );
   nor U15296 ( n15598,n14833,n14622 );
   nor U15297 ( n15597,n15601,n15421 );
   nor U15298 ( n15595,n15602,n15603,n15604,n15605 );
   nor U15299 ( n15605,n15601,n15427 );
   and U15300 ( n15601,n15606,n15607,n15608 );
   not U15301 ( n15608,n15609 );
   nand U15302 ( n15607,n15610,n15570 );
   nand U15303 ( n15606,n15572,n15611 );
   nor U15304 ( n15604,n15426,n14809 );
   nor U15305 ( n15603,n15420,n14809 );
   not U15306 ( n14809,n15612 );
   nor U15307 ( n15602,n15613,n15320 );
   nor U15308 ( n15613,n15609,n15614,n15615 );
   nor U15309 ( n15615,n15616,n15570 );
   nor U15310 ( n15614,n15572,n15617 );
   not U15311 ( n15572,n15570 );
   nand U15312 ( n15570,n15540,n15618 );
   nand U15313 ( n15618,n15539,n15537 );
   nand U15314 ( n15609,n15619,n15620 );
   nand U15315 ( n15620,n15621,n15610 );
   not U15316 ( n15610,n15617 );
   nand U15317 ( n15617,n15622,n15568 );
   nand U15318 ( n15619,n15623,n15611 );
   not U15319 ( n15611,n15616 );
   nand U15320 ( n15616,n15624,n15625 );
   nor U15321 ( n15589,n14996,n15626 );
   nand U15322 ( n15587,n15293,n14405 );
   nand U15323 ( n15586,n14991,n14810 );
   xor U15324 ( n14810,n14812,n15574 );
   not U15325 ( n15574,n15627 );
   nand U15326 ( n15585,n15520,n15612 );
   xor U15327 ( n15612,n15622,n15628 );
   nand U15328 ( n14797,n15637,n15638 );
   nand U15329 ( n15638,n15639,n15640 );
   nand U15330 ( n15639,n15593,n15627 );
   and U15331 ( n15635,n15277,n14798 );
   xor U15332 ( n14798,n15641,n15642 );
   nor U15333 ( n15634,n14795,n15280 );
   nor U15334 ( n15633,n14800,n15282 );
   xor U15335 ( n14800,n15641,n15643 );
   nor U15336 ( n15631,n15644,n15645 );
   nor U15337 ( n15645,n14996,n15646 );
   nor U15338 ( n15644,n14796,n15292 );
   nand U15339 ( n15630,n15293,n14402 );
   nand U15340 ( n15629,n14990,n15647 );
   nor U15341 ( n15655,n15656,n15292 );
   nor U15342 ( n15654,n15657,n15362 );
   nor U15343 ( n15653,n14776,n14995 );
   and U15344 ( n14776,n15658,n15659,n15660,n15661 );
   nor U15345 ( n15661,n15662,n15663,n15664,n15665 );
   nor U15346 ( n15665,n15426,n14782 );
   nor U15347 ( n15664,n15420,n14782 );
   nor U15348 ( n15663,n15437,n14782 );
   nor U15349 ( n15662,n15320,n15666 );
   nor U15350 ( n15660,n15667,n15668 );
   nor U15351 ( n15668,n14811,n14622 );
   not U15352 ( n15666,n15669 );
   nand U15353 ( n15659,n15669,n15466 );
   nand U15354 ( n15658,n15669,n15346 );
   xor U15355 ( n15669,n15670,n15671 );
   nor U15356 ( n15652,n14996,n15672 );
   nand U15357 ( n15650,n15293,n14399 );
   nand U15358 ( n15649,n14991,n14783 );
   xor U15359 ( n14783,n15637,n14784 );
   or U15360 ( n15648,n14986,n14782 );
   nand U15361 ( n14782,n15673,n15674 );
   nand U15362 ( n15674,n15675,n15676,n15677 );
   nand U15363 ( n15675,n15678,n15679 );
   not U15364 ( n15679,n15642 );
   nand U15365 ( n15673,n15680,n15678,n15670 );
   nand U15366 ( n15680,n15642,n15676 );
   nor U15367 ( n15642,n15681,n15682 );
   nor U15368 ( n15686,n15687,n15688,n15689,n15690 );
   nor U15369 ( n15690,n14770,n15260 );
   nand U15370 ( n14773,n15691,n15692 );
   nand U15371 ( n15692,n15693,n15694 );
   nand U15372 ( n15693,n15695,n15656 );
   and U15373 ( n15688,n15277,n14772 );
   xor U15374 ( n14772,n15696,n15697 );
   nor U15375 ( n15687,n14794,n15280 );
   nor U15376 ( n15685,n15698,n15699 );
   nor U15377 ( n15699,n14769,n15292 );
   nor U15378 ( n15698,n15700,n15362 );
   nand U15379 ( n15684,p1_reg2_reg_14_,n14995 );
   nand U15380 ( n14766,n15701,n15702 );
   nand U15381 ( n15702,n15703,n15704,n15466 );
   nand U15382 ( n15703,n15705,n15706 );
   nand U15383 ( n15701,n15707,n15704,n15708 );
   nand U15384 ( n15704,n15697,n15709 );
   or U15385 ( n15707,n15710,n15711,n15709 );
   nor U15386 ( n15715,n15716,n15717,n15718,n15719 );
   nor U15387 ( n15719,n14755,n15260 );
   and U15388 ( n15718,n15277,n14758 );
   xor U15389 ( n14758,n15720,n15721 );
   nor U15390 ( n15717,n14756,n15280 );
   and U15391 ( n15716,n14759,n14991 );
   xor U15392 ( n14759,n15722,n15691 );
   nor U15393 ( n15714,n15723,n15724 );
   nor U15394 ( n15724,n14995,n14749 );
   nand U15395 ( n14749,n15725,n15726,n14626 );
   nand U15396 ( n15726,n15727,n15728 );
   nand U15397 ( n15725,n15729,n15721 );
   nor U15398 ( n15723,n14996,n15730 );
   nand U15399 ( n15713,n14990,n15731 );
   nand U15400 ( n15712,n14994,n15722 );
   nor U15401 ( n15739,n15740,n15292 );
   nor U15402 ( n15738,n15741,n15362 );
   nor U15403 ( n15737,n14737,n14995 );
   and U15404 ( n14737,n15742,n15743 );
   nor U15405 ( n15743,n15744,n15745,n15746,n15747 );
   nor U15406 ( n15747,n15013,n15748,n15749 );
   nor U15407 ( n15749,n15750,n15751 );
   nor U15408 ( n15751,n15752,n15753,n15754 );
   and U15409 ( n15754,n15728,n15729 );
   and U15410 ( n15748,n15752,n15727 );
   nor U15411 ( n15746,n15755,n15320 );
   nor U15412 ( n15745,n14743,n15426 );
   nor U15413 ( n15744,n15755,n15421 );
   nor U15414 ( n15742,n15756,n15757,n15758,n15759 );
   nor U15415 ( n15759,n14743,n15420 );
   nor U15416 ( n15758,n14743,n15437 );
   nor U15417 ( n15757,n15755,n15427 );
   and U15418 ( n15755,n15760,n15761,n15762,n15763 );
   nand U15419 ( n15763,n15764,n15727 );
   nor U15420 ( n15727,n15729,n15753 );
   nand U15421 ( n15762,n15729,n15750 );
   nor U15422 ( n15729,n15705,n15711 );
   nand U15423 ( n15761,n15753,n15750 );
   nor U15424 ( n15750,n15765,n15766 );
   not U15425 ( n15753,n15767 );
   nand U15426 ( n15760,n15768,n15764 );
   nor U15427 ( n15756,n14770,n14622 );
   nor U15428 ( n15736,n14996,n15769 );
   nand U15429 ( n15734,n15293,n14390 );
   or U15430 ( n15733,n15302,n14744 );
   nand U15431 ( n14744,n15770,n15771 );
   nand U15432 ( n15771,n15772,n14745 );
   nand U15433 ( n15772,n15773,n14757 );
   or U15434 ( n15732,n14986,n14743 );
   xor U15435 ( n14743,n15764,n15774 );
   not U15436 ( n15764,n15752 );
   nor U15437 ( n15782,n15783,n15292 );
   nor U15438 ( n15781,n15784,n15362 );
   nor U15439 ( n15780,n14726,n14995 );
   and U15440 ( n14726,n15785,n15786,n15787,n15788 );
   nor U15441 ( n15788,n15789,n15790,n15791,n15792 );
   nor U15442 ( n15792,n15793,n15013 );
   nor U15443 ( n15791,n15793,n15421 );
   nor U15444 ( n15790,n14755,n14622 );
   nor U15445 ( n15789,n15793,n15427 );
   nor U15446 ( n15787,n15794,n15795 );
   nor U15447 ( n15795,n15437,n14732 );
   nor U15448 ( n15794,n15793,n15320 );
   xor U15449 ( n15793,n15796,n15797 );
   nand U15450 ( n15786,n15798,n15514 );
   nand U15451 ( n15785,n15798,n15510 );
   nor U15452 ( n15779,n14996,n15799 );
   nand U15453 ( n15777,n15293,n14387 );
   nand U15454 ( n15776,n14991,n14733 );
   xor U15455 ( n14733,n15770,n14734 );
   nand U15456 ( n15775,n15520,n15798 );
   not U15457 ( n15798,n14732 );
   nand U15458 ( n14732,n15800,n15801 );
   nand U15459 ( n15801,n15802,n15803,n15804 );
   nand U15460 ( n15800,n15805,n15806,n15796 );
   nand U15461 ( n15805,n15803,n15774 );
   nor U15462 ( n15810,n15811,n15812,n15813,n15814 );
   nor U15463 ( n15814,n14996,n15815 );
   nor U15464 ( n15813,n14720,n15292 );
   nor U15465 ( n15812,n15816,n15362 );
   nor U15466 ( n15811,n14718,n15260 );
   nor U15467 ( n15809,n15817,n15818 );
   nor U15468 ( n15818,n14719,n15280 );
   nor U15469 ( n15817,n15819,n15282 );
   not U15470 ( n15819,n14723 );
   xor U15471 ( n14723,n15820,n15821 );
   nand U15472 ( n15808,n14722,n15277 );
   xor U15473 ( n14722,n15820,n15822 );
   nand U15474 ( n15807,n14991,n14721 );
   and U15475 ( n14721,n15823,n15824 );
   nand U15476 ( n15824,n15825,n15826 );
   nand U15477 ( n15825,n15827,n15783 );
   nor U15478 ( n15831,n15832,n15833,n15834,n15835 );
   nor U15479 ( n15835,n14996,n15836 );
   nor U15480 ( n15834,n14705,n15292 );
   nor U15481 ( n15833,n15837,n15362 );
   nor U15482 ( n15832,n14703,n15260 );
   nor U15483 ( n15830,n15838,n15839 );
   and U15484 ( n15839,n14707,n14991 );
   xor U15485 ( n14707,n15840,n15823 );
   nor U15486 ( n15838,n15841,n15282 );
   not U15487 ( n15841,n14706 );
   xor U15488 ( n14706,n15842,n15843 );
   nand U15489 ( n15829,n15844,n14387 );
   nand U15490 ( n15828,n14708,n15277 );
   xor U15491 ( n14708,n15842,n15845 );
   nor U15492 ( n15853,n15854,n15292 );
   nor U15493 ( n15852,n15855,n15362 );
   nor U15494 ( n15851,n14685,n14995 );
   and U15495 ( n14685,n15856,n15857,n15858,n15859 );
   nor U15496 ( n15859,n15860,n15861,n15862,n15863 );
   nor U15497 ( n15863,n15013,n15864 );
   nor U15498 ( n15862,n15421,n15864 );
   nor U15499 ( n15861,n14718,n14622 );
   nor U15500 ( n15860,n15427,n15864 );
   nor U15501 ( n15858,n15865,n15866 );
   nor U15502 ( n15866,n15426,n14691 );
   nor U15503 ( n15865,n15420,n14691 );
   or U15504 ( n15857,n15864,n15320 );
   xor U15505 ( n15864,n15867,n15868 );
   nand U15506 ( n15856,n15869,n15870 );
   and U15507 ( n15850,n14995,p1_reg2_reg_20_ );
   nand U15508 ( n15848,n15293,n14378 );
   or U15509 ( n15847,n15302,n14692 );
   nand U15510 ( n14692,n15871,n15872 );
   nand U15511 ( n15872,n15873,n14693 );
   nand U15512 ( n15873,n15874,n14705 );
   nand U15513 ( n15846,n15520,n15869 );
   not U15514 ( n15869,n14691 );
   nand U15515 ( n14691,n15875,n15876 );
   nand U15516 ( n15876,n15877,n15878,n15879 );
   nand U15517 ( n15877,n15880,n15881 );
   nand U15518 ( n15875,n15867,n15881,n15882 );
   nand U15519 ( n15882,n15845,n15883 );
   nor U15520 ( n15891,n14679,n15292 );
   and U15521 ( n15890,n15892,n14990 );
   and U15522 ( n15889,n14678,n14996 );
   nand U15523 ( n14678,n15893,n15894,n15895,n15896 );
   nor U15524 ( n15896,n15897,n15898 );
   nor U15525 ( n15898,n14703,n14622 );
   nor U15526 ( n15897,n15899,n15900,n15901 );
   nor U15527 ( n15901,n15902,n15903,n15904 );
   nor U15528 ( n15900,n15905,n15906 );
   nand U15529 ( n15895,n14681,n15907 );
   nand U15530 ( n15894,n15510,n15908,n15909,n15910 );
   nand U15531 ( n15893,n15911,n15912,n15466 );
   not U15532 ( n15466,n15421 );
   nand U15533 ( n15912,n15913,n15902 );
   nand U15534 ( n15911,n15914,n15915,n15905 );
   and U15535 ( n15888,n14995,p1_reg2_reg_21_ );
   nand U15536 ( n15886,n15293,n14375 );
   nand U15537 ( n15885,n14991,n14680 );
   xor U15538 ( n14680,n15916,n14679 );
   nand U15539 ( n15884,n15520,n14681 );
   and U15540 ( n14681,n15909,n15910,n15908 );
   nand U15541 ( n15908,n15879,n15845,n15913 );
   nand U15542 ( n15910,n15913,n15917 );
   nand U15543 ( n15909,n15918,n15906,n15919 );
   nand U15544 ( n15918,n15879,n15845 );
   not U15545 ( n15845,n15880 );
   nor U15546 ( n15880,n15920,n15921 );
   nor U15547 ( n15925,n15926,n15927,n15928,n15929 );
   nor U15548 ( n15929,n14641,n15260 );
   nand U15549 ( n14669,n15930,n15931 );
   nand U15550 ( n15931,n15932,n15933 );
   nand U15551 ( n15932,n15916,n14679 );
   and U15552 ( n15927,n15277,n14670 );
   xor U15553 ( n14670,n15934,n15935 );
   nor U15554 ( n15926,n14667,n15280 );
   nor U15555 ( n15924,n15936,n15937 );
   nor U15556 ( n15937,n14995,n14661 );
   nand U15557 ( n14661,n15938,n15939,n14626 );
   nand U15558 ( n15939,n15940,n15941,n15942 );
   nand U15559 ( n15938,n15934,n15943 );
   not U15560 ( n15934,n15944 );
   and U15561 ( n15936,n14995,p1_reg2_reg_22_ );
   nand U15562 ( n15923,n14990,n15945 );
   nand U15563 ( n15922,n14994,n15933 );
   nor U15564 ( n15953,n15954,n15292 );
   and U15565 ( n15952,n15955,n14990 );
   nor U15566 ( n15951,n14649,n14995 );
   and U15567 ( n14649,n15956,n15957,n15958,n15959 );
   nor U15568 ( n15959,n15960,n15961,n15962,n15963 );
   nor U15569 ( n15963,n15013,n15964,n15965 );
   nor U15570 ( n15965,n15966,n15967 );
   nor U15571 ( n15967,n15968,n15969 );
   nor U15572 ( n15968,n15970,n15942 );
   and U15573 ( n15964,n15971,n15941,n15942 );
   nor U15574 ( n15962,n14655,n15420 );
   nor U15575 ( n15961,n15972,n15320 );
   nor U15576 ( n15960,n15972,n15427 );
   nor U15577 ( n15958,n15973,n15974 );
   nor U15578 ( n15974,n15975,n14622 );
   nor U15579 ( n15973,n15972,n15421 );
   and U15580 ( n15972,n15976,n15977 );
   nand U15581 ( n15977,n15978,n15979 );
   nand U15582 ( n15979,n15943,n15940 );
   not U15583 ( n15943,n15942 );
   not U15584 ( n15978,n15969 );
   nand U15585 ( n15969,n15980,n15941 );
   nand U15586 ( n15976,n15966,n15981 );
   nand U15587 ( n15981,n15941,n15942 );
   nand U15588 ( n15942,n15915,n15982 );
   nand U15589 ( n15982,n15905,n15914 );
   and U15590 ( n15966,n15983,n15984 );
   nand U15591 ( n15957,n15510,n15985 );
   nand U15592 ( n15956,n15870,n15985 );
   and U15593 ( n15950,n14995,p1_reg2_reg_23_ );
   nand U15594 ( n15948,n15293,n14369 );
   nand U15595 ( n15947,n14991,n14656 );
   xor U15596 ( n14656,n14657,n15930 );
   nand U15597 ( n15946,n15520,n15985 );
   not U15598 ( n15985,n14655 );
   xor U15599 ( n14655,n15980,n15986 );
   not U15600 ( n15980,n15971 );
   nor U15601 ( n15990,n15991,n15992,n15993,n15994 );
   and U15602 ( n15994,n14995,p1_reg2_reg_24_ );
   nor U15603 ( n15993,n14642,n15292 );
   and U15604 ( n15992,n15995,n14990 );
   nor U15605 ( n15991,n14640,n15260 );
   nor U15606 ( n15989,n15996,n15997 );
   nor U15607 ( n15997,n14641,n15280 );
   nor U15608 ( n15996,n14646,n15282 );
   xor U15609 ( n14646,n15998,n15999 );
   nand U15610 ( n15988,n14644,n15277 );
   xor U15611 ( n14644,n16000,n15999 );
   nand U15612 ( n15987,n14991,n14643 );
   and U15613 ( n14643,n16001,n16002 );
   nand U15614 ( n16002,n16003,n16004 );
   nand U15615 ( n16003,n16005,n15954 );
   nor U15616 ( n16009,n16010,n16011,n16012,n16013 );
   and U15617 ( n16013,n14995,p1_reg2_reg_25_ );
   nor U15618 ( n16012,n14624,n15292 );
   and U15619 ( n16011,n16014,n14990 );
   nor U15620 ( n16010,n14620,n15260 );
   nor U15621 ( n16008,n16015,n16016 );
   and U15622 ( n16016,n14628,n14991 );
   xor U15623 ( n14628,n16001,n16017 );
   nor U15624 ( n16015,n14627,n15282 );
   nand U15625 ( n15282,n14996,n14626 );
   nand U15626 ( n14626,n15899,n15421 );
   not U15627 ( n15899,n15708 );
   nand U15628 ( n15708,n15013,n15320,n15427 );
   xor U15629 ( n14627,n16018,n16019 );
   nand U15630 ( n16007,n15844,n14369 );
   not U15631 ( n15844,n15280 );
   nand U15632 ( n15280,n14996,n14771 );
   not U15633 ( n14771,n14622 );
   nand U15634 ( n16006,n14629,n15277 );
   nand U15635 ( n15277,n14986,n16020 );
   nand U15636 ( n16020,n14996,n15020 );
   not U15637 ( n15020,n14948 );
   nor U15638 ( n14948,n15907,n15510 );
   nand U15639 ( n15907,n15437,n15420 );
   xor U15640 ( n14629,n16021,n16018 );
   nor U15641 ( n16029,n16030,n15292 );
   nor U15642 ( n16028,n16031,n15362 );
   nor U15643 ( n16027,n14600,n14995 );
   and U15644 ( n14600,n16032,n16033,n16034,n16035 );
   nor U15645 ( n16035,n16036,n16037,n16038,n16039 );
   nor U15646 ( n16039,n15320,n16040 );
   nor U15647 ( n16038,n15421,n16040 );
   nor U15648 ( n16037,n14640,n14622 );
   nor U15649 ( n16034,n16041,n16042 );
   nor U15650 ( n16042,n15437,n14606 );
   nor U15651 ( n16041,n15013,n16040 );
   nand U15652 ( n16040,n16043,n16044 );
   nand U15653 ( n16044,n16045,n16046 );
   nand U15654 ( n16043,n16047,n16048 );
   nand U15655 ( n16033,n16049,n15514 );
   nand U15656 ( n16032,n16049,n15510 );
   and U15657 ( n16026,n14995,p1_reg2_reg_26_ );
   nand U15658 ( n16024,n15293,n14360 );
   or U15659 ( n16023,n15302,n14608 );
   nand U15660 ( n14608,n16050,n16051 );
   nand U15661 ( n16051,n16052,n14610 );
   nand U15662 ( n16052,n16053,n14624 );
   nand U15663 ( n16022,n15520,n16049 );
   not U15664 ( n16049,n14606 );
   nand U15665 ( n14606,n16054,n16055 );
   nand U15666 ( n16055,n16056,n16057,n16058 );
   nand U15667 ( n16056,n16059,n16060 );
   not U15668 ( n16059,n16021 );
   nand U15669 ( n16054,n16061,n16060,n16047 );
   not U15670 ( n16047,n16058 );
   nand U15671 ( n16061,n16057,n16021 );
   nand U15672 ( n16021,n16062,n16063 );
   nand U15673 ( n16063,n16064,n16000 );
   nor U15674 ( n16072,n16073,n15292 );
   and U15675 ( n16071,n16074,n14990 );
   nor U15676 ( n16070,n14587,n14995 );
   and U15677 ( n14587,n16075,n16076,n16077,n16078 );
   nor U15678 ( n16078,n16079,n16080,n16081,n16082 );
   nor U15679 ( n16082,n15013,n16083,n16084 );
   nor U15680 ( n16084,n16085,n16086 );
   nor U15681 ( n16085,n16087,n16088 );
   and U15682 ( n16087,n16046,n16048 );
   nor U15683 ( n16083,n16089,n16090 );
   nor U15684 ( n16081,n15420,n14593 );
   and U15685 ( n16080,n16091,n15014 );
   nor U15686 ( n16079,n15426,n14593 );
   not U15687 ( n14593,n16092 );
   nor U15688 ( n16077,n16093,n16094 );
   nor U15689 ( n16094,n14620,n14622 );
   nor U15690 ( n16093,n16095,n15421 );
   xor U15691 ( n16095,n16090,n16086 );
   nand U15692 ( n16076,n16096,n16091 );
   xor U15693 ( n16091,n16090,n16089 );
   and U15694 ( n16090,n16046,n16097 );
   nand U15695 ( n16075,n16092,n15870 );
   and U15696 ( n16069,n14995,p1_reg2_reg_27_ );
   nand U15697 ( n16067,n15293,n14357 );
   nand U15698 ( n16066,n14991,n14594 );
   xor U15699 ( n14594,n16050,n14597 );
   nand U15700 ( n16065,n15520,n16092 );
   xor U15701 ( n16092,n16089,n16098 );
   nand U15702 ( n16098,n16099,n16100,n16101 );
   nand U15703 ( n16099,n16102,n16060,n16103 );
   not U15704 ( n16089,n16086 );
   nor U15705 ( n16111,n16112,n15292 );
   and U15706 ( n16110,n16113,n14990 );
   not U15707 ( n14990,n15362 );
   nand U15708 ( n15362,n14996,n16114 );
   nor U15709 ( n16109,n14575,n14995 );
   and U15710 ( n14575,n16115,n16116,n16117,n16118 );
   nor U15711 ( n16118,n16119,n16120,n16121,n16122 );
   nor U15712 ( n16122,n15320,n16123 );
   nor U15713 ( n16121,n16123,n15013 );
   nor U15714 ( n16120,n16123,n15421 );
   nor U15715 ( n16119,n14582,n15437 );
   nor U15716 ( n16117,n16124,n16125 );
   nor U15717 ( n16125,n16123,n15427 );
   xor U15718 ( n16123,n16126,n15018 );
   nand U15719 ( n15018,n16127,n16128 );
   nand U15720 ( n16127,n16097,n16046,n16129 );
   not U15721 ( n16097,n16045 );
   nor U15722 ( n16045,n16048,n16088 );
   not U15723 ( n16088,n16130 );
   nand U15724 ( n16048,n16131,n16132 );
   nand U15725 ( n16132,n14640,n16133 );
   or U15726 ( n16133,n16019,n16017 );
   nand U15727 ( n16131,n16019,n16017 );
   nand U15728 ( n16019,n16134,n16135 );
   nand U15729 ( n16135,n15998,n16136 );
   and U15730 ( n15998,n16137,n16138 );
   nand U15731 ( n16138,n15984,n16139 );
   nand U15732 ( n16139,n15983,n16140 );
   nand U15733 ( n16140,n15903,n15941 );
   and U15734 ( n15983,n15940,n16141 );
   nand U15735 ( n16141,n15954,n14372 );
   nand U15736 ( n16137,n15905,n16142 );
   not U15737 ( n15905,n15902 );
   nand U15738 ( n15902,n16143,n16144 );
   nand U15739 ( n16144,n16145,n15868 );
   nand U15740 ( n15868,n16146,n16147 );
   nand U15741 ( n16147,n16148,n15843 );
   nand U15742 ( n15843,n16149,n16150 );
   nand U15743 ( n16150,n16151,n15821 );
   nand U15744 ( n15821,n16152,n16153 );
   or U15745 ( n16153,n15797,n16154 );
   nand U15746 ( n15797,n16155,n16156 );
   nand U15747 ( n16156,n16157,n16158 );
   nand U15748 ( n16158,n16159,n16160 );
   nand U15749 ( n16160,n15711,n15767 );
   not U15750 ( n16159,n15765 );
   nand U15751 ( n16155,n15705,n16161 );
   not U15752 ( n16161,n16162 );
   nor U15753 ( n15705,n15709,n15710 );
   or U15754 ( n15709,n16163,n16164 );
   and U15755 ( n16164,n16165,n15671 );
   nand U15756 ( n15671,n16166,n16167 );
   nand U15757 ( n16167,n15643,n16168 );
   and U15758 ( n15643,n16169,n16170 );
   nand U15759 ( n16170,n15539,n15537,n16171 );
   not U15760 ( n16171,n16172 );
   nand U15761 ( n15537,n16173,n16174 );
   nand U15762 ( n16174,n16175,n15501 );
   or U15763 ( n15501,n15508,n15469 );
   nor U15764 ( n15469,n15472,n16176 );
   nand U15765 ( n15472,n15435,n16177 );
   nand U15766 ( n15435,n16178,n15396,n16179 );
   nand U15767 ( n16179,n15395,n15397 );
   nand U15768 ( n15397,n16180,n15369 );
   nand U15769 ( n16180,n15367,n15370 );
   nand U15770 ( n15367,n16181,n16182 );
   nand U15771 ( n16182,n16183,n14432 );
   or U15772 ( n16183,n15349,n14915 );
   nand U15773 ( n16181,n14915,n15349 );
   not U15774 ( n15508,n15470 );
   nand U15775 ( n16175,n14834,n14850 );
   nand U15776 ( n16169,n16184,n15625 );
   nand U15777 ( n16184,n15624,n16185 );
   or U15778 ( n16185,n15540,n15623 );
   not U15779 ( n15623,n15568 );
   and U15780 ( n15624,n15569,n16186 );
   nand U15781 ( n16186,n15593,n14408 );
   nand U15782 ( n16165,n15656,n14402 );
   nand U15783 ( n16143,n14703,n14693 );
   nor U15784 ( n16124,n14609,n14622 );
   nand U15785 ( n16116,n15514,n16189 );
   nand U15786 ( n16115,n15510,n16189 );
   and U15787 ( n16108,n14995,p1_reg2_reg_28_ );
   nand U15788 ( n16106,n15520,n16189 );
   not U15789 ( n16189,n14582 );
   xor U15790 ( n14582,n16126,n15025 );
   nand U15791 ( n15025,n16190,n16191,n16192,n16193 );
   nand U15792 ( n16192,n16103,n16194,n16102,n16060 );
   nand U15793 ( n16103,n16057,n16064 );
   nand U15794 ( n16191,n16195,n16194 );
   not U15795 ( n16195,n16100 );
   nand U15796 ( n16100,n16196,n16062,n16102,n16060 );
   not U15797 ( n16196,n16000 );
   nand U15798 ( n16000,n16197,n16198 );
   nand U15799 ( n16198,n14641,n16199 );
   or U15800 ( n16199,n15986,n15954 );
   nand U15801 ( n16197,n15954,n15986 );
   nand U15802 ( n15986,n16200,n16201 );
   nand U15803 ( n16201,n15975,n16202 );
   nand U15804 ( n16202,n15933,n15935 );
   or U15805 ( n16200,n15935,n15933 );
   nand U15806 ( n15935,n16203,n16204,n16205 );
   nand U15807 ( n16205,n16206,n16207 );
   nand U15808 ( n16207,n15919,n16208 );
   nand U15809 ( n16208,n15920,n15879 );
   not U15810 ( n15919,n15917 );
   nand U15811 ( n15917,n15878,n16209 );
   nand U15812 ( n16209,n16210,n16211 );
   not U15813 ( n16210,n15881 );
   nand U15814 ( n16203,n15879,n16206,n15921 );
   and U15815 ( n15921,n16212,n15822 );
   nand U15816 ( n15822,n16213,n16214 );
   nand U15817 ( n16214,n16215,n16216 );
   nand U15818 ( n16215,n15803,n15802 );
   nand U15819 ( n15802,n16217,n15806 );
   not U15820 ( n16217,n15774 );
   nand U15821 ( n15774,n16218,n16219 );
   nand U15822 ( n16219,n14770,n16220 );
   nand U15823 ( n16220,n15720,n15722 );
   not U15824 ( n15720,n16221 );
   nand U15825 ( n16218,n14757,n16221 );
   nand U15826 ( n16221,n16222,n16223 );
   nand U15827 ( n16223,n14756,n16224 );
   nand U15828 ( n16224,n15694,n15696 );
   not U15829 ( n14756,n14399 );
   or U15830 ( n16222,n15696,n15694 );
   nand U15831 ( n15696,n16225,n16226 );
   nand U15832 ( n16226,n16227,n15678,n15681 );
   and U15833 ( n15681,n15628,n16228 );
   nand U15834 ( n16228,n14795,n15593 );
   nand U15835 ( n15628,n16229,n16230 );
   nand U15836 ( n16230,n16231,n16232 );
   nand U15837 ( n16231,n15580,n15579 );
   nand U15838 ( n15579,n15583,n15584 );
   nand U15839 ( n15584,n16233,n16234 );
   nand U15840 ( n16233,n15521,n16235 );
   nand U15841 ( n15521,n16236,n16237 );
   nand U15842 ( n16237,n16238,n16239 );
   nand U15843 ( n16239,n14872,n15452 );
   nand U15844 ( n16238,n15477,n15476 );
   nand U15845 ( n15476,n15443,n15480 );
   nand U15846 ( n15443,n16240,n16241,n16242 );
   nand U15847 ( n16242,n15391,n15392 );
   not U15848 ( n15391,n16243 );
   nand U15849 ( n16241,n15360,n15390,n16244 );
   nand U15850 ( n16244,n14899,n14885 );
   nand U15851 ( n15360,n16245,n16246 );
   nand U15852 ( n16246,n16247,n16248,n16249 );
   nand U15853 ( n16249,n15337,n15286,n16250 );
   nand U15854 ( n16250,n15306,n14435 );
   nand U15855 ( n15286,n15281,n14438 );
   nand U15856 ( n15337,n16251,n15285 );
   nand U15857 ( n15285,n14927,n14943 );
   not U15858 ( n16251,n15278 );
   nand U15859 ( n16248,n14941,n14928 );
   nand U15860 ( n16247,n14900,n14915 );
   nand U15861 ( n16245,n15338,n14432 );
   nand U15862 ( n16240,n16252,n14426 );
   nand U15863 ( n16252,n14885,n16243 );
   nand U15864 ( n16236,n14861,n14420 );
   nand U15865 ( n16225,n16227,n16253 );
   nand U15866 ( n16253,n16254,n15676,n16255 );
   nand U15867 ( n16255,n15682,n15678 );
   nand U15868 ( n16212,n14704,n14720 );
   and U15869 ( n15879,n15883,n16211 );
   nand U15870 ( n16190,n14363,n16194,n14610 );
   not U15871 ( n15520,n14986 );
   nand U15872 ( n14986,n16256,n14996 );
   nand U15873 ( n16105,n15293,n14354 );
   nand U15874 ( n15260,n14996,n14579 );
   nand U15875 ( n16104,n14991,n14583 );
   nor U15876 ( n14583,n14992,n16257 );
   and U15877 ( n16257,n16258,n14584 );
   nand U15878 ( n16258,n16259,n16073 );
   not U15879 ( n16259,n16050 );
   nand U15880 ( n16263,p1_reg2_reg_30_,n14995 );
   nand U15881 ( n16261,n14560,n14561,n14991 );
   nand U15882 ( n14560,n14558,n16264 );
   nand U15883 ( n16264,n14992,n14993 );
   nand U15884 ( n16260,n14994,n14558 );
   nand U15885 ( n16267,p1_reg2_reg_31_,n14995 );
   nand U15886 ( n16262,n14559,n14996 );
   nor U15887 ( n14559,n15004,n16268 );
   and U15888 ( n15004,n16269,n16270 );
   nand U15889 ( n16270,n14579,n16271 );
   not U15890 ( n14579,n14596 );
   nand U15891 ( n16269,n16273,n16187 );
   nand U15892 ( n16266,n14991,n14552 );
   xor U15893 ( n14552,n14549,n14561 );
   nand U15894 ( n14561,n16274,n14993,n14992 );
   nor U15895 ( n14992,n14597,n14584,n16050 );
   nand U15896 ( n16050,n14624,n16030,n16053 );
   not U15897 ( n16053,n16001 );
   nand U15898 ( n16001,n14642,n15954,n16005 );
   not U15899 ( n16005,n15930 );
   nand U15900 ( n15930,n14679,n14668,n15916 );
   not U15901 ( n15916,n15871 );
   nand U15902 ( n15871,n14705,n15854,n15874 );
   not U15903 ( n15874,n15823 );
   nand U15904 ( n15823,n15783,n14720,n15827 );
   not U15905 ( n15827,n15770 );
   nand U15906 ( n15770,n15740,n14757,n15773 );
   not U15907 ( n15773,n15691 );
   nand U15908 ( n15691,n15656,n14769,n15695 );
   not U15909 ( n15695,n15637 );
   nand U15910 ( n15637,n14796,n15627,n15593 );
   nor U15911 ( n15627,n14823,n15576 );
   nand U15912 ( n15576,n16275,n14835 );
   not U15913 ( n16275,n15516 );
   nand U15914 ( n15516,n15452,n15490,n15519 );
   not U15915 ( n15519,n15439 );
   nand U15916 ( n15439,n14885,n15411,n15442 );
   not U15917 ( n15442,n15373 );
   nand U15918 ( n15373,n14901,n14915,n15377 );
   not U15919 ( n15377,n15303 );
   nand U15920 ( n15303,n14943,n15261,n14928 );
   nand U15921 ( n15302,n16276,n14996 );
   nand U15922 ( n16265,n14994,n14549 );
   not U15923 ( n14994,n15292 );
   nand U15924 ( n16278,n16279,n16280 );
   nand U15925 ( n16280,n16281,n14962,n16282,n14959 );
   nand U15926 ( n16286,n16287,n16288 );
   nor U15927 ( n16285,n16289,n16290 );
   nor U15928 ( n16290,n16291,n16292,n16293 );
   nor U15929 ( n16293,n16294,n16295,n16296 );
   nor U15930 ( n16295,n16297,n15815 );
   xor U15931 ( n16294,p1_reg2_reg_19_,n16288 );
   nor U15932 ( n16292,n16298,n16299,n16297 );
   nor U15933 ( n16297,n16300,n16301 );
   nor U15934 ( n16299,p1_reg2_reg_18_,n16296 );
   nor U15935 ( n16296,n16302,n16303 );
   not U15936 ( n16302,n16301 );
   xor U15937 ( n16298,n16288,n15836 );
   not U15938 ( n15836,p1_reg2_reg_19_ );
   nor U15939 ( n16289,n16304,n16305,n16306 );
   nor U15940 ( n16306,n16307,n16308,n16309 );
   nor U15941 ( n16308,n16310,n16311 );
   xor U15942 ( n16307,p1_reg1_reg_19_,n16288 );
   nor U15943 ( n16305,n16312,n16313,n16310 );
   nor U15944 ( n16310,n16300,n16314 );
   nor U15945 ( n16313,p1_reg1_reg_18_,n16309 );
   nor U15946 ( n16309,n16315,n16303 );
   xor U15947 ( n16312,n16316,p1_reg1_reg_19_ );
   nand U15948 ( n16284,n16317,p1_addr_reg_19_ );
   nand U15949 ( n16283,p1_reg3_reg_19_,p1_u3086 );
   nand U15950 ( n16322,n16323,n16324,n16325 );
   nand U15951 ( n16325,n16326,n16327 );
   xor U15952 ( n16327,n16301,n15815 );
   not U15953 ( n15815,p1_reg2_reg_18_ );
   nand U15954 ( n16323,n16328,n16329 );
   xor U15955 ( n16329,p1_reg1_reg_18_,n16315 );
   nand U15956 ( n16320,n16330,n16303 );
   nand U15957 ( n16330,n16331,n16332 );
   nand U15958 ( n16332,n16333,n16328 );
   xor U15959 ( n16333,n16315,n16311 );
   not U15960 ( n16311,p1_reg1_reg_18_ );
   not U15961 ( n16315,n16314 );
   nand U15962 ( n16314,n16334,n16335,n16336 );
   or U15963 ( n16336,n16337,n16338 );
   nand U15964 ( n16335,p1_reg1_reg_17_,n16339 );
   or U15965 ( n16339,n16340,n16341 );
   nand U15966 ( n16334,n16341,n16340 );
   nand U15967 ( n16331,n16342,n16326 );
   xor U15968 ( n16342,p1_reg2_reg_18_,n16301 );
   nand U15969 ( n16301,n16343,n16344,n16345 );
   or U15970 ( n16345,n16346,n16347 );
   nand U15971 ( n16344,p1_reg2_reg_17_,n16348 );
   or U15972 ( n16348,n16340,n16349 );
   nand U15973 ( n16343,n16349,n16340 );
   nand U15974 ( n16319,p1_addr_reg_18_,n16317 );
   nand U15975 ( n16318,p1_reg3_reg_18_,p1_u3086 );
   nand U15976 ( n16353,n16287,n16340 );
   nor U15977 ( n16352,n16354,n16355 );
   nor U15978 ( n16355,n16291,n16356,n16357 );
   nor U15979 ( n16357,n16358,n16349,n16359 );
   nor U15980 ( n16359,n16360,n16346 );
   nor U15981 ( n16360,p1_reg2_reg_16_,n16361 );
   xor U15982 ( n16358,n16362,n15799 );
   nor U15983 ( n16356,n16347,n16363,n16364 );
   nor U15984 ( n16364,n15799,n16362 );
   nor U15985 ( n16363,n16349,n16365 );
   not U15986 ( n16365,n16346 );
   nor U15987 ( n16349,n16366,n15769 );
   nand U15988 ( n16347,n16367,n16368 );
   nand U15989 ( n16368,n16366,n15769 );
   nand U15990 ( n16367,n16362,n15799 );
   not U15991 ( n15799,p1_reg2_reg_17_ );
   nor U15992 ( n16354,n16304,n16369,n16370 );
   nor U15993 ( n16370,n16371,n16341,n16372 );
   nor U15994 ( n16372,n16373,n16337 );
   nor U15995 ( n16373,p1_reg1_reg_16_,n16361 );
   xor U15996 ( n16371,n16362,n16374 );
   nor U15997 ( n16369,n16338,n16375,n16376 );
   nor U15998 ( n16376,n16374,n16362 );
   nor U15999 ( n16375,n16341,n16377 );
   not U16000 ( n16377,n16337 );
   nor U16001 ( n16341,n16366,n16378 );
   nand U16002 ( n16338,n16379,n16380 );
   nand U16003 ( n16380,n16366,n16378 );
   nand U16004 ( n16379,n16362,n16374 );
   not U16005 ( n16374,p1_reg1_reg_17_ );
   nand U16006 ( n16351,p1_addr_reg_17_,n16317 );
   nand U16007 ( n16350,p1_reg3_reg_17_,p1_u3086 );
   nand U16008 ( n16385,n16386,n16387 );
   nand U16009 ( n16387,n16328,n16388 );
   xor U16010 ( n16388,n16337,n16378 );
   not U16011 ( n16378,p1_reg1_reg_16_ );
   nand U16012 ( n16386,n16326,n16389 );
   xor U16013 ( n16389,n16346,n15769 );
   not U16014 ( n15769,p1_reg2_reg_16_ );
   nand U16015 ( n16383,n16361,n16390 );
   nand U16016 ( n16390,n16391,n16324,n16392 );
   nand U16017 ( n16392,n16393,n16326 );
   xor U16018 ( n16393,p1_reg2_reg_16_,n16346 );
   nand U16019 ( n16346,n16394,n16395 );
   nand U16020 ( n16395,n16396,n15730 );
   or U16021 ( n16396,n16397,n16398 );
   nand U16022 ( n16394,n16397,n16398 );
   nand U16023 ( n16391,n16399,n16328 );
   xor U16024 ( n16399,p1_reg1_reg_16_,n16337 );
   nand U16025 ( n16337,n16400,n16401 );
   nand U16026 ( n16401,n16402,n16403 );
   or U16027 ( n16402,n16404,n16398 );
   nand U16028 ( n16400,n16404,n16398 );
   nand U16029 ( n16382,p1_addr_reg_16_,n16317 );
   nand U16030 ( n16381,p1_reg3_reg_16_,p1_u3086 );
   nand U16031 ( n16410,n16411,n16324,n16412 );
   nand U16032 ( n16412,n16413,n16326 );
   xor U16033 ( n16413,p1_reg2_reg_15_,n16397 );
   nand U16034 ( n16411,n16414,n16328 );
   xor U16035 ( n16414,p1_reg1_reg_15_,n16404 );
   nand U16036 ( n16407,n16415,n16398 );
   nand U16037 ( n16415,n16416,n16417 );
   nand U16038 ( n16417,n16328,n16418 );
   xor U16039 ( n16418,n16404,n16403 );
   not U16040 ( n16403,p1_reg1_reg_15_ );
   nand U16041 ( n16404,n16419,n16420 );
   nand U16042 ( n16420,n16421,n16422 );
   nand U16043 ( n16421,n16423,n16424 );
   or U16044 ( n16419,n16424,n16423 );
   nand U16045 ( n16416,n16326,n16425 );
   xor U16046 ( n16425,n16397,n15730 );
   not U16047 ( n15730,p1_reg2_reg_15_ );
   nand U16048 ( n16397,n16426,n16427 );
   nand U16049 ( n16427,n16428,n16429 );
   nand U16050 ( n16428,n16430,n16424 );
   or U16051 ( n16426,n16424,n16430 );
   nand U16052 ( n16406,p1_addr_reg_15_,n16317 );
   nand U16053 ( n16405,p1_reg3_reg_15_,p1_u3086 );
   nand U16054 ( n16434,n16435,n16436 );
   nand U16055 ( n16436,n16437,n16438 );
   nand U16056 ( n16438,n16328,n16439 );
   xor U16057 ( n16439,n16423,p1_reg1_reg_14_ );
   nand U16058 ( n16437,n16326,n16440 );
   xor U16059 ( n16440,p1_reg2_reg_14_,n16430 );
   nand U16060 ( n16433,n16424,n16441 );
   nand U16061 ( n16441,n16442,n16324,n16443 );
   nand U16062 ( n16443,n16444,n16326 );
   xor U16063 ( n16444,n16430,n16429 );
   not U16064 ( n16429,p1_reg2_reg_14_ );
   nor U16065 ( n16430,n16445,n16446 );
   and U16066 ( n16445,n16447,n16448,n16449 );
   nand U16067 ( n16449,n16450,p1_reg2_reg_13_ );
   nand U16068 ( n16447,n16451,n16452 );
   nand U16069 ( n16442,n16453,n16328 );
   xor U16070 ( n16453,n16422,n16423 );
   nor U16071 ( n16423,n16454,n16455 );
   and U16072 ( n16454,n16456,n16457,n16458 );
   nand U16073 ( n16458,n16450,p1_reg1_reg_13_ );
   nand U16074 ( n16456,n16459,n16460 );
   not U16075 ( n16422,p1_reg1_reg_14_ );
   nand U16076 ( n16432,p1_addr_reg_14_,n16317 );
   nand U16077 ( n16431,p1_reg3_reg_14_,p1_u3086 );
   nand U16078 ( n16464,n16287,n16450 );
   nor U16079 ( n16463,n16465,n16466 );
   nor U16080 ( n16466,n16291,n16467,n16468 );
   nor U16081 ( n16468,n16469,n16470,n16471 );
   xor U16082 ( n16469,n16472,n15672 );
   nor U16083 ( n16467,n16446,n16473,n16474,n16475 );
   nor U16084 ( n16475,n15672,n16472 );
   not U16085 ( n15672,p1_reg2_reg_13_ );
   nor U16086 ( n16474,n16470,n16451 );
   nor U16087 ( n16446,p1_reg2_reg_13_,n16450 );
   nor U16088 ( n16465,n16304,n16476,n16477 );
   nor U16089 ( n16477,n16478,n16479,n16480 );
   xor U16090 ( n16478,n16450,p1_reg1_reg_13_ );
   nor U16091 ( n16476,n16455,n16481,n16482,n16483 );
   and U16092 ( n16483,p1_reg1_reg_13_,n16450 );
   nor U16093 ( n16482,n16479,n16459 );
   nor U16094 ( n16455,p1_reg1_reg_13_,n16450 );
   nand U16095 ( n16462,p1_addr_reg_13_,n16317 );
   nand U16096 ( n16461,p1_reg3_reg_13_,p1_u3086 );
   nor U16097 ( n16489,n16291,n16471,n16490 );
   nor U16098 ( n16490,n16491,n16451 );
   nor U16099 ( n16491,n16473,n16470 );
   not U16100 ( n16470,n16448 );
   nand U16101 ( n16448,n16492,p1_reg2_reg_12_ );
   nor U16102 ( n16471,n16493,n16473 );
   not U16103 ( n16473,n16452 );
   nand U16104 ( n16452,n16494,n15646 );
   nor U16105 ( n16488,n16304,n16480,n16495 );
   nor U16106 ( n16495,n16496,n16459 );
   nor U16107 ( n16496,n16481,n16479 );
   not U16108 ( n16479,n16457 );
   nand U16109 ( n16457,n16492,p1_reg1_reg_12_ );
   nor U16110 ( n16480,n16497,n16481 );
   not U16111 ( n16481,n16460 );
   nand U16112 ( n16460,n16494,n16498 );
   nor U16113 ( n16487,n16499,n16494 );
   nor U16114 ( n16499,n16500,n16287,n16501 );
   nor U16115 ( n16501,n16304,n16497,n16498 );
   not U16116 ( n16498,p1_reg1_reg_12_ );
   not U16117 ( n16497,n16459 );
   nand U16118 ( n16459,n16502,n16503 );
   nand U16119 ( n16503,n16504,n16505 );
   nand U16120 ( n16505,n16506,n16507 );
   nand U16121 ( n16502,n16508,p1_reg1_reg_11_ );
   nor U16122 ( n16500,n16291,n16493,n15646 );
   not U16123 ( n15646,p1_reg2_reg_12_ );
   not U16124 ( n16493,n16451 );
   nand U16125 ( n16451,n16509,n16510 );
   nand U16126 ( n16510,n16511,n16512 );
   nand U16127 ( n16512,n16506,n15626 );
   nand U16128 ( n16509,n16508,p1_reg2_reg_11_ );
   nand U16129 ( n16485,p1_addr_reg_12_,n16317 );
   nand U16130 ( n16484,p1_reg3_reg_12_,p1_u3086 );
   nand U16131 ( n16517,n16518,n16519 );
   nand U16132 ( n16519,n16328,n16520 );
   xor U16133 ( n16520,n16504,p1_reg1_reg_11_ );
   nand U16134 ( n16518,n16326,n16521 );
   xor U16135 ( n16521,n16511,p1_reg2_reg_11_ );
   nand U16136 ( n16515,n16508,n16522 );
   nand U16137 ( n16522,n16523,n16324,n16524 );
   nand U16138 ( n16524,n16525,n16326 );
   xor U16139 ( n16525,n15626,n16511 );
   nor U16140 ( n16511,n16526,n16527 );
   and U16141 ( n16526,n16528,n16529,n16530 );
   nand U16142 ( n16530,n16531,p1_reg2_reg_10_ );
   nand U16143 ( n16528,n16532,n16533 );
   not U16144 ( n15626,p1_reg2_reg_11_ );
   nand U16145 ( n16523,n16534,n16328 );
   xor U16146 ( n16534,n16507,n16504 );
   nor U16147 ( n16504,n16535,n16536 );
   and U16148 ( n16535,n16537,n16538,n16539 );
   nand U16149 ( n16539,n16531,p1_reg1_reg_10_ );
   nand U16150 ( n16537,n16540,n16541 );
   not U16151 ( n16507,p1_reg1_reg_11_ );
   nand U16152 ( n16514,p1_addr_reg_11_,n16317 );
   nand U16153 ( n16513,p1_reg3_reg_11_,p1_u3086 );
   nand U16154 ( n16545,n16287,n16531 );
   nor U16155 ( n16544,n16546,n16547 );
   nor U16156 ( n16547,n16291,n16548,n16549 );
   nor U16157 ( n16549,n16550,n16551,n16552 );
   nor U16158 ( n16552,n16553,n16554 );
   xor U16159 ( n16550,n16555,n15573 );
   nor U16160 ( n16548,n16527,n16554,n16556,n16557 );
   nor U16161 ( n16557,n15573,n16555 );
   not U16162 ( n15573,p1_reg2_reg_10_ );
   nor U16163 ( n16527,n16531,p1_reg2_reg_10_ );
   nor U16164 ( n16546,n16304,n16558,n16559 );
   nor U16165 ( n16559,n16560,n16561,n16562 );
   nor U16166 ( n16562,n16563,n16564 );
   xor U16167 ( n16560,n16531,p1_reg1_reg_10_ );
   nor U16168 ( n16558,n16536,n16564,n16565,n16566 );
   and U16169 ( n16566,p1_reg1_reg_10_,n16531 );
   nor U16170 ( n16536,n16531,p1_reg1_reg_10_ );
   nand U16171 ( n16543,p1_addr_reg_10_,n16317 );
   nand U16172 ( n16542,p1_reg3_reg_10_,p1_u3086 );
   nor U16173 ( n16572,n16291,n16573,n16574 );
   nor U16174 ( n16574,n16554,n16556 );
   nor U16175 ( n16556,n16551,n16532 );
   not U16176 ( n16551,n16529 );
   nand U16177 ( n16529,n16575,p1_reg2_reg_9_ );
   not U16178 ( n16554,n16533 );
   nor U16179 ( n16573,n16532,n16533 );
   nand U16180 ( n16533,n16576,n15543 );
   nor U16181 ( n16571,n16304,n16577,n16578 );
   nor U16182 ( n16578,n16564,n16565 );
   nor U16183 ( n16565,n16561,n16540 );
   not U16184 ( n16561,n16538 );
   nand U16185 ( n16538,n16575,p1_reg1_reg_9_ );
   not U16186 ( n16564,n16541 );
   nor U16187 ( n16577,n16540,n16541 );
   nand U16188 ( n16541,n16576,n16579 );
   nor U16189 ( n16570,n16580,n16576 );
   nor U16190 ( n16580,n16581,n16287,n16582 );
   nor U16191 ( n16582,n16304,n16563,n16579 );
   not U16192 ( n16579,p1_reg1_reg_9_ );
   not U16193 ( n16563,n16540 );
   nand U16194 ( n16540,n16583,n16584 );
   or U16195 ( n16583,n16585,n16586 );
   nor U16196 ( n16581,n16291,n16553,n15543 );
   not U16197 ( n15543,p1_reg2_reg_9_ );
   not U16198 ( n16553,n16532 );
   nand U16199 ( n16532,n16587,n16588 );
   nand U16200 ( n16587,n16589,n16590 );
   nand U16201 ( n16568,p1_addr_reg_9_,n16317 );
   nand U16202 ( n16567,p1_reg3_reg_9_,p1_u3086 );
   nand U16203 ( n16594,n16287,n16595 );
   nor U16204 ( n16593,n16596,n16597 );
   nor U16205 ( n16597,n16291,n16598 );
   xor U16206 ( n16598,n16599,n16590 );
   nand U16207 ( n16590,n16600,n16601 );
   nand U16208 ( n16601,p1_reg2_reg_7_,n16602 );
   or U16209 ( n16602,n16603,n16604 );
   nand U16210 ( n16600,n16604,n16603 );
   nand U16211 ( n16599,n16589,n16588 );
   nand U16212 ( n16588,n16595,p1_reg2_reg_8_ );
   nand U16213 ( n16589,n16605,n15515 );
   not U16214 ( n15515,p1_reg2_reg_8_ );
   nor U16215 ( n16596,n16304,n16606 );
   xor U16216 ( n16606,n16586,n16607 );
   nor U16217 ( n16607,n16608,n16585 );
   nor U16218 ( n16585,n16595,p1_reg1_reg_8_ );
   not U16219 ( n16608,n16584 );
   nand U16220 ( n16584,n16595,p1_reg1_reg_8_ );
   and U16221 ( n16586,n16609,n16610 );
   nand U16222 ( n16610,p1_reg1_reg_7_,n16611 );
   or U16223 ( n16611,n16612,n16604 );
   nand U16224 ( n16609,n16604,n16612 );
   nand U16225 ( n16592,p1_addr_reg_8_,n16317 );
   nand U16226 ( n16591,p1_reg3_reg_8_,p1_u3086 );
   nor U16227 ( n16618,n16291,n16619,n16620 );
   nor U16228 ( n16620,n16621,n16603 );
   nand U16229 ( n16603,n16622,n16623 );
   nand U16230 ( n16623,n16624,n16625 );
   nor U16231 ( n16621,n16604,n15473 );
   nor U16232 ( n16617,n16304,n16626,n16627 );
   nor U16233 ( n16627,n16628,n16612 );
   nand U16234 ( n16612,n16629,n16630 );
   nand U16235 ( n16630,n16631,n16632 );
   and U16236 ( n16628,n16633,p1_reg1_reg_7_ );
   nor U16237 ( n16616,n16634,n16633 );
   nor U16238 ( n16634,n16635,n16287,n16636 );
   nor U16239 ( n16636,n16304,p1_reg1_reg_7_,n16626 );
   and U16240 ( n16626,n16637,n16632,n16638 );
   xor U16241 ( n16638,n16604,p1_reg1_reg_7_ );
   nand U16242 ( n16637,n16639,n16629 );
   nor U16243 ( n16635,n16291,p1_reg2_reg_7_,n16619 );
   and U16244 ( n16619,n16640,n16625,n16641 );
   xor U16245 ( n16641,n16633,n15473 );
   not U16246 ( n15473,p1_reg2_reg_7_ );
   nand U16247 ( n16640,n16642,n16622 );
   nand U16248 ( n16614,p1_addr_reg_7_,n16317 );
   nand U16249 ( n16613,p1_reg3_reg_7_,p1_u3086 );
   nor U16250 ( n16648,n16291,n16649,n16650 );
   nor U16251 ( n16650,n16651,n16624 );
   and U16252 ( n16651,n16625,n16622 );
   nand U16253 ( n16622,n16652,p1_reg2_reg_6_ );
   and U16254 ( n16649,n16625,n16624 );
   nand U16255 ( n16625,n16653,n15438 );
   nor U16256 ( n16647,n16304,n16654,n16655 );
   nor U16257 ( n16655,n16656,n16631 );
   and U16258 ( n16656,n16632,n16629 );
   nand U16259 ( n16629,n16652,p1_reg1_reg_6_ );
   not U16260 ( n16632,n16657 );
   nor U16261 ( n16654,n16657,n16639 );
   not U16262 ( n16639,n16631 );
   nor U16263 ( n16657,n16652,p1_reg1_reg_6_ );
   nor U16264 ( n16646,n16658,n16653 );
   nor U16265 ( n16658,n16659,n16287,n16660 );
   and U16266 ( n16660,n16328,n16631,p1_reg1_reg_6_ );
   nand U16267 ( n16631,n16661,n16662 );
   nand U16268 ( n16662,p1_reg1_reg_5_,n16663 );
   or U16269 ( n16663,n16664,n16665 );
   nand U16270 ( n16661,n16665,n16664 );
   nor U16271 ( n16659,n16291,n16642,n15438 );
   not U16272 ( n15438,p1_reg2_reg_6_ );
   not U16273 ( n16642,n16624 );
   nand U16274 ( n16624,n16666,n16667 );
   nand U16275 ( n16667,p1_reg2_reg_5_,n16668 );
   or U16276 ( n16668,n16669,n16665 );
   nand U16277 ( n16666,n16665,n16669 );
   nand U16278 ( n16644,p1_addr_reg_6_,n16317 );
   nand U16279 ( n16643,p1_reg3_reg_6_,p1_u3086 );
   nor U16280 ( n16675,n16291,n16676,n16677 );
   nor U16281 ( n16677,n16678,n16669 );
   nand U16282 ( n16669,n16679,n16680 );
   nor U16283 ( n16678,n16665,n15401 );
   nor U16284 ( n16674,n16304,n16681,n16682 );
   nor U16285 ( n16682,n16683,n16664 );
   nand U16286 ( n16664,n16684,n16685 );
   and U16287 ( n16683,n16686,p1_reg1_reg_5_ );
   nor U16288 ( n16673,n16687,n16686 );
   nor U16289 ( n16687,n16688,n16287,n16689 );
   nor U16290 ( n16689,n16291,p1_reg2_reg_5_,n16676 );
   and U16291 ( n16676,n16690,n16691,n16692 );
   xor U16292 ( n16692,n16686,n15401 );
   not U16293 ( n15401,p1_reg2_reg_5_ );
   nand U16294 ( n16690,n16693,n16679 );
   nor U16295 ( n16688,n16304,p1_reg1_reg_5_,n16681 );
   and U16296 ( n16681,n16694,n16695,n16696 );
   xor U16297 ( n16696,n16665,p1_reg1_reg_5_ );
   nand U16298 ( n16694,n16697,n16684 );
   nand U16299 ( n16671,p1_addr_reg_5_,n16317 );
   nand U16300 ( n16670,p1_reg3_reg_5_,p1_u3086 );
   nor U16301 ( n16701,n16702,n16703,n16704 );
   nor U16302 ( n16704,n16705,n16706 );
   nor U16303 ( n16703,n16707,n16708 );
   nor U16304 ( n16707,n16709,n16287,n16710 );
   nor U16305 ( n16710,n16291,n16693,n16711 );
   nor U16306 ( n16709,n16304,n16697,n16712 );
   nor U16307 ( n16702,p1_state_reg,n16713 );
   nand U16308 ( n16700,n16714,n16680,n16326 );
   nand U16309 ( n16680,n16715,n16691 );
   nand U16310 ( n16714,n16693,n16716 );
   nand U16311 ( n16716,n16679,n16691 );
   nand U16312 ( n16691,n16708,n16711 );
   not U16313 ( n16711,p1_reg2_reg_4_ );
   nand U16314 ( n16679,n16717,p1_reg2_reg_4_ );
   not U16315 ( n16693,n16715 );
   nand U16316 ( n16715,n16718,n16719 );
   nand U16317 ( n16719,p1_reg2_reg_3_,n16720 );
   nand U16318 ( n16720,n16721,n16722 );
   or U16319 ( n16718,n16722,n16721 );
   nand U16320 ( n16698,n16723,n16685,n16328 );
   nand U16321 ( n16685,n16724,n16695 );
   nand U16322 ( n16723,n16697,n16725 );
   nand U16323 ( n16725,n16684,n16695 );
   nand U16324 ( n16695,n16708,n16712 );
   not U16325 ( n16712,p1_reg1_reg_4_ );
   nand U16326 ( n16684,n16717,p1_reg1_reg_4_ );
   not U16327 ( n16697,n16724 );
   nand U16328 ( n16724,n16726,n16727 );
   nand U16329 ( n16727,p1_reg1_reg_3_,n16728 );
   nand U16330 ( n16728,n16729,n16722 );
   or U16331 ( n16726,n16722,n16729 );
   nand U16332 ( n16733,n16287,n16734 );
   nor U16333 ( n16732,n16735,n16736 );
   nor U16334 ( n16736,n16737,n16291 );
   xor U16335 ( n16737,n16734,n16738 );
   xor U16336 ( n16738,n16721,p1_reg2_reg_3_ );
   nor U16337 ( n16721,n16739,n16740 );
   and U16338 ( n16740,n16741,n16742 );
   nor U16339 ( n16735,n16743,n16304 );
   xor U16340 ( n16743,n16734,n16744 );
   xor U16341 ( n16744,n16729,p1_reg1_reg_3_ );
   nor U16342 ( n16729,n16745,n16746 );
   nor U16343 ( n16746,n16747,n16748 );
   and U16344 ( n16747,n16749,n16750 );
   nand U16345 ( n16731,p1_addr_reg_3_,n16317 );
   nor U16346 ( n16757,n16304,n16758,n16759 );
   nor U16347 ( n16759,n16760,n16761 );
   xor U16348 ( n16761,n16762,p1_reg1_reg_2_ );
   nor U16349 ( n16758,n16747,n16748,n16745 );
   and U16350 ( n16745,n16762,p1_reg1_reg_2_ );
   nor U16351 ( n16748,n16762,p1_reg1_reg_2_ );
   nand U16352 ( n16760,n16749,n16750 );
   nand U16353 ( n16750,p1_reg1_reg_0_,n16763,p1_ir_reg_0_ );
   not U16354 ( n16756,n16699 );
   nand U16355 ( n16699,n16764,n16765,p1_u3973 );
   nand U16356 ( n16765,n16766,n16767,n16188 );
   or U16357 ( n16767,n16768,n16769 );
   nand U16358 ( n16766,n16768,n16770 );
   nand U16359 ( n16764,n16771,n16772 );
   nand U16360 ( n16771,n16188,n16773 );
   nand U16361 ( n16773,n16774,n16775 );
   nor U16362 ( n16755,n16291,n16776,n16777 );
   nor U16363 ( n16777,n16741,n16778 );
   xor U16364 ( n16778,n16779,n15323 );
   and U16365 ( n16776,n16741,n16742,n16780 );
   not U16366 ( n16780,n16739 );
   nor U16367 ( n16739,n16779,n15323 );
   nand U16368 ( n16742,n16779,n15323 );
   not U16369 ( n15323,p1_reg2_reg_2_ );
   nand U16370 ( n16741,n16781,n16782 );
   nand U16371 ( n16782,n16769,n16783 );
   nand U16372 ( n16753,p1_reg3_reg_2_,p1_u3086 );
   nand U16373 ( n16752,n16287,n16762 );
   nand U16374 ( n16751,p1_addr_reg_2_,n16317 );
   nand U16375 ( n16787,n16287,n16788 );
   not U16376 ( n16287,n16324 );
   nor U16377 ( n16786,n16789,n16790 );
   nor U16378 ( n16790,n16791,n16304 );
   xor U16379 ( n16791,n16792,n16793 );
   nand U16380 ( n16793,n16749,n16763 );
   or U16381 ( n16763,n16788,p1_reg1_reg_1_ );
   nand U16382 ( n16749,n16788,p1_reg1_reg_1_ );
   nor U16383 ( n16792,n16794,n16772 );
   nor U16384 ( n16789,n16795,n16291 );
   xor U16385 ( n16795,n16769,n16796 );
   nand U16386 ( n16796,n16781,n16783 );
   nand U16387 ( n16783,n16797,n15291 );
   not U16388 ( n15291,p1_reg2_reg_1_ );
   nand U16389 ( n16781,n16788,p1_reg2_reg_1_ );
   nor U16390 ( n16769,n16772,n16775 );
   nand U16391 ( n16785,p1_addr_reg_1_,n16317 );
   nand U16392 ( n16784,p1_reg3_reg_1_,p1_u3086 );
   nand U16393 ( n16802,n16803,n16324,n16804 );
   nand U16394 ( n16804,n16326,n16775 );
   not U16395 ( n16775,p1_reg2_reg_0_ );
   nand U16396 ( n16324,n16805,n16272 );
   nand U16397 ( n16803,n16328,n16794 );
   not U16398 ( n16794,p1_reg1_reg_0_ );
   nand U16399 ( n16800,n16806,n16772 );
   nand U16400 ( n16806,n16807,n16808 );
   nand U16401 ( n16808,n16328,p1_reg1_reg_0_ );
   not U16402 ( n16328,n16304 );
   nand U16403 ( n16807,n16326,p1_reg2_reg_0_ );
   not U16404 ( n16326,n16291 );
   and U16405 ( n16805,n16809,n16705 );
   nand U16406 ( n16809,n16810,n16811 );
   nand U16407 ( n16811,n14541,n16812 );
   nand U16408 ( n16812,n16813,n16814,n16815 );
   nor U16409 ( n16815,n16816,n16277,n16114 );
   not U16410 ( n16114,n16279 );
   nand U16411 ( n16810,n16817,p1_state_reg );
   not U16412 ( n16774,n16768 );
   nand U16413 ( n16799,p1_addr_reg_0_,n16317 );
   not U16414 ( n16317,n16705 );
   nand U16415 ( n16705,n16818,n16819 );
   nand U16416 ( n16818,n16820,n16821 );
   nand U16417 ( n16798,p1_reg3_reg_0_,p1_u3086 );
   nor U16418 ( n16824,n16825,n16826,n16827,n16828 );
   and U16419 ( n16828,n14966,n15014,n16829,n16817 );
   nor U16420 ( n16827,n14966,n16829,n16821,n14967 );
   nand U16421 ( n16829,n16830,n16831,n16832,n16833 );
   nor U16422 ( n16833,n16834,n16835 );
   nor U16423 ( n16835,n16836,n16837 );
   nor U16424 ( n16834,n16838,n16839 );
   nor U16425 ( n16839,n16840,n16841 );
   nor U16426 ( n16841,n16842,n16843 );
   nor U16427 ( n16840,n16844,n16845,n16846 );
   not U16428 ( n16845,n16847 );
   not U16429 ( n16838,n16848 );
   nand U16430 ( n16832,n16849,n16850 );
   nand U16431 ( n16850,n16851,n16852 );
   nand U16432 ( n16852,n16853,n16854 );
   nand U16433 ( n16851,n16855,n16856 );
   nand U16434 ( n16831,n16857,n16858,n16859,n16860 );
   nand U16435 ( n16860,n16861,n16862 );
   nand U16436 ( n16862,n16863,n16864 );
   nand U16437 ( n16861,n16865,n16866 );
   nand U16438 ( n16866,n16867,n16868 );
   nand U16439 ( n16868,n16869,n16870 );
   nand U16440 ( n16867,n16871,n16872 );
   nand U16441 ( n16872,n16873,n16874,n16875 );
   nand U16442 ( n16875,n16876,n16877 );
   nand U16443 ( n16874,n16878,n16879 );
   or U16444 ( n16879,n16877,n16876 );
   and U16445 ( n16876,n16880,n16881 );
   nand U16446 ( n16881,n16882,n16883 );
   nand U16447 ( n16880,n14378,n16884 );
   nand U16448 ( n16877,n16885,n16886 );
   nand U16449 ( n16886,n16887,n16888 );
   nand U16450 ( n16888,n15854,n16889 );
   not U16451 ( n16887,n16890 );
   nand U16452 ( n16885,n16891,n16892 );
   nand U16453 ( n16892,n16889,n16890,n16893 );
   nand U16454 ( n16893,n14693,n16884 );
   nand U16455 ( n16890,n16894,n16895 );
   nand U16456 ( n16895,n14381,n16884 );
   nand U16457 ( n16894,n14693,n16883 );
   nand U16458 ( n16889,n14381,n16883 );
   nand U16459 ( n16891,n16896,n16897 );
   nand U16460 ( n16897,n16898,n16899,n16900,n16901 );
   nand U16461 ( n16901,n16902,n16903 );
   nor U16462 ( n16900,n16904,n16905 );
   nor U16463 ( n16905,n16906,n16907 );
   nor U16464 ( n16904,n16908,n16909,n16910 );
   not U16465 ( n16909,n16911 );
   nand U16466 ( n16899,n16912,n16913,n16914 );
   nand U16467 ( n16898,n16914,n16915,n16916,n16917 );
   nand U16468 ( n16917,n16918,n16919 );
   nand U16469 ( n16919,n16920,n16921 );
   nand U16470 ( n16918,n16922,n16923 );
   nand U16471 ( n16923,n16924,n16925 );
   nand U16472 ( n16925,n16926,n16927 );
   nand U16473 ( n16924,n16928,n16929 );
   nand U16474 ( n16929,n16930,n16931 );
   nand U16475 ( n16928,n16932,n16933,n16934,n16935 );
   nand U16476 ( n16935,n16936,n16937,n16938 );
   nand U16477 ( n16934,n16939,n16936,n16940 );
   nand U16478 ( n16940,n16941,n16942 );
   nand U16479 ( n16942,n16943,n16944,n16945 );
   nor U16480 ( n16945,n16946,n16947,n16948 );
   nor U16481 ( n16948,n16949,n16950 );
   nor U16482 ( n16947,n16951,n16952,n16953 );
   not U16483 ( n16952,n16954 );
   nor U16484 ( n16946,n16955,n16956,n16957 );
   nand U16485 ( n16944,n16958,n16959,n16960,n16961 );
   nand U16486 ( n16961,n16962,n16963,n16964,n16965 );
   or U16487 ( n16965,n16966,n16967 );
   nand U16488 ( n16964,n16968,n16969 );
   nand U16489 ( n16963,n16970,n16971,n16972,n16973 );
   and U16490 ( n16973,n16974,n16975,n16976 );
   xor U16491 ( n16972,n15287,n16883 );
   nand U16492 ( n16971,n16977,n16978 );
   nand U16493 ( n16962,n16979,n16970 );
   nand U16494 ( n16970,n16967,n16966 );
   nand U16495 ( n16966,n16980,n16981 );
   nand U16496 ( n16981,n15392,n16883 );
   nand U16497 ( n16980,n14426,n16884 );
   and U16498 ( n16967,n16982,n16983 );
   nand U16499 ( n16983,n15392,n16884 );
   nand U16500 ( n16982,n14426,n16883 );
   nand U16501 ( n16979,n16984,n16985 );
   nand U16502 ( n16985,n16986,n16974 );
   nand U16503 ( n16974,n16987,n16988 );
   nand U16504 ( n16986,n16989,n16990 );
   nand U16505 ( n16990,n16991,n16976 );
   nand U16506 ( n16976,n16992,n16993 );
   nand U16507 ( n16991,n16994,n16995 );
   or U16508 ( n16995,n16977,n16996,n16978 );
   nand U16509 ( n16978,n16997,n16998 );
   nand U16510 ( n16998,n15281,n16883 );
   nand U16511 ( n16997,n14438,n16884 );
   not U16512 ( n16996,n16975 );
   nand U16513 ( n16975,n16999,n17000 );
   and U16514 ( n16977,n17001,n17002 );
   nand U16515 ( n17002,n14438,n16883 );
   nand U16516 ( n17001,n15281,n16884 );
   or U16517 ( n16994,n17000,n16999 );
   and U16518 ( n16999,n17003,n17004 );
   nand U16519 ( n17004,n14435,n16883 );
   nand U16520 ( n17003,n15306,n16884 );
   nand U16521 ( n17000,n17005,n17006 );
   nand U16522 ( n17006,n15306,n16883 );
   nand U16523 ( n17005,n14435,n16884 );
   or U16524 ( n16989,n16993,n16992 );
   and U16525 ( n16992,n17007,n17008 );
   nand U16526 ( n17008,n14432,n16883 );
   nand U16527 ( n17007,n15338,n16884 );
   nand U16528 ( n16993,n17009,n17010 );
   nand U16529 ( n17010,n15338,n16883 );
   nand U16530 ( n17009,n14432,n16884 );
   or U16531 ( n16984,n16988,n16987 );
   and U16532 ( n16987,n17011,n17012 );
   nand U16533 ( n17012,n15376,n16884 );
   nand U16534 ( n17011,n14429,n16883 );
   nand U16535 ( n16988,n17013,n17014 );
   nand U16536 ( n17014,n15376,n16883 );
   nand U16537 ( n17013,n14429,n16884 );
   or U16538 ( n16960,n16969,n16968 );
   and U16539 ( n16968,n17015,n17016 );
   nand U16540 ( n17016,n14873,n16883 );
   nand U16541 ( n17015,n14423,n16884 );
   nand U16542 ( n16969,n17017,n17018 );
   nand U16543 ( n17018,n14873,n16884 );
   nand U16544 ( n17017,n14423,n16883 );
   nand U16545 ( n16959,n16956,n16957 );
   nand U16546 ( n16957,n17019,n17020 );
   nand U16547 ( n17020,n14861,n16883 );
   nand U16548 ( n17019,n14420,n16884 );
   and U16549 ( n16956,n17021,n17022 );
   nand U16550 ( n17022,n14420,n16883 );
   nand U16551 ( n17021,n14861,n16884 );
   not U16552 ( n16958,n16955 );
   nand U16553 ( n16955,n17023,n16954 );
   nand U16554 ( n16954,n16949,n16950 );
   nand U16555 ( n16950,n17024,n17025 );
   nand U16556 ( n17025,n15532,n16883 );
   nand U16557 ( n17024,n14414,n16884 );
   and U16558 ( n16949,n17026,n17027 );
   nand U16559 ( n17027,n14414,n16883 );
   nand U16560 ( n17026,n15532,n16884 );
   nand U16561 ( n17023,n16953,n16951 );
   nand U16562 ( n16951,n17028,n17029 );
   nand U16563 ( n17029,n14417,n16884 );
   nand U16564 ( n17028,n14850,n16883 );
   and U16565 ( n16953,n17030,n17031 );
   nand U16566 ( n17031,n14850,n16884 );
   nand U16567 ( n17030,n14417,n16883 );
   nand U16568 ( n16943,n17032,n17033 );
   or U16569 ( n16941,n17033,n17032 );
   and U16570 ( n17032,n17034,n17035 );
   nand U16571 ( n17035,n14823,n16883 );
   nand U16572 ( n17034,n14411,n16884 );
   nand U16573 ( n17033,n17036,n17037 );
   nand U16574 ( n17037,n14411,n16883 );
   nand U16575 ( n17036,n14823,n16884 );
   nand U16576 ( n16936,n17038,n17039 );
   or U16577 ( n16939,n16937,n16938 );
   and U16578 ( n16938,n17040,n17041 );
   nand U16579 ( n17041,n14408,n16883 );
   nand U16580 ( n17040,n14812,n16884 );
   nand U16581 ( n16937,n17042,n17043 );
   nand U16582 ( n17043,n14812,n16883 );
   nand U16583 ( n17042,n14408,n16884 );
   or U16584 ( n16933,n17039,n17038 );
   and U16585 ( n17038,n17044,n17045 );
   nand U16586 ( n17045,n15640,n16883 );
   nand U16587 ( n17044,n14405,n16884 );
   nand U16588 ( n17039,n17046,n17047 );
   nand U16589 ( n17047,n15640,n16884 );
   nand U16590 ( n17046,n14405,n16883 );
   or U16591 ( n16932,n16931,n16930 );
   and U16592 ( n16930,n17048,n17049 );
   nand U16593 ( n17049,n14784,n16883 );
   nand U16594 ( n17048,n14402,n16884 );
   nand U16595 ( n16931,n17050,n17051 );
   nand U16596 ( n17051,n14402,n16883 );
   nand U16597 ( n17050,n14784,n16884 );
   or U16598 ( n16922,n16927,n16926 );
   and U16599 ( n16926,n17052,n17053 );
   nand U16600 ( n17053,n15694,n16884 );
   nand U16601 ( n17052,n14399,n16883 );
   nand U16602 ( n16927,n17054,n17055 );
   nand U16603 ( n17055,n15694,n16883 );
   nand U16604 ( n17054,n14399,n16884 );
   or U16605 ( n16916,n16921,n16920 );
   and U16606 ( n16920,n17056,n17057 );
   nand U16607 ( n17057,n15722,n16884 );
   nand U16608 ( n17056,n14396,n16883 );
   nand U16609 ( n16921,n17058,n17059 );
   nand U16610 ( n17059,n14396,n16884 );
   nand U16611 ( n17058,n15722,n16883 );
   or U16612 ( n16915,n16913,n16912 );
   and U16613 ( n16912,n17060,n17061 );
   nand U16614 ( n17061,n14745,n16884 );
   nand U16615 ( n17060,n14393,n16883 );
   nand U16616 ( n16913,n17062,n17063 );
   nand U16617 ( n17063,n14745,n16883 );
   nand U16618 ( n17062,n14393,n16884 );
   and U16619 ( n16914,n17064,n16911 );
   nand U16620 ( n16911,n16906,n16907 );
   nand U16621 ( n16907,n17065,n17066 );
   nand U16622 ( n17066,n14387,n16883 );
   nand U16623 ( n17065,n15826,n16884 );
   and U16624 ( n16906,n17067,n17068 );
   nand U16625 ( n17068,n15826,n16883 );
   nand U16626 ( n17067,n14387,n16884 );
   nand U16627 ( n17064,n16910,n16908 );
   nand U16628 ( n16908,n17069,n17070 );
   nand U16629 ( n17070,n14734,n16884 );
   nand U16630 ( n17069,n14390,n16883 );
   and U16631 ( n16910,n17071,n17072 );
   nand U16632 ( n17072,n14734,n16883 );
   nand U16633 ( n17071,n14390,n16884 );
   or U16634 ( n16896,n16903,n16902 );
   and U16635 ( n16902,n17073,n17074 );
   nand U16636 ( n17074,n14384,n16883 );
   nand U16637 ( n17073,n15840,n16884 );
   nand U16638 ( n16903,n17075,n17076 );
   nand U16639 ( n17076,n14384,n16884 );
   nand U16640 ( n17075,n15840,n16883 );
   nand U16641 ( n16878,n17077,n17078 );
   nand U16642 ( n17078,n14378,n16883 );
   nand U16643 ( n17077,n16882,n16884 );
   nand U16644 ( n16873,n17079,n17080 );
   or U16645 ( n16871,n17080,n17079 );
   and U16646 ( n17079,n17081,n17082 );
   nand U16647 ( n17082,n15933,n16883 );
   nand U16648 ( n17081,n14375,n16884 );
   nand U16649 ( n17080,n17083,n17084 );
   nand U16650 ( n17084,n15933,n16884 );
   nand U16651 ( n17083,n14375,n16883 );
   or U16652 ( n16865,n16870,n16869 );
   and U16653 ( n16869,n17085,n17086 );
   nand U16654 ( n17086,n14657,n16883 );
   nand U16655 ( n17085,n14372,n16884 );
   nand U16656 ( n16870,n17087,n17088 );
   nand U16657 ( n17088,n14372,n16883 );
   nand U16658 ( n17087,n14657,n16884 );
   or U16659 ( n16859,n16864,n16863 );
   and U16660 ( n16863,n17089,n17090 );
   nand U16661 ( n17090,n16004,n16883 );
   nand U16662 ( n17089,n14369,n16884 );
   nand U16663 ( n16864,n17091,n17092 );
   nand U16664 ( n17092,n14369,n16883 );
   nand U16665 ( n17091,n16004,n16884 );
   nand U16666 ( n16858,n17093,n17094 );
   nand U16667 ( n16830,n16857,n17095 );
   nand U16668 ( n17095,n17096,n17097 );
   or U16669 ( n17097,n17094,n17093 );
   and U16670 ( n17093,n17098,n17099 );
   nand U16671 ( n17099,n16017,n16884 );
   nand U16672 ( n17098,n14366,n16883 );
   nand U16673 ( n17094,n17100,n17101 );
   nand U16674 ( n17101,n16017,n16883 );
   nand U16675 ( n17100,n14366,n16884 );
   nand U16676 ( n17096,n17102,n17103,n17104 );
   nand U16677 ( n17103,n14363,n16884 );
   nand U16678 ( n17102,n14610,n16883 );
   and U16679 ( n16857,n17105,n17106,n16849 );
   and U16680 ( n16849,n17107,n17108,n16847,n16848 );
   nand U16681 ( n16848,n16836,n16837 );
   nand U16682 ( n16837,n17109,n17110 );
   nand U16683 ( n17110,n14348,n16883 );
   nand U16684 ( n17109,n14549,n16884 );
   and U16685 ( n16836,n17111,n17112 );
   nand U16686 ( n17112,n14549,n16883 );
   nand U16687 ( n17111,n14348,n16884 );
   nand U16688 ( n16847,n16842,n16843 );
   nand U16689 ( n16843,n17113,n17114 );
   nand U16690 ( n17114,n17115,n16884 );
   nand U16691 ( n17113,n14558,n16883 );
   and U16692 ( n16842,n17116,n17117 );
   nand U16693 ( n17117,n17115,n16883 );
   nand U16694 ( n17116,n14558,n16884 );
   or U16695 ( n17108,n16854,n16853 );
   and U16696 ( n16853,n17118,n17119 );
   nand U16697 ( n17119,n14357,n16884 );
   nand U16698 ( n17118,n14584,n16883 );
   nand U16699 ( n16854,n17120,n17121 );
   nand U16700 ( n17121,n14584,n16884 );
   nand U16701 ( n17120,n14357,n16883 );
   nand U16702 ( n17107,n16846,n16844 );
   nand U16703 ( n16844,n17122,n17123 );
   nand U16704 ( n17123,n14571,n16883 );
   nand U16705 ( n17122,n14354,n16884 );
   and U16706 ( n16846,n17124,n17125 );
   nand U16707 ( n17125,n14354,n16883 );
   nand U16708 ( n17124,n14571,n16884 );
   nand U16709 ( n17106,n17126,n17127,n17128 );
   not U16710 ( n17128,n17104 );
   nand U16711 ( n17104,n17129,n17130 );
   nand U16712 ( n17130,n14610,n16884 );
   nand U16713 ( n17129,n14363,n16883 );
   nand U16714 ( n17127,n14620,n16884 );
   nand U16715 ( n17126,n16030,n16883 );
   or U16716 ( n17105,n16856,n16855 );
   and U16717 ( n16855,n17131,n17132 );
   nand U16718 ( n17132,n14597,n16883 );
   nand U16719 ( n17131,n14360,n16884 );
   nand U16720 ( n16856,n17133,n17134 );
   nand U16721 ( n17134,n14597,n16884 );
   nand U16722 ( n17133,n14360,n16883 );
   nor U16723 ( n16826,n17135,n17136,n17137 );
   nor U16724 ( n17137,n17138,n16316 );
   and U16725 ( n17138,n17139,n16817 );
   nor U16726 ( n17136,n16288,n17140 );
   nor U16727 ( n17140,n16821,n17139 );
   nand U16728 ( n17139,n17141,n17142,n17143,n17144 );
   nor U16729 ( n17144,n17145,n17146,n17147,n17148 );
   or U16730 ( n17148,n15310,n15288,n15332,n17149 );
   xor U16731 ( n15332,n14432,n15338 );
   nand U16732 ( n15288,n17150,n17151 );
   xor U16733 ( n15310,n14435,n15306 );
   or U16734 ( n17147,n15387,n15471,n15697,n15721 );
   xor U16735 ( n15721,n14396,n15722 );
   xor U16736 ( n15697,n14399,n15694 );
   not U16737 ( n15471,n15478 );
   xor U16738 ( n15478,n14872,n14861 );
   xor U16739 ( n15387,n14426,n15392 );
   nand U16740 ( n17146,n15944,n15971,n16126,n15021 );
   not U16741 ( n15021,n14987 );
   nand U16742 ( n14987,n17152,n17153 );
   xor U16743 ( n16126,n14357,n16112 );
   xor U16744 ( n15971,n14641,n14657 );
   xor U16745 ( n15944,n15975,n15933 );
   nand U16746 ( n17145,n17154,n15263,n15359,n15434 );
   nand U16747 ( n15434,n15480,n15477 );
   nand U16748 ( n15477,n14873,n14423 );
   nand U16749 ( n15480,n14883,n15411 );
   nand U16750 ( n15359,n16243,n15390 );
   nand U16751 ( n15390,n14884,n14901 );
   nand U16752 ( n16243,n15376,n14429 );
   nand U16753 ( n15263,n15278,n17155 );
   nand U16754 ( n17155,n14942,n15261 );
   nand U16755 ( n15278,n14956,n14441 );
   nor U16756 ( n17143,n17156,n17157,n15842,n17158 );
   not U16757 ( n17158,n17159 );
   and U16758 ( n15842,n15883,n15881 );
   nand U16759 ( n15881,n15840,n14384 );
   nand U16760 ( n15883,n14718,n14705 );
   nand U16761 ( n17157,n15530,n15641,n15752 );
   nand U16762 ( n15752,n15806,n15803 );
   nand U16763 ( n15803,n14745,n14393 );
   nand U16764 ( n15806,n14755,n15740 );
   nand U16765 ( n15641,n15676,n15678 );
   nand U16766 ( n15678,n14811,n14796 );
   nand U16767 ( n15676,n14405,n15640 );
   nand U16768 ( n15530,n15580,n15583 );
   nand U16769 ( n15583,n14849,n14835 );
   nand U16770 ( n15580,n14414,n15532 );
   nand U16771 ( n17156,n15999,n16018,n16058,n16086 );
   nand U16772 ( n16086,n16193,n16194 );
   nand U16773 ( n16194,n14609,n16073 );
   nand U16774 ( n16193,n14360,n14597 );
   nand U16775 ( n16058,n16102,n16101 );
   nand U16776 ( n16101,n14610,n14363 );
   nand U16777 ( n16102,n14620,n16030 );
   nand U16778 ( n16018,n16057,n16060 );
   nand U16779 ( n16060,n14640,n14624 );
   nand U16780 ( n16057,n16017,n14366 );
   nand U16781 ( n15999,n16062,n16064 );
   nand U16782 ( n16064,n16004,n14369 );
   nand U16783 ( n16062,n14621,n14642 );
   nor U16784 ( n17142,n15913,n17160,n15820,n15796 );
   not U16785 ( n15796,n15804 );
   nand U16786 ( n15804,n16216,n16213 );
   nand U16787 ( n16213,n14734,n14390 );
   nand U16788 ( n16216,n14719,n15783 );
   nor U16789 ( n15820,n15920,n17161 );
   nor U16790 ( n17161,n14387,n15826 );
   nor U16791 ( n15920,n14704,n14720 );
   not U16792 ( n17160,n15867 );
   nand U16793 ( n15867,n15878,n16211 );
   nand U16794 ( n16211,n14703,n15854 );
   nand U16795 ( n15878,n14693,n14381 );
   not U16796 ( n15913,n15906 );
   nand U16797 ( n15906,n16204,n16206 );
   nand U16798 ( n16206,n14667,n14679 );
   nand U16799 ( n16204,n14378,n16882 );
   nor U16800 ( n17141,n15670,n15622,n15571,n15502 );
   not U16801 ( n15502,n15507 );
   nand U16802 ( n15507,n16234,n16235 );
   nand U16803 ( n16235,n14834,n15490 );
   nand U16804 ( n16234,n14850,n14417 );
   not U16805 ( n15571,n15581 );
   nand U16806 ( n15581,n16232,n16229 );
   nand U16807 ( n16229,n14823,n14411 );
   nand U16808 ( n16232,n14833,n15553 );
   nor U16809 ( n15622,n15682,n17162 );
   nor U16810 ( n17162,n14408,n14812 );
   nor U16811 ( n15682,n15593,n14795 );
   not U16812 ( n15670,n15677 );
   nand U16813 ( n15677,n16254,n16227 );
   nand U16814 ( n16227,n14794,n15656 );
   nand U16815 ( n16254,n14402,n14784 );
   nand U16816 ( n16825,n17163,n17164,n17165 );
   nand U16817 ( n17165,n17166,n17154,n16817,n17167 );
   nor U16818 ( n17167,n17168,n16288 );
   nand U16819 ( n17166,n17169,n17170 );
   nand U16820 ( n17170,n17171,n17172,n17173 );
   or U16821 ( n17173,n17152,n14348 );
   nand U16822 ( n17172,n17174,n17153,n17175,n17176 );
   nand U16823 ( n17176,n17177,n15017,n16129 );
   nand U16824 ( n17177,n17178,n16130 );
   nand U16825 ( n17178,n16046,n17179 );
   nand U16826 ( n17179,n17180,n17181 );
   nand U16827 ( n17181,n17182,n17183,n17184 );
   nand U16828 ( n17182,n16134,n15941,n15984,n17185 );
   nor U16829 ( n17185,n17186,n17187 );
   nor U16830 ( n17187,n15970,n17188 );
   nor U16831 ( n17188,n17189,n17190,n15904 );
   not U16832 ( n15904,n15914 );
   nor U16833 ( n17189,n17191,n17192 );
   nor U16834 ( n17191,n17193,n17194,n15766 );
   not U16835 ( n15766,n16157 );
   nor U16836 ( n17186,n17192,n15970,n17195 );
   nor U16837 ( n17195,n17196,n17197 );
   nor U16838 ( n17197,n17198,n15767 );
   nor U16839 ( n17198,n14755,n14745 );
   nor U16840 ( n17196,n17199,n15765 );
   nand U16841 ( n15765,n15728,n17200 );
   nand U16842 ( n17200,n15740,n14393 );
   not U16843 ( n15740,n14745 );
   nor U16844 ( n17199,n15710,n17201 );
   nor U16845 ( n17201,n17202,n15711,n17203 );
   nor U16846 ( n17203,n16163,n17204 );
   nor U16847 ( n17204,n17205,n17206 );
   nor U16848 ( n17205,n17207,n17208,n17209,n16172 );
   nor U16849 ( n17209,n17210,n15621 );
   nor U16850 ( n17210,n17211,n17212 );
   nor U16851 ( n17211,n17213,n17214 );
   nor U16852 ( n17213,n16176,n17215 );
   nor U16853 ( n17215,n17216,n17217 );
   not U16854 ( n17217,n16178 );
   nor U16855 ( n17216,n17218,n15436,n15430 );
   nor U16856 ( n17218,n17219,n17220 );
   nor U16857 ( n17208,n17221,n17214,n15349 );
   nand U16858 ( n15349,n17222,n15313 );
   not U16859 ( n17222,n15321 );
   nor U16860 ( n15321,n15322,n17223 );
   nand U16861 ( n15322,n17150,n17224 );
   nand U16862 ( n17224,n15287,n17151 );
   not U16863 ( n15287,n15267 );
   nand U16864 ( n17221,n17225,n15569,n17226 );
   not U16865 ( n17207,n16166 );
   nand U16866 ( n17153,n17227,n14571 );
   nand U16867 ( n17171,n17228,n14549 );
   nand U16868 ( n17228,n17152,n17159 );
   or U16869 ( n17169,n16274,n17115 );
   nor U16870 ( n17115,n15003,n16268 );
   and U16871 ( n16823,n14970,n17164,n17163 );
   nand U16872 ( n17163,n17229,n16817,n14970 );
   xor U16873 ( n17229,n16316,n17230 );
   nand U16874 ( n17230,n17154,n17231,n17232 );
   nand U16875 ( n17232,n17233,n16142,n17234,n17235 );
   nor U16876 ( n17235,n17236,n17190,n17237,n17238 );
   nor U16877 ( n17238,n17239,n17192 );
   nand U16878 ( n17192,n16145,n15915,n17240 );
   nand U16879 ( n17240,n17241,n16146 );
   nand U16880 ( n17241,n16151,n17242,n16148 );
   nand U16881 ( n16148,n14705,n14384 );
   nand U16882 ( n17242,n16154,n16149 );
   nor U16883 ( n16154,n14734,n14719 );
   nand U16884 ( n16151,n14720,n14387 );
   not U16885 ( n14720,n15826 );
   nand U16886 ( n16145,n15854,n14381 );
   nor U16887 ( n17239,n17194,n17243 );
   nor U16888 ( n17243,n17244,n17245 );
   nor U16889 ( n17245,n17193,n17246,n16162 );
   nand U16890 ( n16162,n15767,n16157 );
   nand U16891 ( n16157,n14755,n14745 );
   nand U16892 ( n15767,n14770,n15722 );
   nor U16893 ( n17246,n15768,n17247 );
   nor U16894 ( n17247,n17248,n15710 );
   nor U16895 ( n15710,n14399,n14769 );
   nor U16896 ( n17248,n15711,n17249 );
   nor U16897 ( n17249,n17250,n16163 );
   nor U16898 ( n16163,n14402,n15656 );
   nor U16899 ( n17250,n17251,n17252,n17202,n17206 );
   nand U16900 ( n17206,n16168,n17253 );
   nand U16901 ( n17253,n16166,n14408,n15593 );
   nand U16902 ( n16168,n14796,n14405 );
   not U16903 ( n14796,n15640 );
   nor U16904 ( n17202,n14794,n14784 );
   and U16905 ( n17252,n15621,n16166,n15625 );
   not U16906 ( n15621,n15569 );
   nand U16907 ( n15569,n15553,n14411 );
   not U16908 ( n15553,n14823 );
   nor U16909 ( n17251,n17254,n16172,n17212 );
   nand U16910 ( n17212,n15539,n17255 );
   nand U16911 ( n17255,n14850,n15540,n14834 );
   nand U16912 ( n15539,n14849,n15532 );
   not U16913 ( n14849,n14414 );
   nand U16914 ( n16172,n15568,n15625 );
   nand U16915 ( n15625,n14795,n14812 );
   nand U16916 ( n15568,n14833,n14823 );
   nand U16917 ( n17254,n17256,n16166,n17257 );
   nand U16918 ( n17257,n16173,n15540,n16176 );
   nor U16919 ( n16176,n14420,n15452 );
   nand U16920 ( n16166,n14811,n15640 );
   not U16921 ( n14811,n14405 );
   nand U16922 ( n17256,n17225,n17258,n17259 );
   not U16923 ( n17259,n17214 );
   nand U16924 ( n17214,n15540,n15470,n16173 );
   nand U16925 ( n16173,n15490,n14417 );
   not U16926 ( n15490,n14850 );
   nand U16927 ( n15470,n15452,n14420 );
   not U16928 ( n15452,n14861 );
   nand U16929 ( n15540,n14835,n14414 );
   not U16930 ( n14835,n15532 );
   nand U16931 ( n17258,n17220,n17260,n17261,n17262 );
   nand U16932 ( n17262,n17226,n17151,n17263,n15313 );
   nand U16933 ( n15313,n14928,n14435 );
   nand U16934 ( n17263,n17150,n15267,n17264 );
   nand U16935 ( n17264,n17135,n15268 );
   nand U16936 ( n15268,n15261,n14441 );
   not U16937 ( n15261,n14956 );
   nand U16938 ( n15267,n14942,n14956 );
   not U16939 ( n14942,n14441 );
   nand U16940 ( n17150,n14927,n15281 );
   not U16941 ( n14927,n14438 );
   nand U16942 ( n17151,n14943,n14438 );
   nor U16943 ( n17261,n15436,n15430 );
   not U16944 ( n15430,n15395 );
   nand U16945 ( n15395,n14899,n15392 );
   nand U16946 ( n17260,n17223,n17226 );
   and U16947 ( n17226,n15369,n17265 );
   nand U16948 ( n17265,n14915,n14432 );
   not U16949 ( n17223,n15312 );
   nand U16950 ( n15312,n14941,n15306 );
   not U16951 ( n14941,n14435 );
   and U16952 ( n17220,n15370,n17266 );
   nand U16953 ( n17266,n15338,n15369,n14900 );
   not U16954 ( n14900,n14432 );
   nand U16955 ( n15369,n14901,n14429 );
   nand U16956 ( n15370,n14884,n15376 );
   and U16957 ( n17225,n16178,n17267 );
   nand U16958 ( n17267,n17219,n16177 );
   not U16959 ( n16177,n15436 );
   nor U16960 ( n15436,n14423,n15411 );
   not U16961 ( n17219,n15396 );
   nand U16962 ( n15396,n14885,n14426 );
   not U16963 ( n14885,n15392 );
   nand U16964 ( n16178,n15411,n14423 );
   not U16965 ( n15411,n14873 );
   not U16966 ( n15711,n15706 );
   nand U16967 ( n15706,n14769,n14399 );
   not U16968 ( n14769,n15694 );
   not U16969 ( n15768,n15728 );
   nand U16970 ( n15728,n14757,n14396 );
   not U16971 ( n14757,n15722 );
   nor U16972 ( n17244,n17193,n14755,n14745 );
   nand U16973 ( n17193,n16149,n16152 );
   nand U16974 ( n16152,n14719,n14734 );
   nand U16975 ( n16149,n14704,n15826 );
   not U16976 ( n14704,n14387 );
   not U16977 ( n17194,n16146 );
   nand U16978 ( n16146,n14718,n15840 );
   not U16979 ( n17237,n17268 );
   nor U16980 ( n17190,n15854,n15903,n14381 );
   not U16981 ( n15903,n15915 );
   nand U16982 ( n15915,n14679,n14378 );
   not U16983 ( n15854,n14693 );
   not U16984 ( n17236,n16134 );
   and U16985 ( n16142,n15914,n15941,n15984 );
   nand U16986 ( n15941,n15975,n15933 );
   not U16987 ( n15975,n14375 );
   nand U16988 ( n15914,n14667,n16882 );
   nand U16989 ( n17231,n17269,n17268,n17234 );
   not U16990 ( n17234,n17149 );
   nand U16991 ( n17149,n17270,n17175 );
   nand U16992 ( n17175,n17271,n14348 );
   not U16993 ( n17271,n14549 );
   nand U16994 ( n17270,n15003,n14558 );
   not U16995 ( n15003,n14351 );
   nand U16996 ( n17268,n14571,n17159,n17227 );
   not U16997 ( n17227,n14354 );
   nand U16998 ( n17269,n17152,n17159,n17272 );
   nand U16999 ( n17272,n17233,n17273 );
   nand U17000 ( n17273,n17184,n17274,n17183,n17275 );
   nand U17001 ( n17275,n15984,n16134,n15970 );
   not U17002 ( n15970,n15940 );
   nand U17003 ( n15940,n14668,n14375 );
   not U17004 ( n14668,n15933 );
   nand U17005 ( n15984,n14641,n14657 );
   nand U17006 ( n17183,n14372,n16134,n15954 );
   nand U17007 ( n16134,n14621,n16004 );
   and U17008 ( n17184,n17276,n16136 );
   nand U17009 ( n16136,n14642,n14369 );
   nand U17010 ( n17276,n14624,n14366 );
   and U17011 ( n17233,n17174,n17277 );
   nand U17012 ( n17277,n17274,n17278 );
   nand U17013 ( n17278,n16130,n17180 );
   nand U17014 ( n17180,n14640,n16017 );
   nand U17015 ( n16130,n14620,n14610 );
   and U17016 ( n17274,n16046,n15017,n16129 );
   nand U17017 ( n16129,n16073,n14360 );
   nand U17018 ( n16046,n16030,n14363 );
   and U17019 ( n17174,n15011,n17279 );
   nand U17020 ( n17279,n17280,n15017 );
   nand U17021 ( n15017,n16112,n14357 );
   not U17022 ( n16112,n14584 );
   not U17023 ( n17280,n16128 );
   nand U17024 ( n16128,n14609,n14597 );
   nand U17025 ( n15011,n14595,n14584 );
   not U17026 ( n14595,n14357 );
   nand U17027 ( n17159,n16274,n14351 );
   nand U17028 ( n14351,n17281,n17282,n17283 );
   nand U17029 ( n17283,p1_reg2_reg_30_,n17284 );
   nand U17030 ( n17282,p1_reg0_reg_30_,n17285 );
   nand U17031 ( n17281,p1_reg1_reg_30_,n17286 );
   not U17032 ( n16274,n14558 );
   nand U17033 ( n14558,n17287,n17288 );
   nand U17034 ( n17288,n17289,n11804 );
   xor U17035 ( n11804,n17290,n17291 );
   nand U17036 ( n17291,n17292,n17293 );
   nand U17037 ( n17287,n17294,p2_datao_reg_30_ );
   nand U17038 ( n17152,n14993,n14354 );
   not U17039 ( n14993,n14571 );
   nand U17040 ( n14571,n17295,n17296 );
   nand U17041 ( n17296,n17289,n11795 );
   xor U17042 ( n11795,n17297,n17298 );
   and U17043 ( n17297,n17299,n17300 );
   nand U17044 ( n17295,n17294,p2_datao_reg_29_ );
   nand U17045 ( n17154,n16268,n14549 );
   nand U17046 ( n14549,n17301,n17302 );
   nand U17047 ( n17302,n17289,n11811 );
   and U17048 ( n11811,n17303,n17304,n17305,n17306 );
   nand U17049 ( n17306,n17293,n17307,n17308 );
   not U17050 ( n17293,n17309 );
   nand U17051 ( n17305,n17290,n17292,n17310 );
   not U17052 ( n17290,n17307 );
   nand U17053 ( n17307,n17299,n17311 );
   nand U17054 ( n17311,n17298,n17300 );
   nand U17055 ( n17300,n17312,n17313,n17314 );
   not U17056 ( n17314,si_29_ );
   nand U17057 ( n17313,n11808,p1_datao_reg_29_ );
   nand U17058 ( n17312,n11812,p2_datao_reg_29_ );
   and U17059 ( n17298,n17315,n17316 );
   nand U17060 ( n17316,n17317,n17318 );
   not U17061 ( n17318,si_28_ );
   or U17062 ( n17317,n17319,n17320 );
   nand U17063 ( n17315,n17320,n17319 );
   nand U17064 ( n17299,n17321,n17322,si_29_ );
   or U17065 ( n17322,n11808,p2_datao_reg_29_ );
   nand U17066 ( n17321,n11808,n12645 );
   not U17067 ( n12645,p1_datao_reg_29_ );
   nand U17068 ( n17304,n17309,n17310 );
   nor U17069 ( n17309,n17323,si_30_ );
   or U17070 ( n17303,n17292,n17310 );
   not U17071 ( n17310,n17308 );
   xor U17072 ( n17308,si_31_,n17324 );
   nand U17073 ( n17324,n17325,n17326 );
   nand U17074 ( n17326,n11808,p1_datao_reg_31_ );
   nand U17075 ( n17325,n11812,p2_datao_reg_31_ );
   nand U17076 ( n17292,si_30_,n17323 );
   nand U17077 ( n17323,n17327,n17328 );
   nand U17078 ( n17328,n11808,p1_datao_reg_30_ );
   nand U17079 ( n17327,n11812,p2_datao_reg_30_ );
   nand U17080 ( n17301,n17294,p2_datao_reg_31_ );
   not U17081 ( n16268,n14348 );
   nand U17082 ( n14348,n17329,n17330,n17331 );
   nand U17083 ( n17331,p1_reg2_reg_31_,n17284 );
   nand U17084 ( n17330,p1_reg0_reg_31_,n17285 );
   nand U17085 ( n17329,p1_reg1_reg_31_,n17286 );
   and U17086 ( n16822,n17164,p1_u3086 );
   nand U17087 ( n17164,p1_b_reg,n17332 );
   nand U17088 ( n17332,n17333,n17334,p1_state_reg );
   nand U17089 ( n17334,n16821,n17335 );
   nand U17090 ( n17335,n14966,n17336,n16188,n17337 );
   nor U17091 ( n17337,n16768,n17338 );
   nand U17092 ( n17333,n14966,n16817 );
   nor U17093 ( n17342,n17343,n17344,n17345 );
   nor U17094 ( n17345,n14755,n17346 );
   not U17095 ( n14755,n14393 );
   and U17096 ( n17344,n17347,n15731 );
   nor U17097 ( n17343,p1_state_reg,n17348 );
   nand U17098 ( n17341,n17349,n15722 );
   xor U17099 ( n17350,n17352,n17353 );
   xor U17100 ( n17353,n17354,n17355 );
   nand U17101 ( n17339,n17356,n14399 );
   nor U17102 ( n17360,n17361,n17362,n17363 );
   nor U17103 ( n17363,n14609,n17346 );
   nor U17104 ( n17362,n14640,n17364 );
   nor U17105 ( n17361,p1_state_reg,n17365 );
   nand U17106 ( n17359,n17349,n14610 );
   nand U17107 ( n17358,n17366,n17367 );
   xor U17108 ( n17367,n17368,n17369 );
   nand U17109 ( n17369,n17370,n17371 );
   nand U17110 ( n17368,n17372,n17373 );
   nand U17111 ( n17357,n17374,n17375 );
   nor U17112 ( n17379,n17380,n17381,n17382 );
   nor U17113 ( n17382,n14899,n17364 );
   not U17114 ( n14899,n14426 );
   nor U17115 ( n17381,n14872,n17346 );
   nor U17116 ( n17380,p1_state_reg,n17383 );
   nand U17117 ( n17378,n17384,n17347 );
   nand U17118 ( n17377,n17385,n17366 );
   xor U17119 ( n17385,n17386,n17387 );
   xor U17120 ( n17386,n17388,n17389 );
   nand U17121 ( n17376,n17349,n14873 );
   nor U17122 ( n17393,n17394,n17395,n17396 );
   nor U17123 ( n17396,n14718,n17346 );
   nor U17124 ( n17395,n14719,n17364 );
   nor U17125 ( n17394,p1_state_reg,n17397 );
   nand U17126 ( n17392,n17398,n17347 );
   or U17127 ( n17391,n17399,n17351 );
   xor U17128 ( n17399,n17400,n17401 );
   xor U17129 ( n17400,n17402,n17403 );
   nand U17130 ( n17390,n17349,n15826 );
   and U17131 ( n17409,n17410,p1_reg3_reg_2_ );
   nor U17132 ( n17408,n17351,n17411 );
   xor U17133 ( n17411,n17412,n17413 );
   xor U17134 ( n17413,n17414,n17415 );
   nor U17135 ( n17407,n14928,n17416 );
   not U17136 ( n14928,n15306 );
   nand U17137 ( n17405,n17417,n14432 );
   nand U17138 ( n17404,n17356,n14438 );
   nor U17139 ( n17421,n17422,n17423,n17424 );
   nor U17140 ( n17424,n17425,n15594 );
   nor U17141 ( n17423,n15593,n17416 );
   not U17142 ( n15593,n14812 );
   and U17143 ( n17422,p1_u3086,p1_reg3_reg_11_ );
   nand U17144 ( n17420,n17417,n14405 );
   xor U17145 ( n17426,n17427,n17428 );
   xor U17146 ( n17428,n17429,n17430 );
   nand U17147 ( n17418,n17356,n14411 );
   nor U17148 ( n17434,n17435,n17436,n17437 );
   nor U17149 ( n17437,n14641,n17346 );
   not U17150 ( n14641,n14372 );
   nor U17151 ( n17436,n14667,n17364 );
   nor U17152 ( n17435,p1_state_reg,n17438 );
   nand U17153 ( n17433,n17349,n15933 );
   or U17154 ( n17432,n17439,n17351 );
   xor U17155 ( n17439,n17440,n17441 );
   xor U17156 ( n17440,n17442,n17443 );
   nand U17157 ( n17431,n15945,n17375 );
   nor U17158 ( n17447,n17448,n17449,n17450 );
   nor U17159 ( n17450,n17425,n15657 );
   nor U17160 ( n17449,n15656,n17416 );
   not U17161 ( n15656,n14784 );
   and U17162 ( n17448,p1_u3086,p1_reg3_reg_13_ );
   nand U17163 ( n17446,n17356,n14405 );
   nand U17164 ( n17452,n17453,n17454 );
   nand U17165 ( n17454,n17455,n17456 );
   nand U17166 ( n17451,n17455,n17456,n17457 );
   nand U17167 ( n17444,n17417,n14399 );
   nor U17168 ( n17461,n17462,n17463,n17464 );
   nor U17169 ( n17464,n14667,n17346 );
   not U17170 ( n14667,n14378 );
   nor U17171 ( n17463,n14718,n17364 );
   not U17172 ( n14718,n14384 );
   nor U17173 ( n17462,p1_state_reg,n17465 );
   nand U17174 ( n17460,n17349,n14693 );
   nand U17175 ( n17459,n17366,n17466 );
   xor U17176 ( n17466,n17467,n17468 );
   xor U17177 ( n17467,n17469,n17470 );
   nand U17178 ( n17458,n17471,n17375 );
   nand U17179 ( n17475,p1_reg3_reg_0_,n17410 );
   nand U17180 ( n17474,n17366,n16770 );
   not U17181 ( n16770,n17476 );
   xor U17182 ( n17476,n17477,n17478 );
   xor U17183 ( n17478,n17479,n17480 );
   nand U17184 ( n17473,n17349,n14956 );
   nand U17185 ( n17472,n17417,n14438 );
   nor U17186 ( n17484,n17485,n17486,n17487 );
   nor U17187 ( n17487,n14834,n17364 );
   nor U17188 ( n17486,n14833,n17346 );
   not U17189 ( n14833,n14411 );
   and U17190 ( n17485,p1_u3086,p1_reg3_reg_9_ );
   nand U17191 ( n17483,n15544,n17347 );
   nand U17192 ( n17482,n17488,n17366 );
   xor U17193 ( n17488,n17489,n17490 );
   xor U17194 ( n17489,n17491,n17492 );
   nand U17195 ( n17481,n17349,n15532 );
   and U17196 ( n17499,n17366,n17500 );
   xor U17197 ( n17500,n17501,n17502 );
   xor U17198 ( n17501,n17503,n17504 );
   nor U17199 ( n17498,n17425,n15361 );
   not U17200 ( n15361,n17505 );
   nor U17201 ( n17497,n14901,n17416 );
   not U17202 ( n14901,n15376 );
   nand U17203 ( n17495,p1_reg3_reg_4_,p1_u3086 );
   nand U17204 ( n17494,n17417,n14426 );
   nand U17205 ( n17493,n17356,n14432 );
   nor U17206 ( n17509,n17510,n17511,n17512 );
   nor U17207 ( n17512,n14640,n17346 );
   not U17208 ( n14640,n14366 );
   nor U17209 ( n17511,n14642,n17416 );
   not U17210 ( n14642,n16004 );
   nor U17211 ( n17510,p1_state_reg,n17513 );
   nand U17212 ( n17508,n17356,n14372 );
   nand U17213 ( n17507,n17366,n17514 );
   xor U17214 ( n17514,n17515,n17516 );
   nand U17215 ( n17515,n17517,n17518 );
   nand U17216 ( n17506,n15995,n17375 );
   nor U17217 ( n17522,n17523,n17524,n17525 );
   nor U17218 ( n17525,n17425,n15784 );
   not U17219 ( n15784,n17526 );
   nor U17220 ( n17524,n15783,n17416 );
   not U17221 ( n15783,n14734 );
   and U17222 ( n17523,p1_u3086,p1_reg3_reg_17_ );
   nand U17223 ( n17521,n17356,n14393 );
   nand U17224 ( n17528,n17529,n17530 );
   nand U17225 ( n17530,n17531,n17532 );
   nand U17226 ( n17527,n17531,n17532,n17533 );
   nand U17227 ( n17519,n17417,n14387 );
   nor U17228 ( n17537,n17538,n17539,n17540 );
   nor U17229 ( n17540,n14884,n17364 );
   nor U17230 ( n17539,n14883,n17346 );
   and U17231 ( n17538,p1_u3086,p1_reg3_reg_5_ );
   nand U17232 ( n17536,n15402,n17347 );
   nand U17233 ( n17535,n17541,n17366 );
   xor U17234 ( n17541,n17542,n17543 );
   xor U17235 ( n17542,n17544,n17545 );
   nand U17236 ( n17534,n17349,n15392 );
   nor U17237 ( n17549,n17550,n17551,n17552 );
   nor U17238 ( n17552,n14719,n17346 );
   not U17239 ( n14719,n14390 );
   nor U17240 ( n17551,n17425,n15741 );
   not U17241 ( n15741,n17553 );
   nor U17242 ( n17550,p1_state_reg,n17554 );
   nand U17243 ( n17548,n17349,n14745 );
   xor U17244 ( n17555,n17556,n17557 );
   xor U17245 ( n17557,n17558,n17559 );
   nand U17246 ( n17546,n17356,n14396 );
   nor U17247 ( n17563,n17564,n17565,n17566 );
   nor U17248 ( n17566,n14620,n17346 );
   nor U17249 ( n17565,n14624,n17416 );
   not U17250 ( n14624,n16017 );
   and U17251 ( n17564,p1_u3086,p1_reg3_reg_25_ );
   nand U17252 ( n17562,n17356,n14369 );
   nand U17253 ( n17561,n17366,n17567 );
   nand U17254 ( n17567,n17568,n17569 );
   nand U17255 ( n17569,n17570,n17373 );
   not U17256 ( n17570,n17372 );
   nand U17257 ( n17568,n17571,n17572 );
   nand U17258 ( n17572,n17573,n17517 );
   xor U17259 ( n17571,n17574,n17575 );
   nand U17260 ( n17560,n16014,n17375 );
   nor U17261 ( n17579,n17580,n17581,n17582 );
   nor U17262 ( n17582,n14794,n17346 );
   nor U17263 ( n17581,n14795,n17364 );
   nor U17264 ( n17580,p1_state_reg,n17583 );
   nand U17265 ( n17578,n15647,n17347 );
   nand U17266 ( n17577,n17366,n17584 );
   xor U17267 ( n17584,n17585,n17586 );
   xor U17268 ( n17585,n17587,n17588 );
   nand U17269 ( n17576,n17349,n15640 );
   nor U17270 ( n17592,n17593,n17594,n17595 );
   nor U17271 ( n17595,n14679,n17416 );
   not U17272 ( n14679,n16882 );
   nor U17273 ( n17594,n14703,n17364 );
   not U17274 ( n14703,n14381 );
   nor U17275 ( n17593,p1_state_reg,n17596 );
   nand U17276 ( n17591,n17417,n14375 );
   nand U17277 ( n17590,n17597,n17598,n17366 );
   nand U17278 ( n17598,n17599,n17600 );
   nand U17279 ( n17600,n17601,n17602 );
   nand U17280 ( n17597,n17601,n17602,n17603 );
   nand U17281 ( n17589,n15892,n17375 );
   and U17282 ( n17609,n17410,p1_reg3_reg_1_ );
   nand U17283 ( n17410,n17425,p1_state_reg );
   nor U17284 ( n17608,n17351,n17610 );
   xor U17285 ( n17610,n17611,n17612 );
   xor U17286 ( n17611,n17613,n17614 );
   nor U17287 ( n17607,n14943,n17416 );
   not U17288 ( n14943,n15281 );
   nand U17289 ( n17605,n17417,n14435 );
   nand U17290 ( n17604,n17356,n14441 );
   nor U17291 ( n17618,n17619,n17620,n17621 );
   nor U17292 ( n17621,n14872,n17364 );
   not U17293 ( n14872,n14420 );
   nor U17294 ( n17620,n17425,n15491 );
   not U17295 ( n15491,n17622 );
   nor U17296 ( n17619,p1_state_reg,n17623 );
   nand U17297 ( n17617,n17417,n14414 );
   or U17298 ( n17616,n17624,n17351 );
   xor U17299 ( n17624,n17625,n17626 );
   xor U17300 ( n17625,n17627,n17628 );
   nand U17301 ( n17615,n17349,n14850 );
   nor U17302 ( n17632,n17633,n17634,n17635 );
   nor U17303 ( n17635,n14609,n17364 );
   not U17304 ( n14609,n14360 );
   and U17305 ( n17634,n17375,n16113 );
   nor U17306 ( n17633,p1_state_reg,n17636 );
   nand U17307 ( n17631,n17349,n14584 );
   nand U17308 ( n17638,n17639,n17640 );
   nand U17309 ( n17640,n17641,n17642 );
   or U17310 ( n17642,n17643,n17644 );
   not U17311 ( n17639,n17645 );
   nand U17312 ( n17637,n17645,n17646 );
   nand U17313 ( n17646,n17647,n17648 );
   nand U17314 ( n17648,n17643,n17641 );
   not U17315 ( n17641,n17649 );
   xor U17316 ( n17645,n17650,n17651 );
   nand U17317 ( n17651,n17652,n17653 );
   nand U17318 ( n17653,n17654,n14584 );
   nand U17319 ( n17652,n17655,n14357 );
   xor U17320 ( n17650,n17656,n17657 );
   nand U17321 ( n17656,n17658,n17659 );
   nand U17322 ( n17659,n17660,n14584 );
   nand U17323 ( n14584,n17661,n17662 );
   nand U17324 ( n17662,n17289,n11788 );
   xor U17325 ( n11788,n17320,n17663 );
   xor U17326 ( n17663,si_28_,n17319 );
   nand U17327 ( n17319,n17664,n17665 );
   nand U17328 ( n17665,n17666,n17667 );
   not U17329 ( n17667,si_27_ );
   or U17330 ( n17666,n17668,n17669 );
   nand U17331 ( n17664,n17669,n17668 );
   nand U17332 ( n17320,n17670,n17671 );
   or U17333 ( n17671,n11808,p2_datao_reg_28_ );
   nand U17334 ( n17670,n11808,n13754 );
   not U17335 ( n13754,p1_datao_reg_28_ );
   nand U17336 ( n17661,n17294,p2_datao_reg_28_ );
   nand U17337 ( n17658,n17654,n14357 );
   nand U17338 ( n17629,n17417,n14354 );
   nand U17339 ( n14354,n17672,n17673,n17674,n17675 );
   nand U17340 ( n17675,n17676,n14989 );
   nor U17341 ( n14989,n17677,n17678,n17636 );
   not U17342 ( n17636,p1_reg3_reg_28_ );
   nand U17343 ( n17674,p1_reg0_reg_29_,n17285 );
   nand U17344 ( n17673,p1_reg1_reg_29_,n17286 );
   nand U17345 ( n17672,p1_reg2_reg_29_,n17284 );
   nor U17346 ( n17682,n17683,n17684,n17685 );
   nor U17347 ( n17685,n17425,n15837 );
   nor U17348 ( n17684,n14705,n17416 );
   not U17349 ( n14705,n15840 );
   and U17350 ( n17683,p1_u3086,p1_reg3_reg_19_ );
   nand U17351 ( n17681,n17417,n14381 );
   xor U17352 ( n17686,n17687,n17688 );
   xor U17353 ( n17687,n17689,n17690 );
   nand U17354 ( n17679,n17356,n14387 );
   nor U17355 ( n17696,n14915,n17416 );
   not U17356 ( n14915,n15338 );
   nor U17357 ( n17695,n17351,n17697,n17698 );
   nor U17358 ( n17698,n17699,n17700,n17701 );
   not U17359 ( n17699,n17702 );
   nor U17360 ( n17697,n17703,n17702 );
   nor U17361 ( n17703,n17700,n17701 );
   nor U17362 ( n17694,n14884,n17346 );
   not U17363 ( n14884,n14429 );
   nand U17364 ( n17692,n17356,n14435 );
   nand U17365 ( n16730,p1_reg3_reg_3_,p1_u3086 );
   nand U17366 ( n17691,n17347,n15350 );
   nor U17367 ( n17707,n17708,n17709,n17710 );
   nor U17368 ( n17710,n14795,n17346 );
   not U17369 ( n14795,n14408 );
   nor U17370 ( n17709,n17425,n15554 );
   not U17371 ( n17425,n17347 );
   nor U17372 ( n17708,p1_state_reg,n17711 );
   nand U17373 ( n17706,n17349,n14823 );
   xor U17374 ( n17712,n17713,n17714 );
   xor U17375 ( n17714,n17715,n17716 );
   nand U17376 ( n17704,n17356,n14414 );
   nor U17377 ( n17720,n17721,n17722,n17723 );
   nor U17378 ( n17723,n14621,n17346 );
   not U17379 ( n14621,n14369 );
   nor U17380 ( n17722,n15954,n17416 );
   not U17381 ( n15954,n14657 );
   nor U17382 ( n17721,p1_state_reg,n17724 );
   nand U17383 ( n17719,n17356,n14375 );
   or U17384 ( n17718,n17725,n17351 );
   xor U17385 ( n17725,n17726,n17727 );
   xor U17386 ( n17727,n17728,n17729 );
   nand U17387 ( n17717,n15955,n17375 );
   nor U17388 ( n17733,n17734,n17735,n17736 );
   nor U17389 ( n17736,n14770,n17346 );
   not U17390 ( n14770,n14396 );
   nor U17391 ( n17735,n14794,n17364 );
   not U17392 ( n14794,n14402 );
   nor U17393 ( n17734,p1_state_reg,n17737 );
   nand U17394 ( n17732,n17738,n17347 );
   or U17395 ( n17731,n17739,n17351 );
   xor U17396 ( n17739,n17740,n17741 );
   xor U17397 ( n17740,n17742,n17743 );
   nand U17398 ( n17730,n17349,n15694 );
   nor U17399 ( n17747,n17748,n17749,n17750 );
   nor U17400 ( n17750,n14620,n17364 );
   not U17401 ( n14620,n14363 );
   nor U17402 ( n17749,n16073,n17416 );
   not U17403 ( n16073,n14597 );
   nor U17404 ( n17748,p1_state_reg,n17677 );
   nand U17405 ( n17746,n17417,n14357 );
   nand U17406 ( n14357,n17751,n17752,n17753,n17754 );
   nand U17407 ( n17754,n17676,n16113 );
   xor U17408 ( n16113,n17755,p1_reg3_reg_28_ );
   nor U17409 ( n17755,n17678,n17677 );
   nand U17410 ( n17753,p1_reg0_reg_28_,n17285 );
   nand U17411 ( n17752,p1_reg1_reg_28_,n17286 );
   nand U17412 ( n17751,p1_reg2_reg_28_,n17284 );
   nand U17413 ( n17745,n17756,n17366 );
   xor U17414 ( n17756,n17757,n17643 );
   nand U17415 ( n17643,n17371,n17758 );
   nand U17416 ( n17758,n17370,n17373,n17372 );
   nand U17417 ( n17372,n17573,n17517,n17759 );
   nand U17418 ( n17759,n17760,n17575 );
   nand U17419 ( n17517,n17761,n17762 );
   xor U17420 ( n17761,n17763,n17657 );
   nand U17421 ( n17573,n17764,n17518 );
   nand U17422 ( n17518,n17765,n17766 );
   not U17423 ( n17766,n17762 );
   nand U17424 ( n17762,n17767,n17768 );
   nand U17425 ( n17768,n17654,n16004 );
   nand U17426 ( n17767,n17655,n14369 );
   xor U17427 ( n17765,n17479,n17763 );
   nand U17428 ( n17763,n17769,n17770 );
   nand U17429 ( n17770,n17660,n16004 );
   nand U17430 ( n16004,n17771,n17772 );
   nand U17431 ( n17772,n17289,n11751 );
   xor U17432 ( n11751,n17773,n17774 );
   xor U17433 ( n17774,si_24_,n17775 );
   nand U17434 ( n17771,n17294,p2_datao_reg_24_ );
   nand U17435 ( n17769,n17654,n14369 );
   nand U17436 ( n14369,n17776,n17777,n17778,n17779 );
   nand U17437 ( n17779,n15995,n17676 );
   nor U17438 ( n15995,n17780,n17781 );
   and U17439 ( n17780,n17513,n17782 );
   nand U17440 ( n17782,p1_reg3_reg_23_,n17783 );
   nand U17441 ( n17778,p1_reg0_reg_24_,n17285 );
   nand U17442 ( n17777,p1_reg1_reg_24_,n17286 );
   nand U17443 ( n17776,p1_reg2_reg_24_,n17284 );
   not U17444 ( n17764,n17516 );
   nand U17445 ( n17516,n17784,n17785 );
   nand U17446 ( n17785,n17726,n17786 );
   or U17447 ( n17786,n17729,n17728 );
   xor U17448 ( n17726,n17479,n17787 );
   nand U17449 ( n17787,n17788,n17789 );
   nand U17450 ( n17789,n17660,n14657 );
   nand U17451 ( n17788,n17654,n14372 );
   nand U17452 ( n17784,n17728,n17729 );
   nand U17453 ( n17729,n17790,n17791 );
   nand U17454 ( n17791,n17792,n17443 );
   nand U17455 ( n17443,n17793,n17602 );
   nand U17456 ( n17602,n17794,n17795 );
   not U17457 ( n17795,n17796 );
   xor U17458 ( n17794,n17479,n17797 );
   nand U17459 ( n17793,n17599,n17601 );
   nand U17460 ( n17601,n17798,n17796 );
   nand U17461 ( n17796,n17799,n17800 );
   nand U17462 ( n17800,n17654,n16882 );
   nand U17463 ( n17799,n17655,n14378 );
   xor U17464 ( n17798,n17797,n17657 );
   nand U17465 ( n17797,n17801,n17802 );
   nand U17466 ( n17802,n17660,n16882 );
   nand U17467 ( n16882,n17803,n17804 );
   nand U17468 ( n17804,n17289,n11727 );
   xor U17469 ( n11727,n17805,n17806 );
   xor U17470 ( n17806,si_21_,n17807 );
   nand U17471 ( n17803,n17294,p2_datao_reg_21_ );
   nand U17472 ( n17801,n17654,n14378 );
   nand U17473 ( n14378,n17808,n17809,n17810,n17811 );
   nand U17474 ( n17811,n17676,n15892 );
   xor U17475 ( n15892,n17596,n17812 );
   nand U17476 ( n17810,p1_reg0_reg_21_,n17285 );
   nand U17477 ( n17809,p1_reg1_reg_21_,n17286 );
   nand U17478 ( n17808,p1_reg2_reg_21_,n17284 );
   not U17479 ( n17599,n17603 );
   nand U17480 ( n17603,n17813,n17814 );
   nand U17481 ( n17814,n17815,n17470 );
   nand U17482 ( n17470,n17816,n17817 );
   nand U17483 ( n17817,n17654,n14693 );
   nand U17484 ( n17816,n17655,n14381 );
   nand U17485 ( n17815,n17469,n17468 );
   or U17486 ( n17813,n17468,n17469 );
   and U17487 ( n17469,n17818,n17819 );
   nand U17488 ( n17819,n17820,n17821 );
   or U17489 ( n17821,n17690,n17688 );
   not U17490 ( n17820,n17689 );
   nand U17491 ( n17689,n17822,n17823 );
   nand U17492 ( n17823,n17824,n17403 );
   nand U17493 ( n17403,n17825,n17532 );
   nand U17494 ( n17532,n17826,n17827 );
   not U17495 ( n17827,n17828 );
   xor U17496 ( n17826,n17479,n17829 );
   nand U17497 ( n17825,n17529,n17531 );
   nand U17498 ( n17531,n17830,n17828 );
   nand U17499 ( n17828,n17831,n17832 );
   nand U17500 ( n17832,n17654,n14734 );
   nand U17501 ( n17831,n17655,n14390 );
   xor U17502 ( n17830,n17829,n17657 );
   nand U17503 ( n17829,n17833,n17834 );
   nand U17504 ( n17834,n17660,n14734 );
   nand U17505 ( n14734,n17835,n17836,n17837 );
   nand U17506 ( n17837,n17294,p2_datao_reg_17_ );
   nand U17507 ( n17836,n16340,n16273 );
   not U17508 ( n16340,n16362 );
   nand U17509 ( n16362,n17838,n17839,n15151 );
   nand U17510 ( n17839,n15143,n15241 );
   nand U17511 ( n17838,p1_ir_reg_17_,n15135,p1_ir_reg_31_ );
   nand U17512 ( n17835,n17289,n11694 );
   not U17513 ( n11694,n13910 );
   xor U17514 ( n13910,n17840,n17841 );
   xor U17515 ( n17840,n17842,n17843 );
   nand U17516 ( n17833,n17654,n14390 );
   nand U17517 ( n14390,n17844,n17845,n17846,n17847 );
   nand U17518 ( n17847,n17676,n17526 );
   xor U17519 ( n17526,p1_reg3_reg_17_,n17848 );
   nand U17520 ( n17846,p1_reg0_reg_17_,n17285 );
   nand U17521 ( n17845,p1_reg1_reg_17_,n17286 );
   nand U17522 ( n17844,p1_reg2_reg_17_,n17284 );
   not U17523 ( n17529,n17533 );
   nand U17524 ( n17533,n17849,n17850 );
   nand U17525 ( n17850,n17556,n17851 );
   nand U17526 ( n17851,n17558,n17559 );
   xor U17527 ( n17556,n17657,n17852 );
   nand U17528 ( n17852,n17853,n17854 );
   nand U17529 ( n17854,n17660,n14745 );
   nand U17530 ( n17853,n17654,n14393 );
   or U17531 ( n17849,n17559,n17558 );
   and U17532 ( n17558,n17855,n17856 );
   nand U17533 ( n17856,n17654,n14745 );
   nand U17534 ( n14745,n17857,n17858,n17859 );
   nand U17535 ( n17859,n17294,p2_datao_reg_16_ );
   nand U17536 ( n17858,n16361,n16273 );
   not U17537 ( n16361,n16366 );
   nand U17538 ( n16366,n17860,n17861 );
   or U17539 ( n17861,p1_ir_reg_16_,p1_ir_reg_31_ );
   nand U17540 ( n17860,p1_ir_reg_31_,n17862 );
   nand U17541 ( n17862,n15134,n15135 );
   not U17542 ( n15135,n15142 );
   nand U17543 ( n15134,p1_ir_reg_16_,n17863 );
   nand U17544 ( n17857,n17289,n11684 );
   not U17545 ( n11684,n13922 );
   xor U17546 ( n13922,n17864,n17865 );
   xor U17547 ( n17864,n17866,n17867 );
   nand U17548 ( n17855,n17655,n14393 );
   nand U17549 ( n14393,n17868,n17869,n17870,n17871 );
   nand U17550 ( n17871,n17553,n17676 );
   nor U17551 ( n17553,n17872,n17848 );
   and U17552 ( n17872,n17554,n17873 );
   or U17553 ( n17873,n17348,n17874 );
   nand U17554 ( n17870,p1_reg0_reg_16_,n17285 );
   nand U17555 ( n17869,p1_reg1_reg_16_,n17286 );
   nand U17556 ( n17868,p1_reg2_reg_16_,n17284 );
   nand U17557 ( n17559,n17875,n17876 );
   nand U17558 ( n17876,n17352,n17877 );
   nand U17559 ( n17877,n17355,n17354 );
   xor U17560 ( n17352,n17479,n17878 );
   nand U17561 ( n17878,n17879,n17880 );
   nand U17562 ( n17880,n17660,n15722 );
   nand U17563 ( n17879,n17654,n14396 );
   or U17564 ( n17875,n17354,n17355 );
   and U17565 ( n17355,n17881,n17882 );
   nand U17566 ( n17882,n17883,n17743 );
   nand U17567 ( n17743,n17884,n17456 );
   nand U17568 ( n17456,n17885,n17886 );
   not U17569 ( n17886,n17887 );
   xor U17570 ( n17885,n17479,n17888 );
   nand U17571 ( n17884,n17453,n17455 );
   nand U17572 ( n17455,n17889,n17887 );
   nand U17573 ( n17887,n17890,n17891 );
   nand U17574 ( n17891,n17654,n14784 );
   nand U17575 ( n17890,n17655,n14402 );
   xor U17576 ( n17889,n17888,n17657 );
   nand U17577 ( n17888,n17892,n17893 );
   nand U17578 ( n17893,n17660,n14784 );
   nand U17579 ( n14784,n17894,n17895,n17896 );
   nand U17580 ( n17896,n17294,p2_datao_reg_13_ );
   nand U17581 ( n17895,n16450,n16273 );
   not U17582 ( n16450,n16472 );
   nand U17583 ( n16472,n17897,n17898,n17899 );
   nand U17584 ( n17898,n15114,n15241 );
   nand U17585 ( n17897,p1_ir_reg_13_,n15106,p1_ir_reg_31_ );
   nand U17586 ( n17894,n17289,n11660 );
   nand U17587 ( n11660,n17900,n17901 );
   nand U17588 ( n17901,n17902,n17903 );
   nand U17589 ( n17902,n17904,n17905 );
   nand U17590 ( n17900,n17906,n17907 );
   xor U17591 ( n17907,si_13_,n17908 );
   not U17592 ( n17906,n17903 );
   nand U17593 ( n17903,n17909,n17910 );
   nand U17594 ( n17910,n17911,n17912 );
   nand U17595 ( n17892,n17654,n14402 );
   nand U17596 ( n14402,n17913,n17914,n17915,n17916 );
   nand U17597 ( n17916,n17676,n17917 );
   not U17598 ( n17917,n15657 );
   xor U17599 ( n15657,p1_reg3_reg_13_,n17918 );
   nand U17600 ( n17915,p1_reg0_reg_13_,n17285 );
   nand U17601 ( n17914,p1_reg1_reg_13_,n17286 );
   nand U17602 ( n17913,p1_reg2_reg_13_,n17284 );
   not U17603 ( n17453,n17457 );
   nand U17604 ( n17457,n17919,n17920 );
   nand U17605 ( n17920,n17921,n17588 );
   nand U17606 ( n17588,n17922,n17923 );
   nand U17607 ( n17923,n17654,n15640 );
   nand U17608 ( n17922,n17655,n14405 );
   nand U17609 ( n17921,n17587,n17586 );
   or U17610 ( n17919,n17586,n17587 );
   and U17611 ( n17587,n17924,n17925 );
   nand U17612 ( n17925,n17430,n17926 );
   or U17613 ( n17926,n17429,n17427 );
   and U17614 ( n17430,n17927,n17928 );
   nand U17615 ( n17928,n17713,n17929 );
   or U17616 ( n17929,n17716,n17715 );
   xor U17617 ( n17713,n17479,n17930 );
   nand U17618 ( n17930,n17931,n17932 );
   nand U17619 ( n17932,n17660,n14823 );
   nand U17620 ( n17931,n17654,n14411 );
   nand U17621 ( n17927,n17715,n17716 );
   nand U17622 ( n17716,n17933,n17934 );
   nand U17623 ( n17934,n17935,n17936 );
   or U17624 ( n17936,n17491,n17490 );
   not U17625 ( n17935,n17492 );
   nand U17626 ( n17492,n17937,n17938 );
   nand U17627 ( n17938,n17655,n14414 );
   nand U17628 ( n17937,n17654,n15532 );
   nand U17629 ( n17933,n17490,n17491 );
   nand U17630 ( n17491,n17939,n17940 );
   nand U17631 ( n17940,n17941,n17627 );
   nand U17632 ( n17627,n17942,n17943 );
   nand U17633 ( n17942,n17944,n17945 );
   nand U17634 ( n17941,n17626,n17628 );
   or U17635 ( n17939,n17628,n17626 );
   xor U17636 ( n17626,n17657,n17946 );
   nand U17637 ( n17946,n17947,n17948 );
   nand U17638 ( n17948,n17660,n14850 );
   nand U17639 ( n17947,n17654,n14417 );
   nand U17640 ( n17628,n17949,n17950 );
   nand U17641 ( n17950,n17654,n14850 );
   nand U17642 ( n14850,n17951,n17952,n17953 );
   nand U17643 ( n17953,n17294,p2_datao_reg_8_ );
   nand U17644 ( n17952,n16595,n16273 );
   not U17645 ( n16595,n16605 );
   nand U17646 ( n16605,n17954,n17955 );
   or U17647 ( n17955,p1_ir_reg_31_,p1_ir_reg_8_ );
   nand U17648 ( n17954,p1_ir_reg_31_,n17956 );
   nand U17649 ( n17956,n15083,n15084 );
   nand U17650 ( n15083,p1_ir_reg_8_,n17957 );
   nand U17651 ( n17951,n17289,n11617 );
   xor U17652 ( n11617,n17958,n17959 );
   and U17653 ( n17958,n17960,n17961 );
   nand U17654 ( n17949,n17655,n14417 );
   xor U17655 ( n17490,n17479,n17962 );
   nand U17656 ( n17962,n17963,n17964 );
   nand U17657 ( n17964,n17660,n15532 );
   nand U17658 ( n15532,n17965,n17966,n17967 );
   nand U17659 ( n17967,n17294,p2_datao_reg_9_ );
   nand U17660 ( n17966,n16575,n16273 );
   not U17661 ( n16575,n16576 );
   nand U17662 ( n16576,n17968,n17969 );
   nand U17663 ( n17969,n15241,n17970 );
   or U17664 ( n17968,n15089,n15241 );
   xor U17665 ( n15089,p1_ir_reg_9_,n15084 );
   nand U17666 ( n17965,n17289,n11626 );
   xor U17667 ( n11626,n17971,n17972 );
   and U17668 ( n17971,n17973,n17974 );
   nand U17669 ( n17963,n17654,n14414 );
   nand U17670 ( n14414,n17975,n17976,n17977,n17978 );
   nand U17671 ( n17978,n17676,n15544 );
   xor U17672 ( n15544,p1_reg3_reg_9_,n17979 );
   nand U17673 ( n17977,p1_reg0_reg_9_,n17285 );
   nand U17674 ( n17976,p1_reg1_reg_9_,n17286 );
   nand U17675 ( n17975,p1_reg2_reg_9_,n17284 );
   and U17676 ( n17715,n17980,n17981 );
   nand U17677 ( n17981,n17655,n14411 );
   nand U17678 ( n14411,n17982,n17983,n17984,n17985 );
   nand U17679 ( n17985,n17986,n17676 );
   not U17680 ( n17986,n15554 );
   nand U17681 ( n15554,n17987,n17988 );
   nand U17682 ( n17987,n17711,n17989 );
   nand U17683 ( n17989,p1_reg3_reg_9_,n17979 );
   not U17684 ( n17711,p1_reg3_reg_10_ );
   nand U17685 ( n17984,p1_reg0_reg_10_,n17285 );
   nand U17686 ( n17983,p1_reg1_reg_10_,n17286 );
   nand U17687 ( n17982,p1_reg2_reg_10_,n17284 );
   nand U17688 ( n17980,n17654,n14823 );
   nand U17689 ( n14823,n17990,n17991,n17992 );
   nand U17690 ( n17992,n17294,p2_datao_reg_10_ );
   nand U17691 ( n17991,n16531,n16273 );
   not U17692 ( n16531,n16555 );
   nand U17693 ( n16555,n17993,n17994 );
   or U17694 ( n17994,p1_ir_reg_10_,p1_ir_reg_31_ );
   nand U17695 ( n17993,p1_ir_reg_31_,n15095 );
   nand U17696 ( n15095,n17995,n17996 );
   nand U17697 ( n17996,p1_ir_reg_10_,n17997 );
   nand U17698 ( n17997,n17998,n17970 );
   not U17699 ( n17970,p1_ir_reg_9_ );
   nand U17700 ( n17990,n17289,n11633 );
   xor U17701 ( n11633,n17999,n18000 );
   xor U17702 ( n18000,si_10_,n18001 );
   nand U17703 ( n17924,n17427,n17429 );
   nand U17704 ( n17429,n18002,n18003 );
   nand U17705 ( n18003,n17655,n14408 );
   nand U17706 ( n18002,n17654,n14812 );
   xor U17707 ( n17427,n17657,n18004 );
   nand U17708 ( n18004,n18005,n18006 );
   nand U17709 ( n18006,n17660,n14812 );
   nand U17710 ( n14812,n18007,n18008,n18009 );
   nand U17711 ( n18009,n17294,p2_datao_reg_11_ );
   nand U17712 ( n18008,n16508,n16273 );
   not U17713 ( n16508,n16506 );
   nand U17714 ( n16506,n18010,n18011 );
   nand U17715 ( n18011,n18012,n15241 );
   or U17716 ( n18010,n15100,n15241 );
   xor U17717 ( n15100,n18013,n18012 );
   nand U17718 ( n18007,n17289,n11643 );
   xor U17719 ( n11643,n18014,n18015 );
   nor U17720 ( n18014,n18016,n18017 );
   nand U17721 ( n18005,n17654,n14408 );
   nand U17722 ( n14408,n18018,n18019,n18020,n18021 );
   nand U17723 ( n18021,n17676,n18022 );
   not U17724 ( n18022,n15594 );
   xor U17725 ( n15594,p1_reg3_reg_11_,n17988 );
   nand U17726 ( n18020,p1_reg0_reg_11_,n17285 );
   nand U17727 ( n18019,p1_reg1_reg_11_,n17286 );
   nand U17728 ( n18018,p1_reg2_reg_11_,n17284 );
   xor U17729 ( n17586,n17479,n18023 );
   nand U17730 ( n18023,n18024,n18025 );
   nand U17731 ( n18025,n17660,n15640 );
   nand U17732 ( n15640,n18026,n18027,n18028 );
   nand U17733 ( n18028,n17294,p2_datao_reg_12_ );
   nand U17734 ( n18027,n16492,n16273 );
   not U17735 ( n16492,n16494 );
   nand U17736 ( n16494,n18029,n18030 );
   or U17737 ( n18030,p1_ir_reg_12_,p1_ir_reg_31_ );
   nand U17738 ( n18029,p1_ir_reg_31_,n18031 );
   nand U17739 ( n18031,n15105,n15106 );
   not U17740 ( n15106,n15113 );
   nand U17741 ( n15105,p1_ir_reg_12_,n18032 );
   nand U17742 ( n18032,n18013,n18012 );
   not U17743 ( n18012,p1_ir_reg_11_ );
   nand U17744 ( n18026,n17289,n11650 );
   xor U17745 ( n11650,n18033,n17911 );
   nand U17746 ( n17911,n18034,n18035 );
   nand U17747 ( n18035,n18036,n18015 );
   and U17748 ( n18033,n17909,n17912 );
   nand U17749 ( n18024,n17654,n14405 );
   nand U17750 ( n14405,n18037,n18038,n18039,n18040 );
   nand U17751 ( n18040,n15647,n17676 );
   and U17752 ( n15647,n18041,n17918 );
   nand U17753 ( n18041,n17583,n18042 );
   nand U17754 ( n18042,p1_reg3_reg_11_,n18043 );
   not U17755 ( n17583,p1_reg3_reg_12_ );
   nand U17756 ( n18039,p1_reg0_reg_12_,n17285 );
   nand U17757 ( n18038,p1_reg1_reg_12_,n17286 );
   nand U17758 ( n18037,p1_reg2_reg_12_,n17284 );
   nand U17759 ( n17883,n17741,n17742 );
   or U17760 ( n17881,n17742,n17741 );
   xor U17761 ( n17741,n17657,n18044 );
   nand U17762 ( n18044,n18045,n18046 );
   nand U17763 ( n18046,n17660,n15694 );
   nand U17764 ( n18045,n17654,n14399 );
   nand U17765 ( n17742,n18047,n18048 );
   nand U17766 ( n18048,n17654,n15694 );
   nand U17767 ( n15694,n18049,n18050,n18051 );
   nand U17768 ( n18051,n17294,p2_datao_reg_14_ );
   nand U17769 ( n18050,n16424,n16273 );
   not U17770 ( n16424,n16435 );
   nand U17771 ( n16435,n18052,n18053 );
   or U17772 ( n18053,p1_ir_reg_14_,p1_ir_reg_31_ );
   nand U17773 ( n18052,p1_ir_reg_31_,n15120 );
   nand U17774 ( n15120,n15128,n18054 );
   nand U17775 ( n18054,p1_ir_reg_14_,n17899 );
   nand U17776 ( n18049,n17289,n11667 );
   xor U17777 ( n11667,n18055,n18056 );
   xor U17778 ( n18056,si_14_,n18057 );
   nand U17779 ( n18057,n18058,n18059 );
   nand U17780 ( n18047,n17655,n14399 );
   nand U17781 ( n14399,n18060,n18061,n18062,n18063 );
   nand U17782 ( n18063,n17738,n17676 );
   not U17783 ( n17738,n15700 );
   nand U17784 ( n15700,n18064,n17874 );
   nand U17785 ( n18064,n17737,n18065 );
   nand U17786 ( n18065,p1_reg3_reg_13_,n18066 );
   not U17787 ( n17737,p1_reg3_reg_14_ );
   nand U17788 ( n18062,p1_reg0_reg_14_,n17285 );
   nand U17789 ( n18061,p1_reg1_reg_14_,n17286 );
   nand U17790 ( n18060,p1_reg2_reg_14_,n17284 );
   nand U17791 ( n17354,n18067,n18068 );
   nand U17792 ( n18068,n17655,n14396 );
   nand U17793 ( n14396,n18069,n18070,n18071,n18072 );
   nand U17794 ( n18072,n17676,n15731 );
   xor U17795 ( n15731,n17348,n17874 );
   nand U17796 ( n18071,p1_reg0_reg_15_,n17285 );
   nand U17797 ( n18070,p1_reg1_reg_15_,n17286 );
   nand U17798 ( n18069,p1_reg2_reg_15_,n17284 );
   nand U17799 ( n18067,n17654,n15722 );
   nand U17800 ( n15722,n18073,n18074,n18075 );
   nand U17801 ( n18075,n17294,p2_datao_reg_15_ );
   nand U17802 ( n18074,n16409,n16273 );
   not U17803 ( n16409,n16398 );
   nand U17804 ( n16398,n18076,n18077,n17863 );
   nand U17805 ( n18077,n15129,n15241 );
   nand U17806 ( n18076,p1_ir_reg_15_,n15128,p1_ir_reg_31_ );
   not U17807 ( n15128,n15127 );
   nand U17808 ( n18073,n17289,n11677 );
   not U17809 ( n11677,n14056 );
   xor U17810 ( n14056,n18078,n18079 );
   xor U17811 ( n18078,n18080,n18081 );
   nand U17812 ( n17824,n17401,n17402 );
   or U17813 ( n17822,n17402,n17401 );
   xor U17814 ( n17401,n17657,n18082 );
   nand U17815 ( n18082,n18083,n18084 );
   nand U17816 ( n18084,n17660,n15826 );
   nand U17817 ( n18083,n17654,n14387 );
   nand U17818 ( n17402,n18085,n18086 );
   nand U17819 ( n18086,n17654,n15826 );
   nand U17820 ( n15826,n18087,n18088,n18089 );
   nand U17821 ( n18089,n17294,p2_datao_reg_18_ );
   nand U17822 ( n18088,n16300,n16273 );
   not U17823 ( n16300,n16303 );
   nand U17824 ( n16303,n18090,n18091,n18092 );
   nand U17825 ( n18091,n15152,n15241 );
   nand U17826 ( n18090,p1_ir_reg_18_,n15151,p1_ir_reg_31_ );
   nand U17827 ( n18087,n17289,n11704 );
   xor U17828 ( n11704,n18093,n18094 );
   xor U17829 ( n18094,si_18_,n18095 );
   nand U17830 ( n18085,n17655,n14387 );
   nand U17831 ( n14387,n18096,n18097,n18098,n18099 );
   nand U17832 ( n18099,n17398,n17676 );
   not U17833 ( n17398,n15816 );
   nand U17834 ( n15816,n18100,n18101 );
   nand U17835 ( n18100,n17397,n18102 );
   nand U17836 ( n18102,p1_reg3_reg_17_,n17848 );
   not U17837 ( n17397,p1_reg3_reg_18_ );
   nand U17838 ( n18098,p1_reg0_reg_18_,n17285 );
   nand U17839 ( n18097,p1_reg1_reg_18_,n17286 );
   nand U17840 ( n18096,p1_reg2_reg_18_,n17284 );
   nand U17841 ( n17818,n17688,n17690 );
   nand U17842 ( n17690,n18103,n18104 );
   nand U17843 ( n18104,n17655,n14384 );
   nand U17844 ( n18103,n17654,n15840 );
   xor U17845 ( n17688,n17657,n18105 );
   nand U17846 ( n18105,n18106,n18107 );
   nand U17847 ( n18107,n17660,n15840 );
   nand U17848 ( n15840,n18108,n18109,n18110 );
   nand U17849 ( n18110,n16273,n16288 );
   nand U17850 ( n18109,n17289,n11711 );
   xor U17851 ( n11711,n18111,n18112 );
   xor U17852 ( n18112,si_19_,n18113 );
   nand U17853 ( n18108,n17294,p2_datao_reg_19_ );
   nand U17854 ( n18106,n17654,n14384 );
   nand U17855 ( n14384,n18114,n18115,n18116,n18117 );
   nand U17856 ( n18117,n17676,n18118 );
   not U17857 ( n18118,n15837 );
   xor U17858 ( n15837,p1_reg3_reg_19_,n18101 );
   nand U17859 ( n18116,p1_reg0_reg_19_,n17285 );
   nand U17860 ( n18115,p1_reg1_reg_19_,n17286 );
   nand U17861 ( n18114,p1_reg2_reg_19_,n17284 );
   xor U17862 ( n17468,n17479,n18119 );
   nand U17863 ( n18119,n18120,n18121 );
   nand U17864 ( n18121,n17660,n14693 );
   nand U17865 ( n14693,n18122,n18123 );
   nand U17866 ( n18123,n17289,n11718 );
   xor U17867 ( n11718,n18124,n18125 );
   xor U17868 ( n18125,si_20_,n18126 );
   nand U17869 ( n18122,n17294,p2_datao_reg_20_ );
   nand U17870 ( n18120,n17654,n14381 );
   nand U17871 ( n14381,n18127,n18128,n18129,n18130 );
   nand U17872 ( n18130,n17471,n17676 );
   not U17873 ( n17471,n15855 );
   nand U17874 ( n15855,n18131,n17812 );
   nand U17875 ( n18131,n17465,n18132 );
   nand U17876 ( n18132,p1_reg3_reg_19_,n18133 );
   not U17877 ( n17465,p1_reg3_reg_20_ );
   nand U17878 ( n18129,p1_reg0_reg_20_,n17285 );
   nand U17879 ( n18128,p1_reg1_reg_20_,n17286 );
   nand U17880 ( n18127,p1_reg2_reg_20_,n17284 );
   nand U17881 ( n17792,n17441,n17442 );
   or U17882 ( n17790,n17442,n17441 );
   xor U17883 ( n17441,n17657,n18134 );
   nand U17884 ( n18134,n18135,n18136 );
   nand U17885 ( n18136,n17660,n15933 );
   nand U17886 ( n18135,n17654,n14375 );
   nand U17887 ( n17442,n18137,n18138 );
   nand U17888 ( n18138,n17654,n15933 );
   nand U17889 ( n15933,n18139,n18140 );
   nand U17890 ( n18140,n17289,n11734 );
   xor U17891 ( n11734,n18141,n18142 );
   xor U17892 ( n18142,si_22_,n18143 );
   nand U17893 ( n18139,n17294,p2_datao_reg_22_ );
   nand U17894 ( n18137,n17655,n14375 );
   nand U17895 ( n14375,n18144,n18145,n18146,n18147 );
   nand U17896 ( n18147,n15945,n17676 );
   and U17897 ( n15945,n18148,n18149 );
   nand U17898 ( n18148,n17438,n18150 );
   or U17899 ( n18150,n17596,n17812 );
   nand U17900 ( n18146,p1_reg0_reg_22_,n17285 );
   nand U17901 ( n18145,p1_reg1_reg_22_,n17286 );
   nand U17902 ( n18144,p1_reg2_reg_22_,n17284 );
   and U17903 ( n17728,n18151,n18152 );
   nand U17904 ( n18152,n17655,n14372 );
   nand U17905 ( n14372,n18153,n18154,n18155,n18156 );
   nand U17906 ( n18156,n17676,n15955 );
   xor U17907 ( n15955,n17724,n18149 );
   nand U17908 ( n18155,p1_reg0_reg_23_,n17285 );
   nand U17909 ( n18154,p1_reg1_reg_23_,n17286 );
   nand U17910 ( n18153,p1_reg2_reg_23_,n17284 );
   nand U17911 ( n18151,n17654,n14657 );
   nand U17912 ( n14657,n18157,n18158 );
   nand U17913 ( n18158,n17289,n11744 );
   xor U17914 ( n11744,n18159,n18160 );
   xor U17915 ( n18160,si_23_,n18161 );
   nand U17916 ( n18157,n17294,p2_datao_reg_23_ );
   or U17917 ( n17373,n17575,n17760 );
   not U17918 ( n17760,n17574 );
   xor U17919 ( n17574,n17479,n18162 );
   nand U17920 ( n18162,n18163,n18164 );
   nand U17921 ( n18164,n17660,n16017 );
   nand U17922 ( n18163,n17654,n14366 );
   nand U17923 ( n17575,n18165,n18166 );
   nand U17924 ( n18166,n17654,n16017 );
   nand U17925 ( n16017,n18167,n18168 );
   nand U17926 ( n18168,n17289,n11761 );
   xor U17927 ( n11761,n18169,n18170 );
   xor U17928 ( n18170,si_25_,n18171 );
   nand U17929 ( n18167,n17294,p2_datao_reg_25_ );
   nand U17930 ( n18165,n17655,n14366 );
   nand U17931 ( n14366,n18172,n18173,n18174,n18175 );
   nand U17932 ( n18175,n17676,n16014 );
   xor U17933 ( n16014,p1_reg3_reg_25_,n17781 );
   nand U17934 ( n18174,p1_reg0_reg_25_,n17285 );
   nand U17935 ( n18173,p1_reg1_reg_25_,n17286 );
   nand U17936 ( n18172,p1_reg2_reg_25_,n17284 );
   nand U17937 ( n17370,n18176,n18177,n18178 );
   xor U17938 ( n18178,n17479,n18179 );
   nand U17939 ( n18177,n17654,n14610 );
   nand U17940 ( n17371,n18180,n18181,n18182 );
   xor U17941 ( n18182,n18179,n17657 );
   nand U17942 ( n18179,n18183,n18184 );
   nand U17943 ( n18184,n17660,n14610 );
   nand U17944 ( n18183,n17654,n14363 );
   nand U17945 ( n18181,n18176,n18185 );
   nand U17946 ( n18176,n17655,n14363 );
   nand U17947 ( n14363,n18186,n18187,n18188,n18189 );
   nand U17948 ( n18189,n17374,n17676 );
   not U17949 ( n17374,n16031 );
   nand U17950 ( n16031,n17678,n18190 );
   nand U17951 ( n18190,n18191,n17365 );
   nand U17952 ( n18188,p1_reg0_reg_26_,n17285 );
   nand U17953 ( n18187,p1_reg1_reg_26_,n17286 );
   nand U17954 ( n18186,p1_reg2_reg_26_,n17284 );
   nand U17955 ( n18180,n16030,n18192 );
   not U17956 ( n16030,n14610 );
   nand U17957 ( n14610,n18193,n18194 );
   nand U17958 ( n18194,n17289,n11768 );
   xor U17959 ( n11768,n18195,n18196 );
   xor U17960 ( n18196,si_26_,n18197 );
   nand U17961 ( n18193,n17294,p2_datao_reg_26_ );
   nor U17962 ( n17757,n17644,n17649 );
   nor U17963 ( n17649,n18198,n18199 );
   not U17964 ( n17644,n17647 );
   nand U17965 ( n17647,n18199,n18198 );
   nand U17966 ( n18198,n18200,n18201 );
   nand U17967 ( n18201,n17654,n14597 );
   nand U17968 ( n18200,n17655,n14360 );
   xor U17969 ( n18199,n17657,n18202 );
   nand U17970 ( n18202,n18203,n18204 );
   nand U17971 ( n18204,n17660,n14597 );
   nand U17972 ( n14597,n18205,n18206 );
   nand U17973 ( n18206,n17289,n11778 );
   xor U17974 ( n11778,n17669,n18207 );
   xor U17975 ( n18207,si_27_,n17668 );
   nand U17976 ( n17668,n18208,n18209 );
   nand U17977 ( n18209,n18210,n18211 );
   not U17978 ( n18211,si_26_ );
   or U17979 ( n18210,n18197,n18195 );
   nand U17980 ( n18208,n18195,n18197 );
   nand U17981 ( n18197,n18212,n18213 );
   nand U17982 ( n18213,n18214,n18215 );
   not U17983 ( n18215,si_25_ );
   or U17984 ( n18214,n18171,n18169 );
   nand U17985 ( n18212,n18169,n18171 );
   nand U17986 ( n18171,n18216,n18217 );
   nand U17987 ( n18217,n18218,n18219 );
   not U17988 ( n18219,si_24_ );
   or U17989 ( n18218,n17775,n17773 );
   nand U17990 ( n18216,n17773,n17775 );
   nand U17991 ( n17775,n18220,n18221 );
   nand U17992 ( n18221,n18222,n18223 );
   not U17993 ( n18223,si_23_ );
   or U17994 ( n18222,n18161,n18159 );
   nand U17995 ( n18220,n18159,n18161 );
   nand U17996 ( n18161,n18224,n18225 );
   nand U17997 ( n18225,n18226,n18227 );
   not U17998 ( n18227,si_22_ );
   or U17999 ( n18226,n18143,n18141 );
   nand U18000 ( n18224,n18141,n18143 );
   nand U18001 ( n18143,n18228,n18229 );
   nand U18002 ( n18229,n18230,n18231 );
   not U18003 ( n18231,si_21_ );
   or U18004 ( n18230,n17807,n17805 );
   nand U18005 ( n18228,n17805,n17807 );
   nand U18006 ( n17807,n18232,n18233 );
   nand U18007 ( n18233,n18234,n18235 );
   not U18008 ( n18235,si_20_ );
   or U18009 ( n18234,n18126,n18124 );
   nand U18010 ( n18232,n18124,n18126 );
   nand U18011 ( n18126,n18236,n18237 );
   nand U18012 ( n18237,n18238,n18239 );
   not U18013 ( n18239,si_19_ );
   or U18014 ( n18238,n18113,n18111 );
   nand U18015 ( n18236,n18111,n18113 );
   nand U18016 ( n18113,n18240,n18241 );
   nand U18017 ( n18241,n18242,n18243 );
   not U18018 ( n18243,si_18_ );
   or U18019 ( n18242,n18095,n18093 );
   nand U18020 ( n18240,n18093,n18095 );
   nand U18021 ( n18095,n18244,n18245 );
   nand U18022 ( n18245,n18246,n17843 );
   not U18023 ( n17843,si_17_ );
   or U18024 ( n18246,n17842,n17841 );
   nand U18025 ( n18244,n17841,n17842 );
   nand U18026 ( n17842,n18247,n18248 );
   nand U18027 ( n18248,n18249,n17867 );
   not U18028 ( n17867,si_16_ );
   or U18029 ( n18249,n17866,n17865 );
   nand U18030 ( n18247,n17865,n17866 );
   nand U18031 ( n17866,n18250,n18251 );
   nand U18032 ( n18251,n18252,n18080 );
   not U18033 ( n18080,si_15_ );
   nand U18034 ( n18252,n18079,n18081 );
   or U18035 ( n18250,n18081,n18079 );
   nand U18036 ( n18079,n18253,n18254 );
   nand U18037 ( n18254,n11808,p1_datao_reg_15_ );
   nand U18038 ( n18253,n11812,p2_datao_reg_15_ );
   nand U18039 ( n18081,n18255,n18256,n18257 );
   or U18040 ( n18257,n18058,n18258 );
   nand U18041 ( n18256,n18259,n18260 );
   or U18042 ( n18260,n18055,si_14_ );
   not U18043 ( n18055,n18258 );
   not U18044 ( n18259,n18059 );
   nand U18045 ( n18059,n18036,n18015,n17912,n17905 );
   nand U18046 ( n18015,n18261,n18262 );
   nand U18047 ( n18262,si_10_,n18263 );
   or U18048 ( n18263,n18001,n17999 );
   nand U18049 ( n18261,n17999,n18001 );
   nand U18050 ( n18001,n17973,n18264 );
   nand U18051 ( n18264,n17972,n17974 );
   nand U18052 ( n17974,n18265,n18266,n18267 );
   not U18053 ( n18267,si_9_ );
   nand U18054 ( n18266,n11808,p1_datao_reg_9_ );
   nand U18055 ( n18265,n11812,p2_datao_reg_9_ );
   nand U18056 ( n17972,n17960,n18268 );
   nand U18057 ( n18268,n17959,n17961 );
   nand U18058 ( n17961,n18269,n18270,n18271 );
   not U18059 ( n18271,si_8_ );
   nand U18060 ( n18270,n11808,p1_datao_reg_8_ );
   nand U18061 ( n18269,n11812,p2_datao_reg_8_ );
   nand U18062 ( n17959,n18272,n18273 );
   nand U18063 ( n18273,n18274,n18275 );
   nand U18064 ( n17960,n18276,n18277,si_8_ );
   or U18065 ( n18277,n11808,p2_datao_reg_8_ );
   nand U18066 ( n18276,n11808,n13990 );
   not U18067 ( n13990,p1_datao_reg_8_ );
   nand U18068 ( n17973,n18278,n18279,si_9_ );
   or U18069 ( n18279,n11808,p2_datao_reg_9_ );
   nand U18070 ( n18278,n11808,n13997 );
   not U18071 ( n13997,p1_datao_reg_9_ );
   and U18072 ( n17999,n18280,n18281 );
   or U18073 ( n18281,n11808,p2_datao_reg_10_ );
   or U18074 ( n18280,n11812,p1_datao_reg_10_ );
   not U18075 ( n18036,n18016 );
   nor U18076 ( n18016,n18282,si_11_ );
   nand U18077 ( n18255,si_14_,n18283 );
   nand U18078 ( n18283,n18258,n18058 );
   nand U18079 ( n18058,n17905,n18284 );
   nand U18080 ( n18284,n17904,n17909,n18285 );
   nand U18081 ( n18285,n18017,n17912 );
   nand U18082 ( n17912,n18286,n18287,n18288 );
   not U18083 ( n18288,si_12_ );
   nand U18084 ( n18287,n11808,p1_datao_reg_12_ );
   nand U18085 ( n18286,n11812,p2_datao_reg_12_ );
   not U18086 ( n18017,n18034 );
   nand U18087 ( n18034,si_11_,n18282 );
   nand U18088 ( n18282,n18289,n18290 );
   nand U18089 ( n18290,n11808,p1_datao_reg_11_ );
   nand U18090 ( n18289,n11812,p2_datao_reg_11_ );
   nand U18091 ( n17909,n18291,n18292,si_12_ );
   or U18092 ( n18292,n11808,p2_datao_reg_12_ );
   nand U18093 ( n18291,n11808,n14027 );
   not U18094 ( n14027,p1_datao_reg_12_ );
   nand U18095 ( n17904,si_13_,n17908 );
   or U18096 ( n17905,n17908,si_13_ );
   and U18097 ( n17908,n18293,n18294 );
   or U18098 ( n18294,n11808,p2_datao_reg_13_ );
   or U18099 ( n18293,n11812,p1_datao_reg_13_ );
   nand U18100 ( n18258,n18295,n18296 );
   or U18101 ( n18296,n11808,p2_datao_reg_14_ );
   or U18102 ( n18295,n11812,p1_datao_reg_14_ );
   nand U18103 ( n17865,n18297,n18298 );
   or U18104 ( n18298,n11808,p2_datao_reg_16_ );
   nand U18105 ( n18297,n11808,n13923 );
   not U18106 ( n13923,p1_datao_reg_16_ );
   nand U18107 ( n17841,n18299,n18300 );
   or U18108 ( n18300,n11808,p2_datao_reg_17_ );
   nand U18109 ( n18299,n11808,n13911 );
   not U18110 ( n13911,p1_datao_reg_17_ );
   nand U18111 ( n18093,n18301,n18302 );
   or U18112 ( n18302,n11808,p2_datao_reg_18_ );
   nand U18113 ( n18301,n11808,n14065 );
   not U18114 ( n14065,p1_datao_reg_18_ );
   nand U18115 ( n18111,n18303,n18304 );
   or U18116 ( n18304,n11808,p2_datao_reg_19_ );
   nand U18117 ( n18303,n11808,n14080 );
   not U18118 ( n14080,p1_datao_reg_19_ );
   nand U18119 ( n18124,n18305,n18306 );
   or U18120 ( n18306,n11808,p2_datao_reg_20_ );
   nand U18121 ( n18305,n11808,n14083 );
   not U18122 ( n14083,p1_datao_reg_20_ );
   nand U18123 ( n17805,n18307,n18308 );
   or U18124 ( n18308,n11808,p2_datao_reg_21_ );
   nand U18125 ( n18307,n11808,n13878 );
   not U18126 ( n13878,p1_datao_reg_21_ );
   nand U18127 ( n18141,n18309,n18310 );
   or U18128 ( n18310,n11808,p2_datao_reg_22_ );
   nand U18129 ( n18309,n11808,n14086 );
   not U18130 ( n14086,p1_datao_reg_22_ );
   nand U18131 ( n18159,n18311,n18312 );
   or U18132 ( n18312,n11808,p2_datao_reg_23_ );
   nand U18133 ( n18311,n11808,n13853 );
   not U18134 ( n13853,p1_datao_reg_23_ );
   nand U18135 ( n17773,n18313,n18314 );
   or U18136 ( n18314,n11808,p2_datao_reg_24_ );
   nand U18137 ( n18313,n11808,n14123 );
   not U18138 ( n14123,p1_datao_reg_24_ );
   nand U18139 ( n18169,n18315,n18316 );
   or U18140 ( n18316,n11808,p2_datao_reg_25_ );
   nand U18141 ( n18315,n11808,n14115 );
   not U18142 ( n14115,p1_datao_reg_25_ );
   nand U18143 ( n18195,n18317,n18318 );
   or U18144 ( n18318,n11808,p2_datao_reg_26_ );
   nand U18145 ( n18317,n11808,n14098 );
   not U18146 ( n14098,p1_datao_reg_26_ );
   nand U18147 ( n17669,n18319,n18320 );
   or U18148 ( n18320,n11808,p2_datao_reg_27_ );
   nand U18149 ( n18319,n11808,n14128 );
   not U18150 ( n14128,p1_datao_reg_27_ );
   nand U18151 ( n18205,n17294,p2_datao_reg_27_ );
   nand U18152 ( n18203,n17654,n14360 );
   nand U18153 ( n14360,n18321,n18322,n18323,n18324 );
   nand U18154 ( n18324,n17676,n16074 );
   nand U18155 ( n18323,p1_reg0_reg_27_,n17285 );
   nand U18156 ( n18322,p1_reg1_reg_27_,n17286 );
   nand U18157 ( n18321,p1_reg2_reg_27_,n17284 );
   nand U18158 ( n17744,n16074,n17375 );
   nand U18159 ( n17375,n18325,n18326 );
   nand U18160 ( n18325,n18327,p1_state_reg );
   xor U18161 ( n16074,n17677,n17678 );
   or U18162 ( n17678,n17365,n18191 );
   nand U18163 ( n18191,p1_reg3_reg_25_,n17781 );
   nor U18164 ( n17781,n17724,n18149,n17513 );
   not U18165 ( n17513,p1_reg3_reg_24_ );
   not U18166 ( n18149,n17783 );
   nor U18167 ( n17783,n17596,n17812,n17438 );
   not U18168 ( n17438,p1_reg3_reg_22_ );
   nand U18169 ( n17812,p1_reg3_reg_19_,n18133,p1_reg3_reg_20_ );
   not U18170 ( n18133,n18101 );
   nand U18171 ( n18101,p1_reg3_reg_17_,n17848,p1_reg3_reg_18_ );
   nor U18172 ( n17848,n17348,n17874,n17554 );
   not U18173 ( n17554,p1_reg3_reg_16_ );
   nand U18174 ( n17874,p1_reg3_reg_13_,n18066,p1_reg3_reg_14_ );
   not U18175 ( n18066,n17918 );
   nand U18176 ( n17918,p1_reg3_reg_11_,n18043,p1_reg3_reg_12_ );
   not U18177 ( n18043,n17988 );
   nand U18178 ( n17988,p1_reg3_reg_10_,n17979,p1_reg3_reg_9_ );
   not U18179 ( n17348,p1_reg3_reg_15_ );
   not U18180 ( n17596,p1_reg3_reg_21_ );
   not U18181 ( n17724,p1_reg3_reg_23_ );
   not U18182 ( n17365,p1_reg3_reg_26_ );
   not U18183 ( n17677,p1_reg3_reg_27_ );
   nor U18184 ( n18331,n18332,n18333,n18334 );
   nor U18185 ( n18334,n14883,n17364 );
   not U18186 ( n17364,n17356 );
   nor U18187 ( n17356,n18335,n16272,n18336 );
   not U18188 ( n14883,n14423 );
   nor U18189 ( n18333,n14834,n17346 );
   nor U18190 ( n17417,n16188,n18335,n18336 );
   not U18191 ( n14834,n14417 );
   nand U18192 ( n14417,n18337,n18338,n18339,n18340 );
   nand U18193 ( n18340,n17622,n17676 );
   nor U18194 ( n17622,n18341,n17979 );
   nor U18195 ( n17979,n18342,n18343,n17623 );
   and U18196 ( n18341,n17623,n18344 );
   or U18197 ( n18344,n18342,n18343 );
   not U18198 ( n17623,p1_reg3_reg_8_ );
   nand U18199 ( n18339,p1_reg0_reg_8_,n17285 );
   nand U18200 ( n18338,p1_reg1_reg_8_,n17286 );
   nand U18201 ( n18337,p1_reg2_reg_8_,n17284 );
   nor U18202 ( n18332,p1_state_reg,n18342 );
   nand U18203 ( n18330,n15453,n17347 );
   nand U18204 ( n17347,n18345,n18326 );
   nand U18205 ( n18326,n18346,p1_state_reg );
   nand U18206 ( n18346,n16821,n18347,n16282,n17336 );
   nand U18207 ( n16282,n16187,n14965 );
   nand U18208 ( n18347,n18348,n18335 );
   nand U18209 ( n18345,n18327,n14541 );
   and U18210 ( n18327,n18335,n18349 );
   nand U18211 ( n18349,n18336,n18350 );
   nand U18212 ( n18336,n14966,n14541,n18351 );
   nand U18213 ( n18329,n18352,n18353,n17366 );
   not U18214 ( n17366,n17351 );
   nand U18215 ( n17351,n14541,n18348,n18354 );
   nand U18216 ( n18348,n18355,n18356,n18357 );
   nor U18217 ( n18357,n16276,n15510,n15514 );
   not U18218 ( n15514,n15420 );
   nand U18219 ( n15420,n18351,n14968 );
   not U18220 ( n18351,n17338 );
   not U18221 ( n15510,n15426 );
   nand U18222 ( n15426,n14967,n14966,n16816 );
   nor U18223 ( n16276,n14607,n16288 );
   nand U18224 ( n14607,n18358,n14970 );
   or U18225 ( n18356,n17135,n16814 );
   nor U18226 ( n16814,n15345,n15870 );
   not U18227 ( n15870,n15437 );
   nand U18228 ( n15345,n15427,n15421 );
   nand U18229 ( n15421,n18360,n14966,n16288 );
   nand U18230 ( n15427,n16288,n14966,n14970 );
   or U18231 ( n18355,n14966,n16813 );
   nor U18232 ( n16813,n15346,n15014,n16256 );
   not U18233 ( n16256,n18361 );
   not U18234 ( n15014,n15320 );
   not U18235 ( n15346,n15013 );
   nand U18236 ( n18353,n17944,n18362 );
   nand U18237 ( n18362,n17945,n17943 );
   not U18238 ( n17944,n18363 );
   nand U18239 ( n18352,n17945,n17943,n18363 );
   nand U18240 ( n18363,n18364,n18365 );
   nand U18241 ( n18365,n17388,n18366 );
   nand U18242 ( n18366,n17389,n17387 );
   and U18243 ( n17388,n18367,n18368 );
   nand U18244 ( n18368,n17543,n18369 );
   nand U18245 ( n18369,n18370,n17544 );
   xor U18246 ( n17543,n17479,n18371 );
   nand U18247 ( n18371,n18372,n18373 );
   nand U18248 ( n18373,n17660,n15392 );
   nand U18249 ( n18372,n17654,n14426 );
   or U18250 ( n18367,n17544,n18370 );
   not U18251 ( n18370,n17545 );
   nand U18252 ( n17545,n18374,n18375 );
   nand U18253 ( n18375,n18376,n18377 );
   nand U18254 ( n18377,n17503,n17502 );
   not U18255 ( n18376,n17504 );
   nand U18256 ( n17504,n18378,n18379 );
   nand U18257 ( n18379,n17654,n15376 );
   nand U18258 ( n18378,n17655,n14429 );
   or U18259 ( n18374,n17502,n17503 );
   nor U18260 ( n17503,n18380,n17700 );
   nor U18261 ( n17700,n18381,n18382 );
   nor U18262 ( n18380,n17702,n17701 );
   and U18263 ( n17701,n18381,n18382 );
   nand U18264 ( n18382,n18383,n18384 );
   nand U18265 ( n18384,n17654,n15338 );
   nand U18266 ( n18383,n17655,n14432 );
   xor U18267 ( n18381,n17657,n18385 );
   nand U18268 ( n18385,n18386,n18387 );
   nand U18269 ( n18387,n17660,n15338 );
   nand U18270 ( n15338,n18388,n18389,n18390 );
   nand U18271 ( n18390,n17294,p2_datao_reg_3_ );
   nand U18272 ( n18389,n16734,n16273 );
   not U18273 ( n16734,n16722 );
   nand U18274 ( n16722,n18391,n18392 );
   or U18275 ( n18392,p1_ir_reg_31_,p1_ir_reg_3_ );
   or U18276 ( n18391,n15049,n15241 );
   xor U18277 ( n15049,p1_ir_reg_3_,n15044 );
   nand U18278 ( n18388,n17289,n11578 );
   xor U18279 ( n11578,n18393,n18394 );
   xor U18280 ( n18393,n18395,n18396 );
   nand U18281 ( n18395,n18397,n18398 );
   nand U18282 ( n18398,n18399,n18400 );
   nand U18283 ( n18386,n17654,n14432 );
   nand U18284 ( n14432,n18401,n18402,n18403,n18404 );
   nand U18285 ( n18404,p1_reg0_reg_3_,n17285 );
   nand U18286 ( n18403,p1_reg1_reg_3_,n17286 );
   nand U18287 ( n18402,p1_reg2_reg_3_,n17284 );
   nand U18288 ( n18401,n17676,n15350 );
   nand U18289 ( n17702,n18405,n18406 );
   nand U18290 ( n18406,n17412,n18407 );
   nand U18291 ( n18407,n18408,n17415 );
   xor U18292 ( n17412,n17657,n18409 );
   nand U18293 ( n18409,n18410,n18411 );
   nand U18294 ( n18411,n17660,n15306 );
   nand U18295 ( n18410,n17654,n14435 );
   or U18296 ( n18405,n17415,n18408 );
   not U18297 ( n18408,n17414 );
   nand U18298 ( n17414,n18412,n18413 );
   nand U18299 ( n18413,n17654,n15306 );
   nand U18300 ( n15306,n18414,n18415,n18416 );
   nand U18301 ( n18416,n17294,p2_datao_reg_2_ );
   nand U18302 ( n18415,n16762,n16273 );
   not U18303 ( n16762,n16779 );
   nand U18304 ( n16779,n18417,n18418 );
   or U18305 ( n18418,p1_ir_reg_2_,p1_ir_reg_31_ );
   nand U18306 ( n18417,p1_ir_reg_31_,n18419 );
   nand U18307 ( n18419,n15043,n15044 );
   nand U18308 ( n15043,p1_ir_reg_2_,n18420 );
   nand U18309 ( n18420,n16772,n18421 );
   nand U18310 ( n18414,n17289,n11568 );
   nand U18311 ( n11568,n18422,n18423,n18424 );
   nand U18312 ( n18424,n18425,n18426 );
   xor U18313 ( n18425,n18427,n18400 );
   or U18314 ( n18423,n18426,n18427,n18400 );
   nand U18315 ( n18422,n18428,n18400 );
   not U18316 ( n18428,n18397 );
   nand U18317 ( n18412,n17655,n14435 );
   nand U18318 ( n14435,n18429,n18430,n18431,n18432 );
   nand U18319 ( n18432,p1_reg0_reg_2_,n17285 );
   nand U18320 ( n18431,p1_reg1_reg_2_,n17286 );
   nand U18321 ( n18430,p1_reg2_reg_2_,n17284 );
   nand U18322 ( n18429,p1_reg3_reg_2_,n17676 );
   nand U18323 ( n17415,n18433,n18434 );
   nand U18324 ( n18434,n17612,n18435 );
   or U18325 ( n18435,n17614,n17613 );
   xor U18326 ( n17612,n17479,n18436 );
   nand U18327 ( n18436,n18437,n18438 );
   nand U18328 ( n18438,n17660,n15281 );
   nand U18329 ( n18437,n17654,n14438 );
   nand U18330 ( n18433,n17613,n17614 );
   nand U18331 ( n17614,n18439,n18440 );
   nand U18332 ( n18440,n17479,n18441 );
   nand U18333 ( n18441,n17477,n17480 );
   or U18334 ( n18439,n17477,n17480 );
   nand U18335 ( n17480,n18442,n18443,n18444 );
   nand U18336 ( n18444,p1_ir_reg_0_,n16820 );
   nand U18337 ( n18443,n17655,n14441 );
   nand U18338 ( n18442,n17654,n14956 );
   xor U18339 ( n17477,n17657,n18445 );
   nand U18340 ( n18445,n18446,n18447,n18448 );
   nand U18341 ( n18448,p1_reg1_reg_0_,n16820 );
   nand U18342 ( n18447,n17654,n14441 );
   nand U18343 ( n14441,n18449,n18450,n18451,n18452 );
   nand U18344 ( n18452,p1_reg0_reg_0_,n17285 );
   nand U18345 ( n18451,p1_reg1_reg_0_,n17286 );
   nand U18346 ( n18450,p1_reg2_reg_0_,n17284 );
   nand U18347 ( n18449,p1_reg3_reg_0_,n17676 );
   nand U18348 ( n18446,n17660,n14956 );
   nand U18349 ( n14956,n18453,n18454,n18455 );
   nand U18350 ( n18455,p1_ir_reg_0_,n16273 );
   nand U18351 ( n18454,n17289,n11551 );
   and U18352 ( n11551,n18456,n18457 );
   nand U18353 ( n18456,n18458,n18459 );
   nand U18354 ( n18453,n17294,p2_datao_reg_0_ );
   and U18355 ( n17613,n18460,n18461 );
   nand U18356 ( n18461,n17654,n15281 );
   nand U18357 ( n15281,n18462,n18463,n18464 );
   nand U18358 ( n18464,n17294,p2_datao_reg_1_ );
   nand U18359 ( n18463,n16788,n16273 );
   not U18360 ( n16788,n16797 );
   nand U18361 ( n16797,n18465,n18466 );
   nand U18362 ( n18466,n18421,n15241 );
   or U18363 ( n18465,n15038,n15241 );
   xor U18364 ( n15038,n16772,n18421 );
   not U18365 ( n18421,p1_ir_reg_1_ );
   not U18366 ( n16772,p1_ir_reg_0_ );
   nand U18367 ( n18462,n17289,n11561 );
   xor U18368 ( n11561,n18467,n18468 );
   xor U18369 ( n18467,si_1_,n18457 );
   nand U18370 ( n18460,n17655,n14438 );
   nand U18371 ( n14438,n18469,n18470,n18471,n18472 );
   nand U18372 ( n18472,p1_reg0_reg_1_,n17285 );
   nand U18373 ( n18471,p1_reg1_reg_1_,n17286 );
   nand U18374 ( n18470,p1_reg2_reg_1_,n17284 );
   nand U18375 ( n18469,p1_reg3_reg_1_,n17676 );
   xor U18376 ( n17502,n17657,n18473 );
   nand U18377 ( n18473,n18474,n18475 );
   nand U18378 ( n18475,n17660,n15376 );
   nand U18379 ( n15376,n18476,n18477,n18478 );
   nand U18380 ( n18478,n17294,p2_datao_reg_4_ );
   nand U18381 ( n18477,n17289,n11585 );
   xor U18382 ( n11585,n18479,n18480 );
   and U18383 ( n18479,n18481,n18482 );
   nand U18384 ( n18476,n16717,n16273 );
   not U18385 ( n16717,n16708 );
   nand U18386 ( n16708,n18483,n18484 );
   or U18387 ( n18484,p1_ir_reg_31_,p1_ir_reg_4_ );
   nand U18388 ( n18483,p1_ir_reg_31_,n18485 );
   nand U18389 ( n18485,n15055,n15054 );
   nand U18390 ( n15054,p1_ir_reg_4_,n18486 );
   nand U18391 ( n18474,n17654,n14429 );
   nand U18392 ( n14429,n18487,n18488,n18489,n18490 );
   nand U18393 ( n18490,n17505,n17676 );
   nor U18394 ( n17505,n18491,n18492 );
   nor U18395 ( n18491,p1_reg3_reg_4_,p1_reg3_reg_3_ );
   nand U18396 ( n18489,p1_reg0_reg_4_,n17285 );
   nand U18397 ( n18488,p1_reg1_reg_4_,n17286 );
   nand U18398 ( n18487,p1_reg2_reg_4_,n17284 );
   nand U18399 ( n17544,n18493,n18494 );
   nand U18400 ( n18494,n17654,n15392 );
   nand U18401 ( n15392,n18495,n18496,n18497 );
   nand U18402 ( n18497,n17294,p2_datao_reg_5_ );
   nand U18403 ( n18496,n17289,n11594 );
   xor U18404 ( n11594,n18498,n18499 );
   and U18405 ( n18498,n18500,n18501 );
   nand U18406 ( n18495,n16665,n16273 );
   not U18407 ( n16665,n16686 );
   nand U18408 ( n16686,n18502,n18503,n18504 );
   nand U18409 ( n18503,n15241,n15064 );
   nand U18410 ( n18502,p1_ir_reg_31_,n15055,p1_ir_reg_5_ );
   not U18411 ( n15055,n15063 );
   nand U18412 ( n18493,n17655,n14426 );
   nand U18413 ( n14426,n18505,n18506,n18507,n18508 );
   nand U18414 ( n18508,n17676,n15402 );
   xor U18415 ( n15402,p1_reg3_reg_5_,n18492 );
   nand U18416 ( n18507,p1_reg0_reg_5_,n17285 );
   nand U18417 ( n18506,p1_reg1_reg_5_,n17286 );
   nand U18418 ( n18505,p1_reg2_reg_5_,n17284 );
   or U18419 ( n18364,n17387,n17389 );
   and U18420 ( n17389,n18509,n18510 );
   nand U18421 ( n18510,n17654,n14873 );
   nand U18422 ( n18509,n17655,n14423 );
   xor U18423 ( n17387,n17479,n18511 );
   nand U18424 ( n18511,n18512,n18513 );
   nand U18425 ( n18513,n17660,n14873 );
   nand U18426 ( n14873,n18514,n18515,n18516 );
   nand U18427 ( n18516,n17294,p2_datao_reg_6_ );
   nand U18428 ( n18515,n16652,n16273 );
   not U18429 ( n16652,n16653 );
   nand U18430 ( n16653,n18517,n18518 );
   or U18431 ( n18518,p1_ir_reg_31_,p1_ir_reg_6_ );
   nand U18432 ( n18517,p1_ir_reg_31_,n18519 );
   nand U18433 ( n18519,n15069,n15070 );
   nand U18434 ( n15069,p1_ir_reg_6_,n18504 );
   nand U18435 ( n18514,n17289,n11601 );
   xor U18436 ( n11601,n18520,n18521 );
   xor U18437 ( n18520,n18522,si_6_ );
   nand U18438 ( n18512,n17654,n14423 );
   nand U18439 ( n14423,n18523,n18524,n18525,n18526 );
   nand U18440 ( n18526,p1_reg0_reg_6_,n17285 );
   nand U18441 ( n18525,p1_reg1_reg_6_,n17286 );
   nand U18442 ( n18524,p1_reg2_reg_6_,n17284 );
   nand U18443 ( n18523,n17384,n17676 );
   not U18444 ( n17384,n15412 );
   nand U18445 ( n15412,n18527,n18343 );
   nand U18446 ( n18527,n17383,n18528 );
   nand U18447 ( n18528,p1_reg3_reg_5_,n18492 );
   not U18448 ( n17383,p1_reg3_reg_6_ );
   nand U18449 ( n17943,n18529,n18530 );
   not U18450 ( n18530,n18531 );
   xor U18451 ( n18529,n17479,n18532 );
   nand U18452 ( n17945,n18533,n18531 );
   nand U18453 ( n18531,n18534,n18535 );
   nand U18454 ( n18535,n17655,n14420 );
   nand U18455 ( n18534,n17654,n14861 );
   xor U18456 ( n18533,n18532,n17657 );
   nand U18457 ( n18537,n16288,n14967 );
   nand U18458 ( n18536,n18360,n17135 );
   nand U18459 ( n18532,n18539,n18540 );
   nand U18460 ( n18540,n17654,n14420 );
   nand U18461 ( n14420,n18541,n18542,n18543,n18544 );
   nand U18462 ( n18544,n17676,n15453 );
   xor U18463 ( n15453,n18342,n18343 );
   nand U18464 ( n18343,p1_reg3_reg_5_,n18492,p1_reg3_reg_6_ );
   nor U18465 ( n18492,n16713,n15350 );
   not U18466 ( n15350,p1_reg3_reg_3_ );
   not U18467 ( n16713,p1_reg3_reg_4_ );
   not U18468 ( n18342,p1_reg3_reg_7_ );
   nand U18469 ( n18543,p1_reg0_reg_7_,n17285 );
   not U18470 ( n18545,n18547 );
   nand U18471 ( n18542,p1_reg1_reg_7_,n17286 );
   nand U18472 ( n18541,p1_reg2_reg_7_,n17284 );
   xor U18473 ( n18546,n15241,n15237 );
   not U18474 ( n15237,p1_ir_reg_30_ );
   xor U18475 ( n18547,p1_ir_reg_31_,n15228 );
   not U18476 ( n15228,p1_ir_reg_29_ );
   nand U18477 ( n18185,n18548,n17336 );
   nand U18478 ( n18548,n17338,n18361 );
   nand U18479 ( n18361,n16288,n17135,n14970 );
   nand U18480 ( n17338,n16816,n17135 );
   not U18481 ( n16816,n14965 );
   nand U18482 ( n14965,n14970,n16316 );
   nand U18483 ( n18539,n17660,n14861 );
   nand U18484 ( n18538,n18358,n17336 );
   nand U18485 ( n18192,n18549,n17336 );
   not U18486 ( n17336,n16820 );
   nand U18487 ( n18549,n18550,n15320,n14968 );
   nand U18488 ( n18328,n17349,n14861 );
   nand U18489 ( n14861,n18551,n18552,n18553 );
   nand U18490 ( n18553,n17294,p2_datao_reg_7_ );
   nand U18491 ( n18552,n16604,n16273 );
   not U18492 ( n16604,n16633 );
   nand U18493 ( n16633,n18554,n18555,n17957 );
   nand U18494 ( n18555,n15241,n15078 );
   nand U18495 ( n18554,p1_ir_reg_31_,n15070,p1_ir_reg_7_ );
   not U18496 ( n15070,n15077 );
   nand U18497 ( n18551,n17289,n11610 );
   xor U18498 ( n11610,n18556,n18274 );
   nand U18499 ( n18274,n18557,n18558 );
   nand U18500 ( n18558,si_6_,n18559 );
   nand U18501 ( n18559,n18522,n18521 );
   or U18502 ( n18557,n18521,n18522 );
   and U18503 ( n18522,n18501,n18560 );
   nand U18504 ( n18560,n18499,n18500 );
   nand U18505 ( n18500,n18561,n18562,n18563 );
   not U18506 ( n18563,si_5_ );
   nand U18507 ( n18562,n11808,p1_datao_reg_5_ );
   nand U18508 ( n18561,n11812,p2_datao_reg_5_ );
   nand U18509 ( n18499,n18481,n18564 );
   nand U18510 ( n18564,n18480,n18482 );
   or U18511 ( n18482,n18565,si_4_ );
   nand U18512 ( n18480,n18566,n18567,n18568 );
   or U18513 ( n18568,n18397,n18394 );
   nand U18514 ( n18567,n18569,n18400,n18399 );
   nand U18515 ( n18399,n18570,n18426 );
   not U18516 ( n18426,si_2_ );
   not U18517 ( n18570,n18427 );
   nand U18518 ( n18400,n18571,n18572 );
   nand U18519 ( n18572,si_1_,n18573 );
   nand U18520 ( n18573,n18468,n18457 );
   or U18521 ( n18571,n18457,n18468 );
   nand U18522 ( n18468,n18574,n18575 );
   or U18523 ( n18575,n11808,p2_datao_reg_1_ );
   or U18524 ( n18574,n11812,p1_datao_reg_1_ );
   or U18525 ( n18457,n18459,n18458 );
   and U18526 ( n18458,n18576,n18577 );
   nand U18527 ( n18577,n11808,p1_datao_reg_0_ );
   nand U18528 ( n18576,n11812,p2_datao_reg_0_ );
   not U18529 ( n18459,si_0_ );
   nand U18530 ( n18569,n18394,n18396 );
   not U18531 ( n18396,si_3_ );
   nand U18532 ( n18566,si_3_,n18578 );
   nand U18533 ( n18578,n18394,n18397 );
   nand U18534 ( n18397,si_2_,n18427 );
   nand U18535 ( n18427,n18579,n18580 );
   nand U18536 ( n18580,n11808,p1_datao_reg_2_ );
   nand U18537 ( n18579,n11812,p2_datao_reg_2_ );
   nand U18538 ( n18394,n18581,n18582 );
   or U18539 ( n18582,n11808,p2_datao_reg_3_ );
   or U18540 ( n18581,n11812,p1_datao_reg_3_ );
   nand U18541 ( n18481,si_4_,n18565 );
   nand U18542 ( n18565,n18583,n18584 );
   nand U18543 ( n18584,n11808,p1_datao_reg_4_ );
   nand U18544 ( n18583,n11812,p2_datao_reg_4_ );
   nand U18545 ( n18501,n18585,n18586,si_5_ );
   or U18546 ( n18586,n11808,p2_datao_reg_5_ );
   nand U18547 ( n18585,n11808,n14262 );
   not U18548 ( n14262,p1_datao_reg_5_ );
   nand U18549 ( n18521,n18587,n18588 );
   or U18550 ( n18588,n11808,p2_datao_reg_6_ );
   or U18551 ( n18587,n11812,p1_datao_reg_6_ );
   and U18552 ( n18556,n18272,n18275 );
   or U18553 ( n18275,n18589,si_7_ );
   nand U18554 ( n18272,si_7_,n18589 );
   nand U18555 ( n18589,n18590,n18591 );
   nand U18556 ( n18591,n11808,p1_datao_reg_7_ );
   nand U18557 ( n18590,n11812,p2_datao_reg_7_ );
   or U18558 ( n18594,p1_addr_reg_19_,p1_rd_reg,p2_addr_reg_19_ );
   nand U18559 ( n18593,p1_addr_reg_19_,n10452,p2_addr_reg_19_ );
   not U18560 ( n10452,p2_rd_reg );
   not U18561 ( n17349,n17416 );
   nand U18562 ( n17416,n18595,n14541 );
   not U18563 ( n16817,n16821 );
   nand U18564 ( n18595,n16279,n18596 );
   nand U18565 ( n18596,n18354,n16277 );
   not U18566 ( n16277,n18350 );
   nand U18567 ( n18350,n18360,n14550 );
   nand U18568 ( n14550,n18597,n18598 );
   nand U18569 ( n18598,n18359,n18358 );
   nor U18570 ( n18358,n17135,n14966 );
   not U18571 ( n18359,n18550 );
   nand U18572 ( n18550,n16316,n18360 );
   not U18573 ( n16316,n16288 );
   nand U18574 ( n18597,n14967,n16884 );
   not U18575 ( n18354,n18335 );
   nand U18576 ( n18335,n14540,n14962,n16281 );
   not U18577 ( n16281,n14961 );
   nand U18578 ( n14961,n14975,n18599 );
   or U18579 ( n18599,n15252,p1_d_reg_1_ );
   nand U18580 ( n14975,n18600,n18601 );
   and U18581 ( n14962,n18602,n18603,n18604,n18605 );
   nor U18582 ( n18605,n18606,n18607,n18608,n18609 );
   nor U18583 ( n18609,n15252,n15243 );
   not U18584 ( n15243,p1_d_reg_6_ );
   nor U18585 ( n18608,n15252,n15245 );
   not U18586 ( n15245,p1_d_reg_13_ );
   nor U18587 ( n18607,n15252,n15247 );
   not U18588 ( n15247,p1_d_reg_17_ );
   nor U18589 ( n18606,n18610,n15252 );
   nor U18590 ( n18610,p1_d_reg_22_,p1_d_reg_24_,p1_d_reg_23_ );
   nor U18591 ( n18604,n18611,n18612,n18613,n18614 );
   nor U18592 ( n18614,n15252,n15249 );
   not U18593 ( n15249,p1_d_reg_19_ );
   nor U18594 ( n18613,n15252,n15246 );
   not U18595 ( n15246,p1_d_reg_16_ );
   nor U18596 ( n18612,n18615,n15252 );
   nor U18597 ( n18615,p1_d_reg_7_,p1_d_reg_9_,p1_d_reg_8_ );
   nor U18598 ( n18611,n15252,n15244 );
   not U18599 ( n15244,p1_d_reg_10_ );
   nor U18600 ( n18603,n18616,n18617,n18618,n18619 );
   nor U18601 ( n18619,n15252,n15251 );
   not U18602 ( n15251,p1_d_reg_29_ );
   nor U18603 ( n18618,n15252,n15242 );
   not U18604 ( n15242,p1_d_reg_2_ );
   nor U18605 ( n18617,n15252,n15250 );
   not U18606 ( n15250,p1_d_reg_27_ );
   nor U18607 ( n18616,n15252,n15248 );
   not U18608 ( n15248,p1_d_reg_18_ );
   nor U18609 ( n18602,n18620,n18621,n18622,n18623 );
   nor U18610 ( n18623,n18624,n15252 );
   nor U18611 ( n18624,p1_d_reg_5_,p1_d_reg_4_,p1_d_reg_3_,p1_d_reg_30_ );
   nor U18612 ( n18622,n18625,n15252 );
   nor U18613 ( n18625,p1_d_reg_20_,p1_d_reg_26_,p1_d_reg_25_ );
   nor U18614 ( n18621,n18626,n15252 );
   nor U18615 ( n18626,p1_d_reg_15_,p1_d_reg_14_,p1_d_reg_12_,p1_d_reg_11_ );
   nor U18616 ( n18620,n18627,n15252 );
   nor U18617 ( n18627,p1_d_reg_21_,p1_d_reg_31_,p1_d_reg_28_ );
   not U18618 ( n14540,n14959 );
   nand U18619 ( n14959,n14978,n18628 );
   or U18620 ( n18628,n15252,p1_d_reg_0_ );
   nand U18621 ( n18630,n18632,n16271 );
   not U18622 ( n16271,p1_b_reg );
   nand U18623 ( n18629,n18633,n18601,p1_b_reg );
   nand U18624 ( n14978,n18600,n18633 );
   nand U18625 ( n16279,n14682,n14967 );
   not U18626 ( n14682,n14568 );
   nand U18627 ( n18635,p1_ir_reg_19_,n15241 );
   nand U18628 ( n18634,n15157,n15158,p1_ir_reg_31_ );
   nand U18629 ( n15157,p1_ir_reg_19_,n18092 );
   not U18630 ( n14968,n14966 );
   not U18631 ( n14970,n18360 );
   nand U18632 ( n18360,n18636,n18637 );
   nand U18633 ( n18637,p1_ir_reg_20_,n15241 );
   nand U18634 ( n18636,n15163,n15164,p1_ir_reg_31_ );
   nand U18635 ( n15163,p1_ir_reg_20_,n15158 );
   nor U18636 ( n16820,n18601,n18633,n18600 );
   not U18637 ( n18600,n18631 );
   nand U18638 ( n18631,n18639,n18640 );
   nand U18639 ( n18640,p1_ir_reg_26_,n15241 );
   nand U18640 ( n18639,n15205,n15206,p1_ir_reg_31_ );
   nand U18641 ( n15205,p1_ir_reg_26_,n18641 );
   nand U18642 ( n18641,n15199,n15200 );
   not U18643 ( n15200,p1_ir_reg_25_ );
   not U18644 ( n18633,n18632 );
   nand U18645 ( n18632,n18642,n18643 );
   nand U18646 ( n18643,p1_ir_reg_24_,n15241 );
   nand U18647 ( n18642,n15191,n15192,p1_ir_reg_31_ );
   nand U18648 ( n15191,p1_ir_reg_24_,n18644 );
   nand U18649 ( n18644,n15185,n15186 );
   xor U18650 ( n18601,p1_ir_reg_25_,n18645 );
   nand U18651 ( n18645,p1_ir_reg_31_,n15192 );
   nand U18652 ( n18638,n18646,p1_state_reg );
   nand U18653 ( n18646,n18647,n18592 );
   nand U18654 ( n18592,n16768,n16272 );
   not U18655 ( n16272,n16188 );
   nand U18656 ( n16188,n18648,n18649 );
   nand U18657 ( n18649,p1_ir_reg_28_,n15241 );
   nand U18658 ( n18648,n15219,n15220,p1_ir_reg_31_ );
   not U18659 ( n15220,n15227 );
   nor U18660 ( n15227,p1_ir_reg_27_,p1_ir_reg_28_,n15206 );
   not U18661 ( n15206,n15213 );
   nand U18662 ( n15219,p1_ir_reg_28_,n18650 );
   nand U18663 ( n18650,n15213,n15214 );
   xor U18664 ( n16768,n18651,n15214 );
   not U18665 ( n15214,p1_ir_reg_27_ );
   nor U18666 ( n18651,n15213,n15241 );
   nor U18667 ( n15213,p1_ir_reg_25_,p1_ir_reg_26_,n15192 );
   not U18668 ( n15192,n15199 );
   nor U18669 ( n15199,p1_ir_reg_23_,p1_ir_reg_24_,n15178 );
   nand U18670 ( n18647,n16187,n16821 );
   xor U18671 ( n16821,n18652,n15186 );
   not U18672 ( n15186,p1_ir_reg_23_ );
   nor U18673 ( n18652,n15185,n15241 );
   not U18674 ( n16187,n17168 );
   nand U18675 ( n17168,n14966,n17135 );
   not U18676 ( n17135,n14967 );
   xor U18677 ( n14967,p1_ir_reg_21_,n18653 );
   nand U18678 ( n18653,p1_ir_reg_31_,n15164 );
   nand U18679 ( n14966,n18654,n18655 );
   nand U18680 ( n18655,p1_ir_reg_22_,n15241 );
   nand U18681 ( n18654,n15177,n15178,p1_ir_reg_31_ );
   not U18682 ( n15178,n15185 );
   nor U18683 ( n15185,p1_ir_reg_21_,p1_ir_reg_22_,n15164 );
   not U18684 ( n15164,n15171 );
   nand U18685 ( n15177,p1_ir_reg_22_,n18656 );
   nand U18686 ( n18656,n15171,n15172 );
   not U18687 ( n15172,p1_ir_reg_21_ );
   nor U18688 ( n15171,n15158,p1_ir_reg_20_ );
   or U18689 ( n15158,n18092,p1_ir_reg_19_ );
   nand U18690 ( n18092,n15150,n15152 );
   not U18691 ( n15152,p1_ir_reg_18_ );
   not U18692 ( n15150,n15151 );
   nand U18693 ( n15151,n15142,n15143 );
   not U18694 ( n15143,p1_ir_reg_17_ );
   nor U18695 ( n15142,n17863,p1_ir_reg_16_ );
   nand U18696 ( n17863,n15127,n15129 );
   not U18697 ( n15129,p1_ir_reg_15_ );
   nor U18698 ( n15127,n17899,p1_ir_reg_14_ );
   nand U18699 ( n17899,n15113,n15114 );
   not U18700 ( n15114,p1_ir_reg_13_ );
   nor U18701 ( n15113,p1_ir_reg_11_,p1_ir_reg_12_,n17995 );
   not U18702 ( n17995,n18013 );
   nor U18703 ( n18013,p1_ir_reg_10_,p1_ir_reg_9_,n15084 );
   not U18704 ( n15084,n17998 );
   nor U18705 ( n17998,n17957,p1_ir_reg_8_ );
   nand U18706 ( n17957,n15077,n15078 );
   not U18707 ( n15078,p1_ir_reg_7_ );
   nor U18708 ( n15077,n18504,p1_ir_reg_6_ );
   nand U18709 ( n18504,n15063,n15064 );
   not U18710 ( n15064,p1_ir_reg_5_ );
   nor U18711 ( n15063,n18486,p1_ir_reg_4_ );
   or U18712 ( n18486,n15044,p1_ir_reg_3_ );
   or U18713 ( n15044,p1_ir_reg_1_,p1_ir_reg_2_,p1_ir_reg_0_ );
   xor U18714 ( n18657,p1_addr_reg_10_,n13043 );
   xor U18715 ( n18659,p1_addr_reg_11_,n18661 );
   xor U18716 ( n18662,p1_addr_reg_12_,n18664 );
   xor U18717 ( n18665,p1_addr_reg_13_,n18667 );
   xor U18718 ( n18668,p1_addr_reg_14_,n18670 );
   xor U18719 ( n18671,p1_addr_reg_15_,n12844 );
   xor U18720 ( n18673,p1_addr_reg_16_,n18675 );
   xor U18721 ( n18676,p1_addr_reg_17_,n18678 );
   xor U18722 ( n18679,n18681,p2_addr_reg_18_ );
   xor U18723 ( n18682,p1_addr_reg_2_,n18684 );
   xor U18724 ( n18685,p1_addr_reg_3_,n18687 );
   xor U18725 ( n18688,p1_addr_reg_4_,n18690 );
   xor U18726 ( n18691,p1_addr_reg_5_,n18693 );
   xor U18727 ( n18694,p1_addr_reg_6_,n13196 );
   xor U18728 ( n18698,p1_addr_reg_7_,n13161 );
   xor U18729 ( n18700,p1_addr_reg_8_,n13117 );
   xor U18730 ( n18702,p1_addr_reg_9_,n18704 );
   nand U18731 ( n18706,n18707,n18708 );
   nand U18732 ( n18708,p2_addr_reg_18_,n18709 );
   nand U18733 ( n18709,n18681,n18680 );
   or U18734 ( n18707,n18680,n18681 );
   not U18735 ( n18681,p1_addr_reg_18_ );
   nand U18736 ( n18680,n18710,n18711 );
   nand U18737 ( n18711,n18712,n18678 );
   not U18738 ( n18678,p2_addr_reg_17_ );
   or U18739 ( n18712,n18677,n18713 );
   nand U18740 ( n18710,n18677,n18713 );
   not U18741 ( n18713,p1_addr_reg_17_ );
   nand U18742 ( n18677,n18714,n18715 );
   nand U18743 ( n18715,n18716,n18675 );
   not U18744 ( n18675,p2_addr_reg_16_ );
   or U18745 ( n18716,n18674,n18717 );
   nand U18746 ( n18714,n18674,n18717 );
   not U18747 ( n18717,p1_addr_reg_16_ );
   nand U18748 ( n18674,n18718,n18719 );
   nand U18749 ( n18719,n18720,n12844 );
   not U18750 ( n12844,p2_addr_reg_15_ );
   or U18751 ( n18720,n18672,n18721 );
   nand U18752 ( n18718,n18672,n18721 );
   not U18753 ( n18721,p1_addr_reg_15_ );
   nand U18754 ( n18672,n18722,n18723 );
   nand U18755 ( n18723,n18724,n18670 );
   not U18756 ( n18670,p2_addr_reg_14_ );
   or U18757 ( n18724,n18669,n18725 );
   nand U18758 ( n18722,n18669,n18725 );
   not U18759 ( n18725,p1_addr_reg_14_ );
   nand U18760 ( n18669,n18726,n18727 );
   nand U18761 ( n18727,n18728,n18667 );
   not U18762 ( n18667,p2_addr_reg_13_ );
   or U18763 ( n18728,n18666,n18729 );
   nand U18764 ( n18726,n18666,n18729 );
   not U18765 ( n18729,p1_addr_reg_13_ );
   nand U18766 ( n18666,n18730,n18731 );
   nand U18767 ( n18731,n18732,n18664 );
   not U18768 ( n18664,p2_addr_reg_12_ );
   or U18769 ( n18732,n18663,n18733 );
   nand U18770 ( n18730,n18663,n18733 );
   not U18771 ( n18733,p1_addr_reg_12_ );
   nand U18772 ( n18663,n18734,n18735 );
   nand U18773 ( n18735,n18736,n18661 );
   not U18774 ( n18661,p2_addr_reg_11_ );
   or U18775 ( n18736,n18660,n18737 );
   nand U18776 ( n18734,n18660,n18737 );
   not U18777 ( n18737,p1_addr_reg_11_ );
   nand U18778 ( n18660,n18738,n18739 );
   nand U18779 ( n18739,n18740,n13043 );
   not U18780 ( n13043,p2_addr_reg_10_ );
   or U18781 ( n18740,n18658,n18741 );
   nand U18782 ( n18738,n18658,n18741 );
   not U18783 ( n18741,p1_addr_reg_10_ );
   nand U18784 ( n18658,n18742,n18743 );
   nand U18785 ( n18743,n18744,n18704 );
   not U18786 ( n18704,p2_addr_reg_9_ );
   nand U18787 ( n18744,n18745,p1_addr_reg_9_ );
   or U18788 ( n18742,n18745,p1_addr_reg_9_ );
   not U18789 ( n18745,n18703 );
   nand U18790 ( n18703,n18746,n18747 );
   nand U18791 ( n18747,n18748,n13117 );
   not U18792 ( n13117,p2_addr_reg_8_ );
   nand U18793 ( n18748,n18749,p1_addr_reg_8_ );
   or U18794 ( n18746,n18749,p1_addr_reg_8_ );
   not U18795 ( n18749,n18701 );
   nand U18796 ( n18701,n18750,n18751 );
   nand U18797 ( n18751,n18752,n13161 );
   not U18798 ( n13161,p2_addr_reg_7_ );
   nand U18799 ( n18752,n18753,p1_addr_reg_7_ );
   or U18800 ( n18750,n18753,p1_addr_reg_7_ );
   not U18801 ( n18753,n18699 );
   nand U18802 ( n18699,n18754,n18755 );
   nand U18803 ( n18755,n18756,n13196 );
   not U18804 ( n13196,p2_addr_reg_6_ );
   nand U18805 ( n18756,n18757,p1_addr_reg_6_ );
   or U18806 ( n18754,n18757,p1_addr_reg_6_ );
   not U18807 ( n18757,n18695 );
   nand U18808 ( n18695,n18758,n18759 );
   nand U18809 ( n18759,n18760,n18693 );
   not U18810 ( n18693,p2_addr_reg_5_ );
   nand U18811 ( n18760,n18761,p1_addr_reg_5_ );
   or U18812 ( n18758,n18761,p1_addr_reg_5_ );
   not U18813 ( n18761,n18692 );
   nand U18814 ( n18692,n18762,n18763 );
   nand U18815 ( n18763,n18764,n18690 );
   not U18816 ( n18690,p2_addr_reg_4_ );
   or U18817 ( n18764,n18689,n16706 );
   nand U18818 ( n18762,n18689,n16706 );
   not U18819 ( n16706,p1_addr_reg_4_ );
   nand U18820 ( n18689,n18765,n18766 );
   nand U18821 ( n18766,n18767,n18687 );
   not U18822 ( n18687,p2_addr_reg_3_ );
   nand U18823 ( n18767,n18768,p1_addr_reg_3_ );
   or U18824 ( n18765,n18768,p1_addr_reg_3_ );
   not U18825 ( n18768,n18686 );
   nand U18826 ( n18686,n18769,n18770 );
   nand U18827 ( n18770,n18771,n18684 );
   not U18828 ( n18684,p2_addr_reg_2_ );
   nand U18829 ( n18771,n18772,p1_addr_reg_2_ );
   or U18830 ( n18769,n18772,p1_addr_reg_2_ );
   not U18831 ( n18772,n18683 );
   nand U18832 ( n18683,n18773,n18774 );
   nand U18833 ( n18774,n18775,n18776 );
   not U18834 ( n18776,p2_addr_reg_1_ );
   nand U18835 ( n18775,n18696,p1_addr_reg_1_ );
   or U18836 ( n18773,n18696,p1_addr_reg_1_ );
   and U18837 ( n18696,p1_addr_reg_0_,p2_addr_reg_0_ );
   xor U18838 ( n18705,p2_addr_reg_19_,p1_addr_reg_19_ );
endmodule
