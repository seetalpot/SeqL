
module b14 ( datai_31_, datai_30_, datai_29_, datai_28_, datai_27_, datai_26_,
datai_25_, datai_24_, datai_23_, datai_22_, datai_21_, datai_20_,
datai_19_, datai_18_, datai_17_, datai_16_, datai_15_, datai_14_,
datai_13_, datai_12_, datai_11_, datai_10_, datai_9_, datai_8_,
datai_7_, datai_6_, datai_5_, datai_4_, datai_3_, datai_2_, datai_1_,
datai_0_, ir_reg_0_, ir_reg_1_, ir_reg_2_, ir_reg_3_, ir_reg_4_,
ir_reg_5_, ir_reg_6_, ir_reg_7_, ir_reg_8_, ir_reg_9_, ir_reg_10_,
ir_reg_11_, ir_reg_12_, ir_reg_13_, ir_reg_14_, ir_reg_15_, ir_reg_16_,
ir_reg_17_, ir_reg_18_, ir_reg_19_, ir_reg_20_, ir_reg_21_, ir_reg_22_,
ir_reg_23_, ir_reg_24_, ir_reg_25_, ir_reg_26_, ir_reg_27_, ir_reg_28_,
ir_reg_29_, ir_reg_30_, ir_reg_31_, d_reg_0_, d_reg_1_, d_reg_2_,
d_reg_3_, d_reg_4_, d_reg_5_, d_reg_6_, d_reg_7_, d_reg_8_, d_reg_9_,
d_reg_10_, d_reg_11_, d_reg_12_, d_reg_13_, d_reg_14_, d_reg_15_,
d_reg_16_, d_reg_17_, d_reg_18_, d_reg_19_, d_reg_20_, d_reg_21_,
d_reg_22_, d_reg_23_, d_reg_24_, d_reg_25_, d_reg_26_, d_reg_27_,
d_reg_28_, d_reg_29_, d_reg_30_, d_reg_31_, reg0_reg_0_, reg0_reg_1_,
reg0_reg_2_, reg0_reg_3_, reg0_reg_4_, reg0_reg_5_, reg0_reg_6_,
reg0_reg_7_, reg0_reg_8_, reg0_reg_9_, reg0_reg_10_, reg0_reg_11_,
reg0_reg_12_, reg0_reg_13_, reg0_reg_14_, reg0_reg_15_, reg0_reg_16_,
reg0_reg_17_, reg0_reg_18_, reg0_reg_19_, reg0_reg_20_, reg0_reg_21_,
reg0_reg_22_, reg0_reg_23_, reg0_reg_24_, reg0_reg_25_, reg0_reg_26_,
reg0_reg_27_, reg0_reg_28_, reg0_reg_29_, reg0_reg_30_, reg0_reg_31_,
reg1_reg_0_, reg1_reg_1_, reg1_reg_2_, reg1_reg_3_, reg1_reg_4_,
reg1_reg_5_, reg1_reg_6_, reg1_reg_7_, reg1_reg_8_, reg1_reg_9_,
reg1_reg_10_, reg1_reg_11_, reg1_reg_12_, reg1_reg_13_, reg1_reg_14_,
reg1_reg_15_, reg1_reg_16_, reg1_reg_17_, reg1_reg_18_, reg1_reg_19_,
reg1_reg_20_, reg1_reg_21_, reg1_reg_22_, reg1_reg_23_, reg1_reg_24_,
reg1_reg_25_, reg1_reg_26_, reg1_reg_27_, reg1_reg_28_, reg1_reg_29_,
reg1_reg_30_, reg1_reg_31_, reg2_reg_0_, reg2_reg_1_, reg2_reg_2_,
reg2_reg_3_, reg2_reg_4_, reg2_reg_5_, reg2_reg_6_, reg2_reg_7_,
reg2_reg_8_, reg2_reg_9_, reg2_reg_10_, reg2_reg_11_, reg2_reg_12_,
reg2_reg_13_, reg2_reg_14_, reg2_reg_15_, reg2_reg_16_, reg2_reg_17_,
reg2_reg_18_, reg2_reg_19_, reg2_reg_20_, reg2_reg_21_, reg2_reg_22_,
reg2_reg_23_, reg2_reg_24_, reg2_reg_25_, reg2_reg_26_, reg2_reg_27_,
reg2_reg_28_, reg2_reg_29_, reg2_reg_30_, reg2_reg_31_, addr_reg_19_,
addr_reg_18_, addr_reg_17_, addr_reg_16_, addr_reg_15_, addr_reg_14_,
addr_reg_13_, addr_reg_12_, addr_reg_11_, addr_reg_10_, addr_reg_9_,
addr_reg_8_, addr_reg_7_, addr_reg_6_, addr_reg_5_, addr_reg_4_,
addr_reg_3_, addr_reg_2_, addr_reg_1_, addr_reg_0_, datao_reg_0_,
datao_reg_1_, datao_reg_2_, datao_reg_3_, datao_reg_4_, datao_reg_5_,
datao_reg_6_, datao_reg_7_, datao_reg_8_, datao_reg_9_, datao_reg_10_,
datao_reg_11_, datao_reg_12_, datao_reg_13_, datao_reg_14_,
datao_reg_15_, datao_reg_16_, datao_reg_17_, datao_reg_18_,
datao_reg_19_, datao_reg_20_, datao_reg_21_, datao_reg_22_,
datao_reg_23_, datao_reg_24_, datao_reg_25_, datao_reg_26_,
datao_reg_27_, datao_reg_28_, datao_reg_29_, datao_reg_30_,
datao_reg_31_, b_reg, reg3_reg_15_, reg3_reg_26_, reg3_reg_6_,
reg3_reg_18_, reg3_reg_2_, reg3_reg_11_, reg3_reg_22_, reg3_reg_13_,
reg3_reg_20_, reg3_reg_0_, reg3_reg_9_, reg3_reg_4_, reg3_reg_24_,
reg3_reg_17_, reg3_reg_5_, reg3_reg_16_, reg3_reg_25_, reg3_reg_12_,
reg3_reg_21_, reg3_reg_1_, reg3_reg_8_, reg3_reg_28_, reg3_reg_19_,
reg3_reg_3_, reg3_reg_10_, reg3_reg_23_, reg3_reg_14_, reg3_reg_27_,
reg3_reg_7_, state_reg, u3352, u3351, u3350, u3349, u3348, u3347,
u3346, u3345, u3344, u3343, u3342, u3341, u3340, u3339, u3338, u3337,
u3336, u3335, u3334, u3333, u3332, u3331, u3330, u3329, u3328, u3327,
u3326, u3325, u3324, u3323, u3322, u3321, u3458, u3459, u3320, u3319,
u3318, u3317, u3316, u3315, u3314, u3313, u3312, u3311, u3310, u3309,
u3308, u3307, u3306, u3305, u3304, u3303, u3302, u3301, u3300, u3299,
u3298, u3297, u3296, u3295, u3294, u3293, u3292, u3291, u3467, u3469,
u3471, u3473, u3475, u3477, u3479, u3481, u3483, u3485, u3487, u3489,
u3491, u3493, u3495, u3497, u3499, u3501, u3503, u3505, u3506, u3507,
u3508, u3509, u3510, u3511, u3512, u3513, u3514, u3515, u3516, u3517,
u3518, u3519, u3520, u3521, u3522, u3523, u3524, u3525, u3526, u3527,
u3528, u3529, u3530, u3531, u3532, u3533, u3534, u3535, u3536, u3537,
u3538, u3539, u3540, u3541, u3542, u3543, u3544, u3545, u3546, u3547,
u3548, u3549, u3290, u3289, u3288, u3287, u3286, u3285, u3284, u3283,
u3282, u3281, u3280, u3279, u3278, u3277, u3276, u3275, u3274, u3273,
u3272, u3271, u3270, u3269, u3268, u3267, u3266, u3265, u3264, u3263,
u3262, u3354, u3261, u3260, u3259, u3258, u3257, u3256, u3255, u3254,
u3253, u3252, u3251, u3250, u3249, u3248, u3247, u3246, u3245, u3244,
u3243, u3242, u3241, u3240, u3550, u3551, u3552, u3553, u3554, u3555,
u3556, u3557, u3558, u3559, u3560, u3561, u3562, u3563, u3564, u3565,
u3566, u3567, u3568, u3569, u3570, u3571, u3572, u3573, u3574, u3575,
u3576, u3577, u3578, u3579, u3580, u3581, u3239, u3238, u3237, u3236,
u3235, u3234, u3233, u3232, u3231, u3230, u3229, u3228, u3227, u3226,
u3225, u3224, u3223, u3222, u3221, u3220, u3219, u3218, u3217, u3216,
u3215, u3214, u3213, u3212, u3211, u3210, u3149, u3148, u4043 );
input datai_31_, datai_30_, datai_29_, datai_28_, datai_27_, datai_26_,
datai_25_, datai_24_, datai_23_, datai_22_, datai_21_, datai_20_,
datai_19_, datai_18_, datai_17_, datai_16_, datai_15_, datai_14_,
datai_13_, datai_12_, datai_11_, datai_10_, datai_9_, datai_8_,
datai_7_, datai_6_, datai_5_, datai_4_, datai_3_, datai_2_, datai_1_,
datai_0_, ir_reg_0_, ir_reg_1_, ir_reg_2_, ir_reg_3_, ir_reg_4_,
ir_reg_5_, ir_reg_6_, ir_reg_7_, ir_reg_8_, ir_reg_9_, ir_reg_10_,
ir_reg_11_, ir_reg_12_, ir_reg_13_, ir_reg_14_, ir_reg_15_,
ir_reg_16_, ir_reg_17_, ir_reg_18_, ir_reg_19_, ir_reg_20_,
ir_reg_21_, ir_reg_22_, ir_reg_23_, ir_reg_24_, ir_reg_25_,
ir_reg_26_, ir_reg_27_, ir_reg_28_, ir_reg_29_, ir_reg_30_,
ir_reg_31_, d_reg_0_, d_reg_1_, d_reg_2_, d_reg_3_, d_reg_4_,
d_reg_5_, d_reg_6_, d_reg_7_, d_reg_8_, d_reg_9_, d_reg_10_,
d_reg_11_, d_reg_12_, d_reg_13_, d_reg_14_, d_reg_15_, d_reg_16_,
d_reg_17_, d_reg_18_, d_reg_19_, d_reg_20_, d_reg_21_, d_reg_22_,
d_reg_23_, d_reg_24_, d_reg_25_, d_reg_26_, d_reg_27_, d_reg_28_,
d_reg_29_, d_reg_30_, d_reg_31_, reg0_reg_0_, reg0_reg_1_,
reg0_reg_2_, reg0_reg_3_, reg0_reg_4_, reg0_reg_5_, reg0_reg_6_,
reg0_reg_7_, reg0_reg_8_, reg0_reg_9_, reg0_reg_10_, reg0_reg_11_,
reg0_reg_12_, reg0_reg_13_, reg0_reg_14_, reg0_reg_15_, reg0_reg_16_,
reg0_reg_17_, reg0_reg_18_, reg0_reg_19_, reg0_reg_20_, reg0_reg_21_,
reg0_reg_22_, reg0_reg_23_, reg0_reg_24_, reg0_reg_25_, reg0_reg_26_,
reg0_reg_27_, reg0_reg_28_, reg0_reg_29_, reg0_reg_30_, reg0_reg_31_,
reg1_reg_0_, reg1_reg_1_, reg1_reg_2_, reg1_reg_3_, reg1_reg_4_,
reg1_reg_5_, reg1_reg_6_, reg1_reg_7_, reg1_reg_8_, reg1_reg_9_,
reg1_reg_10_, reg1_reg_11_, reg1_reg_12_, reg1_reg_13_, reg1_reg_14_,
reg1_reg_15_, reg1_reg_16_, reg1_reg_17_, reg1_reg_18_, reg1_reg_19_,
reg1_reg_20_, reg1_reg_21_, reg1_reg_22_, reg1_reg_23_, reg1_reg_24_,
reg1_reg_25_, reg1_reg_26_, reg1_reg_27_, reg1_reg_28_, reg1_reg_29_,
reg1_reg_30_, reg1_reg_31_, reg2_reg_0_, reg2_reg_1_, reg2_reg_2_,
reg2_reg_3_, reg2_reg_4_, reg2_reg_5_, reg2_reg_6_, reg2_reg_7_,
reg2_reg_8_, reg2_reg_9_, reg2_reg_10_, reg2_reg_11_, reg2_reg_12_,
reg2_reg_13_, reg2_reg_14_, reg2_reg_15_, reg2_reg_16_, reg2_reg_17_,
reg2_reg_18_, reg2_reg_19_, reg2_reg_20_, reg2_reg_21_, reg2_reg_22_,
reg2_reg_23_, reg2_reg_24_, reg2_reg_25_, reg2_reg_26_, reg2_reg_27_,
reg2_reg_28_, reg2_reg_29_, reg2_reg_30_, reg2_reg_31_, addr_reg_19_,
addr_reg_18_, addr_reg_17_, addr_reg_16_, addr_reg_15_, addr_reg_14_,
addr_reg_13_, addr_reg_12_, addr_reg_11_, addr_reg_10_, addr_reg_9_,
addr_reg_8_, addr_reg_7_, addr_reg_6_, addr_reg_5_, addr_reg_4_,
addr_reg_3_, addr_reg_2_, addr_reg_1_, addr_reg_0_, datao_reg_0_,
datao_reg_1_, datao_reg_2_, datao_reg_3_, datao_reg_4_, datao_reg_5_,
datao_reg_6_, datao_reg_7_, datao_reg_8_, datao_reg_9_, datao_reg_10_,
datao_reg_11_, datao_reg_12_, datao_reg_13_, datao_reg_14_,
datao_reg_15_, datao_reg_16_, datao_reg_17_, datao_reg_18_,
datao_reg_19_, datao_reg_20_, datao_reg_21_, datao_reg_22_,
datao_reg_23_, datao_reg_24_, datao_reg_25_, datao_reg_26_,
datao_reg_27_, datao_reg_28_, datao_reg_29_, datao_reg_30_,
datao_reg_31_, b_reg, reg3_reg_15_, reg3_reg_26_, reg3_reg_6_,
reg3_reg_18_, reg3_reg_2_, reg3_reg_11_, reg3_reg_22_, reg3_reg_13_,
reg3_reg_20_, reg3_reg_0_, reg3_reg_9_, reg3_reg_4_, reg3_reg_24_,
reg3_reg_17_, reg3_reg_5_, reg3_reg_16_, reg3_reg_25_, reg3_reg_12_,
reg3_reg_21_, reg3_reg_1_, reg3_reg_8_, reg3_reg_28_, reg3_reg_19_,
reg3_reg_3_, reg3_reg_10_, reg3_reg_23_, reg3_reg_14_, reg3_reg_27_,
reg3_reg_7_, state_reg;
output u3352, u3351, u3350, u3349, u3348, u3347, u3346, u3345, u3344, u3343,
u3342, u3341, u3340, u3339, u3338, u3337, u3336, u3335, u3334, u3333,
u3332, u3331, u3330, u3329, u3328, u3327, u3326, u3325, u3324, u3323,
u3322, u3321, u3458, u3459, u3320, u3319, u3318, u3317, u3316, u3315,
u3314, u3313, u3312, u3311, u3310, u3309, u3308, u3307, u3306, u3305,
u3304, u3303, u3302, u3301, u3300, u3299, u3298, u3297, u3296, u3295,
u3294, u3293, u3292, u3291, u3467, u3469, u3471, u3473, u3475, u3477,
u3479, u3481, u3483, u3485, u3487, u3489, u3491, u3493, u3495, u3497,
u3499, u3501, u3503, u3505, u3506, u3507, u3508, u3509, u3510, u3511,
u3512, u3513, u3514, u3515, u3516, u3517, u3518, u3519, u3520, u3521,
u3522, u3523, u3524, u3525, u3526, u3527, u3528, u3529, u3530, u3531,
u3532, u3533, u3534, u3535, u3536, u3537, u3538, u3539, u3540, u3541,
u3542, u3543, u3544, u3545, u3546, u3547, u3548, u3549, u3290, u3289,
u3288, u3287, u3286, u3285, u3284, u3283, u3282, u3281, u3280, u3279,
u3278, u3277, u3276, u3275, u3274, u3273, u3272, u3271, u3270, u3269,
u3268, u3267, u3266, u3265, u3264, u3263, u3262, u3354, u3261, u3260,
u3259, u3258, u3257, u3256, u3255, u3254, u3253, u3252, u3251, u3250,
u3249, u3248, u3247, u3246, u3245, u3244, u3243, u3242, u3241, u3240,
u3550, u3551, u3552, u3553, u3554, u3555, u3556, u3557, u3558, u3559,
u3560, u3561, u3562, u3563, u3564, u3565, u3566, u3567, u3568, u3569,
u3570, u3571, u3572, u3573, u3574, u3575, u3576, u3577, u3578, u3579,
u3580, u3581, u3239, u3238, u3237, u3236, u3235, u3234, u3233, u3232,
u3231, u3230, u3229, u3228, u3227, u3226, u3225, u3224, u3223, u3222,
u3221, u3220, u3219, u3218, u3217, u3216, u3215, u3214, u3213, u3212,
u3211, u3210, u3149, u3148, u4043;
wire   n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
n10805, n10806, n10807, n5442, n5444, n5446, n5448, n5449, n5450,
n5451, n5452, n5454, n5456, n5458, n5460, n5462, n5464, n5466, n5468,
n5470, n5472, n5474, n5476, n5478, n5480, n5482, n5484, n5486, n5488,
n5490, n5492, n5494, n5496, n5498, n5500, n5502, n5504, n5506, n5508,
n5510, n5512, n5514, n5516, n5518, n5520, n5522, n5524, n5526, n5528,
n5530, n5532, n5534, n5536, n5538, n5540, n5542, n5544, n5546, n5548,
n5550, n5552, n5554, n5556, n5558, n5560, n5562, n5564, n5566, n5568,
n5570, n5572, n5574, n5576, n5578, n5580, n5582, n5584, n5586, n5588,
n5590, n5592, n5594, n5596, n5598, n5600, n5602, n5604, n5606, n5608,
n5610, n5612, n5614, n5616, n5618, n5620, n5622, n5624, n5626, n5628,
n5630, n5632, n5634, n5636, n5638, n5640, n5642, n5644, n5646, n5648,
n5650, n5652, n5654, n5656, n5658, n5660, n5662, n5664, n5666, n5668,
n5670, n5672, n5674, n5676, n5678, n5680, n5682, n5684, n5686, n5688,
n5690, n5692, n5694, n5696, n5698, n5700, n5702, n5704, n5706, n5708,
n5710, n5712, n5714, n5716, n5718, n5720, n5722, n5724, n5726, n5728,
n5730, n5732, n5734, n5736, n5738, n5740, n5742, n5744, n5746, n5748,
n5750, n5752, n5754, n5756, n5758, n5760, n5762, n5764, n5766, n5768,
n5770, n5772, n5774, n5776, n5778, n5780, n5782, n5784, n5786, n5788,
n5790, n5792, n5794, n5796, n5798, n5800, n5802, n5804, n5806, n5808,
n5810, n5812, n5814, n5816, n5818, n5820, n5822, n5824, n5826, n5828,
n5830, n5832, n5834, n5836, n5838, n5840, n5842, n5844, n5846, n5848,
n5850, n5852, n5854, n5856, n5858, n5860, n5862, n5864, n5866, n5868,
n5870, n5872, n5874, n5876, n5878, n5880, n5882, n5884, n5886, n5888,
n5890, n5892, n5894, n5896, n5898, n5900, n5902, n5904, n5906, n5908,
n5910, n5912, n5914, n5916, n5918, n5920, n5922, n5924, n5926, n5928,
n5930, n5932, n5933, n5934, n5935, n5936, n5937, n5939, n5940, n5941,
n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
n5972, n5973, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
n10794, n10795, n10796;

   not U5687 ( n5442,n6016 );
   not U5688 ( u4043,n6016 );
   nor U5689 ( n5444,n8692,n8693 );
   not U5690 ( u3243,n5444 );
   nor U5691 ( n5446,n8635,n8636 );
   not U5692 ( u3245,n5446 );
   not U5693 ( n5448,n5451 );
   buf U5694 ( n5449,n8268 );
   not U5695 ( n5450,n8282 );
   buf U5696 ( n5451,n6744 );
   nor U5697 ( n5452,n8608,n8609 );
   not U5698 ( u3246,n5452 );
   nor U5699 ( n5454,n8578,n8579 );
   not U5700 ( u3247,n5454 );
   nor U5701 ( n5456,n8551,n8552 );
   not U5702 ( u3248,n5456 );
   nor U5703 ( n5458,n8523,n8524 );
   not U5704 ( u3249,n5458 );
   nor U5705 ( n5460,n8495,n8496 );
   not U5706 ( u3250,n5460 );
   nor U5707 ( n5462,n8468,n8469 );
   not U5708 ( u3251,n5462 );
   nor U5709 ( n5464,n8438,n8439 );
   not U5710 ( u3252,n5464 );
   nor U5711 ( n5466,n8411,n8412 );
   not U5712 ( u3253,n5466 );
   nor U5713 ( n5468,n8383,n8384 );
   not U5714 ( u3254,n5468 );
   nor U5715 ( n5470,n8355,n8356 );
   not U5716 ( u3255,n5470 );
   nor U5717 ( n5472,n8328,n8329 );
   not U5718 ( u3256,n5472 );
   nor U5719 ( n5474,n8299,n8300 );
   not U5720 ( u3257,n5474 );
   nor U5721 ( n5476,n8269,n8270 );
   not U5722 ( u3258,n5476 );
   and U5723 ( n5478,n8238,n8239 );
   not U5724 ( u3259,n5478 );
   and U5725 ( n5480,n8208,n8209 );
   not U5726 ( u3260,n5480 );
   and U5727 ( n5482,n8198,n8199 );
   not U5728 ( u3261,n5482 );
   and U5729 ( n5484,n6677,n6678 );
   not U5730 ( u3354,n5484 );
   and U5731 ( n5486,n8004,n8005 );
   not U5732 ( u3262,n5486 );
   and U5733 ( n5488,n7959,n7960 );
   not U5734 ( u3263,n5488 );
   and U5735 ( n5490,n7897,n7898 );
   not U5736 ( u3264,n5490 );
   and U5737 ( n5492,n7866,n7867 );
   not U5738 ( u3265,n5492 );
   and U5739 ( n5494,n7836,n7837 );
   not U5740 ( u3266,n5494 );
   and U5741 ( n5496,n7776,n7777 );
   not U5742 ( u3267,n5496 );
   and U5743 ( n5498,n7732,n7733 );
   not U5744 ( u3268,n5498 );
   and U5745 ( n5500,n7694,n7695 );
   not U5746 ( u3269,n5500 );
   and U5747 ( n5502,n7654,n7655 );
   not U5748 ( u3270,n5502 );
   and U5749 ( n5504,n7632,n7633 );
   not U5750 ( u3271,n5504 );
   and U5751 ( n5506,n7606,n7607 );
   not U5752 ( u3272,n5506 );
   and U5753 ( n5508,n7570,n7571 );
   not U5754 ( u3273,n5508 );
   and U5755 ( n5510,n7534,n7535 );
   not U5756 ( u3274,n5510 );
   and U5757 ( n5512,n7497,n7498 );
   not U5758 ( u3275,n5512 );
   and U5759 ( n5514,n7465,n7466 );
   not U5760 ( u3276,n5514 );
   and U5761 ( n5516,n7430,n7431 );
   not U5762 ( u3277,n5516 );
   and U5763 ( n5518,n7403,n7404 );
   not U5764 ( u3278,n5518 );
   and U5765 ( n5520,n7369,n7370 );
   not U5766 ( u3279,n5520 );
   and U5767 ( n5522,n7319,n7320 );
   not U5768 ( u3280,n5522 );
   and U5769 ( n5524,n7291,n7292 );
   not U5770 ( u3281,n5524 );
   and U5771 ( n5526,n7248,n7249 );
   not U5772 ( u3282,n5526 );
   and U5773 ( n5528,n7204,n7205 );
   not U5774 ( u3283,n5528 );
   and U5775 ( n5530,n7167,n7168 );
   not U5776 ( u3284,n5530 );
   and U5777 ( n5532,n7129,n7130 );
   not U5778 ( u3285,n5532 );
   and U5779 ( n5534,n7098,n7099 );
   not U5780 ( u3286,n5534 );
   and U5781 ( n5536,n7068,n7069 );
   not U5782 ( u3287,n5536 );
   and U5783 ( n5538,n7024,n7025 );
   not U5784 ( u3288,n5538 );
   and U5785 ( n5540,n6997,n6998 );
   not U5786 ( u3289,n5540 );
   and U5787 ( n5542,n6981,n6982 );
   not U5788 ( u3290,n5542 );
   and U5789 ( n5544,n6111,n6112 );
   not U5790 ( u3549,n5544 );
   and U5791 ( n5546,n6116,n6117 );
   not U5792 ( u3548,n5546 );
   and U5793 ( n5548,n6119,n6120 );
   not U5794 ( u3547,n5548 );
   and U5795 ( n5550,n6122,n6123 );
   not U5796 ( u3546,n5550 );
   and U5797 ( n5552,n6125,n6126 );
   not U5798 ( u3545,n5552 );
   and U5799 ( n5554,n6128,n6129 );
   not U5800 ( u3544,n5554 );
   and U5801 ( n5556,n6131,n6132 );
   not U5802 ( u3543,n5556 );
   and U5803 ( n5558,n6134,n6135 );
   not U5804 ( u3542,n5558 );
   and U5805 ( n5560,n6137,n6138 );
   not U5806 ( u3541,n5560 );
   and U5807 ( n5562,n6140,n6141 );
   not U5808 ( u3540,n5562 );
   and U5809 ( n5564,n6143,n6144 );
   not U5810 ( u3539,n5564 );
   and U5811 ( n5566,n6146,n6147 );
   not U5812 ( u3538,n5566 );
   and U5813 ( n5568,n6149,n6150 );
   not U5814 ( u3537,n5568 );
   and U5815 ( n5570,n6152,n6153 );
   not U5816 ( u3536,n5570 );
   and U5817 ( n5572,n6155,n6156 );
   not U5818 ( u3535,n5572 );
   and U5819 ( n5574,n6158,n6159 );
   not U5820 ( u3534,n5574 );
   and U5821 ( n5576,n6161,n6162 );
   not U5822 ( u3533,n5576 );
   and U5823 ( n5578,n6164,n6165 );
   not U5824 ( u3532,n5578 );
   and U5825 ( n5580,n6167,n6168 );
   not U5826 ( u3531,n5580 );
   and U5827 ( n5582,n6170,n6171 );
   not U5828 ( u3530,n5582 );
   and U5829 ( n5584,n6173,n6174 );
   not U5830 ( u3529,n5584 );
   and U5831 ( n5586,n6176,n6177 );
   not U5832 ( u3528,n5586 );
   and U5833 ( n5588,n6179,n6180 );
   not U5834 ( u3527,n5588 );
   and U5835 ( n5590,n6182,n6183 );
   not U5836 ( u3526,n5590 );
   and U5837 ( n5592,n6185,n6186 );
   not U5838 ( u3525,n5592 );
   and U5839 ( n5594,n6188,n6189 );
   not U5840 ( u3524,n5594 );
   and U5841 ( n5596,n6191,n6192 );
   not U5842 ( u3523,n5596 );
   and U5843 ( n5598,n6194,n6195 );
   not U5844 ( u3522,n5598 );
   and U5845 ( n5600,n6197,n6198 );
   not U5846 ( u3521,n5600 );
   and U5847 ( n5602,n6200,n6201 );
   not U5848 ( u3520,n5602 );
   and U5849 ( n5604,n6203,n6204 );
   not U5850 ( u3519,n5604 );
   and U5851 ( n5606,n6206,n6207 );
   not U5852 ( u3518,n5606 );
   and U5853 ( n5608,n6213,n6214 );
   not U5854 ( u3517,n5608 );
   and U5855 ( n5610,n6225,n6226 );
   not U5856 ( u3516,n5610 );
   and U5857 ( n5612,n6232,n6233 );
   not U5858 ( u3515,n5612 );
   and U5859 ( n5614,n6245,n6246 );
   not U5860 ( u3514,n5614 );
   and U5861 ( n5616,n6262,n6263 );
   not U5862 ( u3513,n5616 );
   and U5863 ( n5618,n6276,n6277 );
   not U5864 ( u3512,n5618 );
   and U5865 ( n5620,n6290,n6291 );
   not U5866 ( u3511,n5620 );
   and U5867 ( n5622,n6304,n6305 );
   not U5868 ( u3510,n5622 );
   and U5869 ( n5624,n6318,n6319 );
   not U5870 ( u3509,n5624 );
   and U5871 ( n5626,n6332,n6333 );
   not U5872 ( u3508,n5626 );
   and U5873 ( n5628,n6346,n6347 );
   not U5874 ( u3507,n5628 );
   and U5875 ( n5630,n6360,n6361 );
   not U5876 ( u3506,n5630 );
   and U5877 ( n5632,n6374,n6375 );
   not U5878 ( u3505,n5632 );
   and U5879 ( n5634,n6388,n6389 );
   not U5880 ( u3503,n5634 );
   and U5881 ( n5636,n6402,n6403 );
   not U5882 ( u3501,n5636 );
   and U5883 ( n5638,n6416,n6417 );
   not U5884 ( u3499,n5638 );
   and U5885 ( n5640,n6430,n6431 );
   not U5886 ( u3497,n5640 );
   and U5887 ( n5642,n6444,n6445 );
   not U5888 ( u3495,n5642 );
   and U5889 ( n5644,n6458,n6459 );
   not U5890 ( u3493,n5644 );
   and U5891 ( n5646,n6472,n6473 );
   not U5892 ( u3491,n5646 );
   and U5893 ( n5648,n6486,n6487 );
   not U5894 ( u3489,n5648 );
   and U5895 ( n5650,n6500,n6501 );
   not U5896 ( u3487,n5650 );
   and U5897 ( n5652,n6514,n6515 );
   not U5898 ( u3485,n5652 );
   and U5899 ( n5654,n6528,n6529 );
   not U5900 ( u3483,n5654 );
   and U5901 ( n5656,n6542,n6543 );
   not U5902 ( u3481,n5656 );
   and U5903 ( n5658,n6556,n6557 );
   not U5904 ( u3479,n5658 );
   and U5905 ( n5660,n6570,n6571 );
   not U5906 ( u3477,n5660 );
   and U5907 ( n5662,n6584,n6585 );
   not U5908 ( u3475,n5662 );
   and U5909 ( n5664,n6598,n6599 );
   not U5910 ( u3473,n5664 );
   and U5911 ( n5666,n6612,n6613 );
   not U5912 ( u3471,n5666 );
   and U5913 ( n5668,n6626,n6627 );
   not U5914 ( u3469,n5668 );
   and U5915 ( n5670,n6640,n6641 );
   not U5916 ( u3467,n5670 );
   not U5917 ( n5672,n10806 );
   not U5918 ( u3291,n5672 );
   not U5919 ( n5674,n10805 );
   not U5920 ( u3292,n5674 );
   not U5921 ( n5676,n10804 );
   not U5922 ( u3293,n5676 );
   not U5923 ( n5678,n10803 );
   not U5924 ( u3294,n5678 );
   nand U5925 ( n5680,n6671,d_reg_27_ );
   not U5926 ( u3295,n5680 );
   nand U5927 ( n5682,n6671,d_reg_26_ );
   not U5928 ( u3296,n5682 );
   nand U5929 ( n5684,n6671,d_reg_25_ );
   not U5930 ( u3297,n5684 );
   not U5931 ( n5686,n10802 );
   not U5932 ( u3298,n5686 );
   not U5933 ( n5688,n10801 );
   not U5934 ( u3299,n5688 );
   nand U5935 ( n5690,n6671,d_reg_22_ );
   not U5936 ( u3300,n5690 );
   nand U5937 ( n5692,n6671,d_reg_21_ );
   not U5938 ( u3301,n5692 );
   nand U5939 ( n5694,n6671,d_reg_20_ );
   not U5940 ( u3302,n5694 );
   not U5941 ( n5696,n10800 );
   not U5942 ( u3303,n5696 );
   not U5943 ( n5698,n10799 );
   not U5944 ( u3304,n5698 );
   nand U5945 ( n5700,n6671,d_reg_17_ );
   not U5946 ( u3305,n5700 );
   nand U5947 ( n5702,n6671,d_reg_16_ );
   not U5948 ( u3306,n5702 );
   not U5949 ( n5704,n10798 );
   not U5950 ( u3307,n5704 );
   or U5951 ( n5706,n5935,n6969 );
   not U5952 ( u3308,n5706 );
   nand U5953 ( n5708,n6671,d_reg_13_ );
   not U5954 ( u3309,n5708 );
   not U5955 ( n5710,n10797 );
   not U5956 ( u3310,n5710 );
   or U5957 ( n5712,n6672,n6967 );
   not U5958 ( u3311,n5712 );
   or U5959 ( n5714,n6672,n6966 );
   not U5960 ( u3312,n5714 );
   nand U5961 ( n5716,n6671,d_reg_9_ );
   not U5962 ( u3313,n5716 );
   nand U5963 ( n5718,n6671,d_reg_8_ );
   not U5964 ( u3314,n5718 );
   or U5965 ( n5720,n6672,n6965 );
   not U5966 ( u3315,n5720 );
   or U5967 ( n5722,n5935,n6964 );
   not U5968 ( u3316,n5722 );
   or U5969 ( n5724,n6672,n6963 );
   not U5970 ( u3317,n5724 );
   or U5971 ( n5726,n5935,n6962 );
   not U5972 ( u3318,n5726 );
   nand U5973 ( n5728,n6671,d_reg_3_ );
   not U5974 ( u3319,n5728 );
   nand U5975 ( n5730,n6671,d_reg_2_ );
   not U5976 ( u3320,n5730 );
   and U5977 ( n5732,n6669,n6670 );
   not U5978 ( u3459,n5732 );
   and U5979 ( n5734,n6674,n6675 );
   not U5980 ( u3458,n5734 );
   and U5981 ( n5736,n6959,n6960 );
   not U5982 ( u3321,n5736 );
   and U5983 ( n5738,n6953,n6954 );
   not U5984 ( u3322,n5738 );
   and U5985 ( n5740,n6944,n6945 );
   not U5986 ( u3323,n5740 );
   and U5987 ( n5742,n6938,n6939 );
   not U5988 ( u3324,n5742 );
   and U5989 ( n5744,n6929,n6930 );
   not U5990 ( u3325,n5744 );
   and U5991 ( n5746,n6922,n6923 );
   not U5992 ( u3326,n5746 );
   and U5993 ( n5748,n6916,n6917 );
   not U5994 ( u3327,n5748 );
   and U5995 ( n5750,n6907,n6908 );
   not U5996 ( u3328,n5750 );
   and U5997 ( n5752,n6901,n6902 );
   not U5998 ( u3329,n5752 );
   and U5999 ( n5754,n6892,n6893 );
   not U6000 ( u3330,n5754 );
   and U6001 ( n5756,n6886,n6887 );
   not U6002 ( u3331,n5756 );
   and U6003 ( n5758,n6877,n6878 );
   not U6004 ( u3332,n5758 );
   and U6005 ( n5760,n6871,n6872 );
   not U6006 ( u3333,n5760 );
   and U6007 ( n5762,n6862,n6863 );
   not U6008 ( u3334,n5762 );
   and U6009 ( n5764,n6856,n6857 );
   not U6010 ( u3335,n5764 );
   and U6011 ( n5766,n6847,n6848 );
   not U6012 ( u3336,n5766 );
   and U6013 ( n5768,n6841,n6842 );
   not U6014 ( u3337,n5768 );
   and U6015 ( n5770,n6832,n6833 );
   not U6016 ( u3338,n5770 );
   and U6017 ( n5772,n6826,n6827 );
   not U6018 ( u3339,n5772 );
   and U6019 ( n5774,n6817,n6818 );
   not U6020 ( u3340,n5774 );
   and U6021 ( n5776,n6811,n6812 );
   not U6022 ( u3341,n5776 );
   and U6023 ( n5778,n6802,n6803 );
   not U6024 ( u3342,n5778 );
   and U6025 ( n5780,n6796,n6797 );
   not U6026 ( u3343,n5780 );
   and U6027 ( n5782,n6787,n6788 );
   not U6028 ( u3344,n5782 );
   and U6029 ( n5784,n6781,n6782 );
   not U6030 ( u3345,n5784 );
   and U6031 ( n5786,n6772,n6773 );
   not U6032 ( u3346,n5786 );
   and U6033 ( n5788,n6766,n6767 );
   not U6034 ( u3347,n5788 );
   and U6035 ( n5790,n6758,n6759 );
   not U6036 ( u3348,n5790 );
   and U6037 ( n5792,n6751,n6752 );
   not U6038 ( u3349,n5792 );
   and U6039 ( n5794,n6745,n6746 );
   not U6040 ( u3350,n5794 );
   and U6041 ( n5796,n6735,n6736 );
   not U6042 ( u3351,n5796 );
   and U6043 ( n5798,n6731,n6732 );
   not U6044 ( u3352,n5798 );
   and U6045 ( n5800,n8663,n8664 );
   not U6046 ( u3244,n5800 );
   and U6047 ( n5802,n8725,n8726 );
   not U6048 ( u3242,n5802 );
   and U6049 ( n5804,n8768,n8769 );
   not U6050 ( u3241,n5804 );
   and U6051 ( n5806,n8796,n8797 );
   not U6052 ( u3240,n5806 );
   and U6053 ( n5808,n6108,n6109 );
   not U6054 ( u3550,n5808 );
   and U6055 ( n5810,n6105,n6106 );
   not U6056 ( u3551,n5810 );
   and U6057 ( n5812,n6102,n6103 );
   not U6058 ( u3552,n5812 );
   and U6059 ( n5814,n6099,n6100 );
   not U6060 ( u3553,n5814 );
   and U6061 ( n5816,n6096,n6097 );
   not U6062 ( u3554,n5816 );
   and U6063 ( n5818,n6093,n6094 );
   not U6064 ( u3555,n5818 );
   and U6065 ( n5820,n6090,n6091 );
   not U6066 ( u3556,n5820 );
   and U6067 ( n5822,n6087,n6088 );
   not U6068 ( u3557,n5822 );
   and U6069 ( n5824,n6084,n6085 );
   not U6070 ( u3558,n5824 );
   and U6071 ( n5826,n6081,n6082 );
   not U6072 ( u3559,n5826 );
   and U6073 ( n5828,n6078,n6079 );
   not U6074 ( u3560,n5828 );
   and U6075 ( n5830,n6075,n6076 );
   not U6076 ( u3561,n5830 );
   and U6077 ( n5832,n6072,n6073 );
   not U6078 ( u3562,n5832 );
   and U6079 ( n5834,n6069,n6070 );
   not U6080 ( u3563,n5834 );
   and U6081 ( n5836,n6066,n6067 );
   not U6082 ( u3564,n5836 );
   and U6083 ( n5838,n6063,n6064 );
   not U6084 ( u3565,n5838 );
   and U6085 ( n5840,n6060,n6061 );
   not U6086 ( u3566,n5840 );
   and U6087 ( n5842,n6057,n6058 );
   not U6088 ( u3567,n5842 );
   and U6089 ( n5844,n6054,n6055 );
   not U6090 ( u3568,n5844 );
   and U6091 ( n5846,n6051,n6052 );
   not U6092 ( u3569,n5846 );
   and U6093 ( n5848,n6048,n6049 );
   not U6094 ( u3570,n5848 );
   and U6095 ( n5850,n6045,n6046 );
   not U6096 ( u3571,n5850 );
   and U6097 ( n5852,n6042,n6043 );
   not U6098 ( u3572,n5852 );
   and U6099 ( n5854,n6039,n6040 );
   not U6100 ( u3573,n5854 );
   and U6101 ( n5856,n6036,n6037 );
   not U6102 ( u3574,n5856 );
   and U6103 ( n5858,n6033,n6034 );
   not U6104 ( u3575,n5858 );
   and U6105 ( n5860,n6030,n6031 );
   not U6106 ( u3576,n5860 );
   and U6107 ( n5862,n6027,n6028 );
   not U6108 ( u3577,n5862 );
   and U6109 ( n5864,n6024,n6025 );
   not U6110 ( u3578,n5864 );
   and U6111 ( n5866,n6021,n6022 );
   not U6112 ( u3579,n5866 );
   and U6113 ( n5868,n6018,n6019 );
   not U6114 ( u3580,n5868 );
   and U6115 ( n5870,n6014,n6015 );
   not U6116 ( u3581,n5870 );
   and U6117 ( n5872,n8827,n8828 );
   not U6118 ( u3239,n5872 );
   and U6119 ( n5874,n9442,n9443 );
   not U6120 ( u3238,n5874 );
   and U6121 ( n5876,n9463,n9464 );
   not U6122 ( u3237,n5876 );
   and U6123 ( n5878,n9497,n9498 );
   not U6124 ( u3236,n5878 );
   and U6125 ( n5880,n9518,n9519 );
   not U6126 ( u3235,n5880 );
   and U6127 ( n5882,n9535,n9536 );
   not U6128 ( u3234,n5882 );
   and U6129 ( n5884,n9558,n9559 );
   not U6130 ( u3233,n5884 );
   and U6131 ( n5886,n9580,n9581 );
   not U6132 ( u3232,n5886 );
   and U6133 ( n5888,n9597,n9598 );
   not U6134 ( u3231,n5888 );
   and U6135 ( n5890,n9624,n9625 );
   not U6136 ( u3230,n5890 );
   and U6137 ( n5892,n9649,n9650 );
   not U6138 ( u3229,n5892 );
   and U6139 ( n5894,n9658,n9659 );
   not U6140 ( u3228,n5894 );
   and U6141 ( n5896,n9673,n9674 );
   not U6142 ( u3227,n5896 );
   and U6143 ( n5898,n9689,n9690 );
   not U6144 ( u3226,n5898 );
   and U6145 ( n5900,n9706,n9707 );
   not U6146 ( u3225,n5900 );
   and U6147 ( n5902,n9730,n9731 );
   not U6148 ( u3224,n5902 );
   and U6149 ( n5904,n9746,n9747 );
   not U6150 ( u3223,n5904 );
   and U6151 ( n5906,n9770,n9771 );
   not U6152 ( u3222,n5906 );
   and U6153 ( n5908,n9790,n9791 );
   not U6154 ( u3221,n5908 );
   and U6155 ( n5910,n9816,n9817 );
   not U6156 ( u3220,n5910 );
   and U6157 ( n5912,n9843,n9844 );
   not U6158 ( u3219,n5912 );
   and U6159 ( n5914,n9856,n9857 );
   not U6160 ( u3218,n5914 );
   and U6161 ( n5916,n9873,n9874 );
   not U6162 ( u3217,n5916 );
   and U6163 ( n5918,n9908,n9909 );
   not U6164 ( u3216,n5918 );
   and U6165 ( n5920,n9931,n9932 );
   not U6166 ( u3215,n5920 );
   and U6167 ( n5922,n9952,n9953 );
   not U6168 ( u3214,n5922 );
   and U6169 ( n5924,n9967,n9968 );
   not U6170 ( u3213,n5924 );
   and U6171 ( n5926,n9983,n9984 );
   not U6172 ( u3212,n5926 );
   and U6173 ( n5928,n9999,n10000 );
   not U6174 ( u3211,n5928 );
   and U6175 ( n5930,n10461,n10462 );
   not U6176 ( u3210,n5930 );
   not U6177 ( n5932,n5972 );
   buf U6178 ( n5933,n6115 );
   buf U6179 ( n5934,n6224 );
   buf U6180 ( n5935,n6672 );
   not U6181 ( n5936,n5442 );
   nand U6182 ( n5937,n10764,n5936 );
   not U6183 ( u3148,n5937 );
   not U6184 ( n5939,n5937 );
   buf U6185 ( n5940,n10021 );
   buf U6186 ( n5941,n6113 );
   buf U6187 ( n5942,n6215 );
   nand U6188 ( n5944,n6666,n8040 );
   nand U6189 ( n5943,n6666,n8040 );
   buf U6190 ( n5945,n6740 );
   not U6191 ( n5946,n5945 );
   not U6192 ( n5948,n5945 );
   not U6193 ( n5947,n5945 );
   not U6194 ( n5949,n8819 );
   not U6195 ( n5950,n5949 );
   not U6196 ( n5951,n5949 );
   and U6197 ( n5952,n10666,n10665 );
   not U6198 ( n5953,n5952 );
   not U6199 ( n5956,n5952 );
   not U6200 ( n5954,n5952 );
   not U6201 ( n5955,n5952 );
   and U6202 ( n5957,n10664,n10665 );
   not U6203 ( n5958,n5957 );
   not U6204 ( n5961,n5957 );
   not U6205 ( n5959,n5957 );
   not U6206 ( n5960,n5957 );
   or U6207 ( n5962,n8734,n8732 );
   not U6208 ( n5963,n5962 );
   not U6209 ( n5966,n5962 );
   not U6210 ( n5964,n5962 );
   not U6211 ( n5965,n5962 );
   or U6212 ( n5967,n9270,n5951 );
   not U6213 ( n5968,n5967 );
   not U6214 ( n5971,n5967 );
   not U6215 ( n5969,n5967 );
   not U6216 ( n5970,n5967 );
   buf U6217 ( n5972,state_reg );
   not U6218 ( n5973,n5972 );
   not U6219 ( n5975,n5972 );
   not U6220 ( u3149,n5972 );
   not U6221 ( n5976,n6683 );
   not U6222 ( n5977,n6692 );
   not U6223 ( n5978,n6685 );
   not U6224 ( n5979,n10125 );
   buf U6225 ( n5980,n8282 );
   not U6226 ( n5981,n6730 );
   nand U6227 ( n5982,n10636,n10637 );
   not U6228 ( n5983,n9489 );
   not U6229 ( n5984,n9449 );
   not U6230 ( n5985,n9494 );
   buf U6231 ( n5986,n6718 );
   not U6232 ( n5987,ir_reg_31_ );
   not U6233 ( n5988,n8265 );
   buf U6234 ( n5989,n6700 );
   not U6235 ( n5991,n10033 );
   not U6236 ( n5990,n10033 );
   not U6237 ( n5992,n6729 );
   not U6238 ( n5993,n9557 );
   not U6239 ( n5994,n6240 );
   buf U6240 ( n5995,n10125 );
   not U6241 ( n5996,n9889 );
   not U6242 ( n5997,n6223 );
   nor U6243 ( n5999,n7834,n7522 );
   nor U6244 ( n5998,n7834,n7522 );
   not U6245 ( n6000,n6989 );
   nor U6246 ( n6001,n8734,n8806 );
   nand U6247 ( n6002,n6210,n8232 );
   nor U6248 ( n6003,n10665,n10664 );
   not U6249 ( n6004,n6003 );
   not U6250 ( n6006,n6003 );
   not U6251 ( n6005,n6003 );
   buf U6252 ( n6007,n10015 );
   not U6253 ( n6008,n6007 );
   not U6254 ( n6011,n6007 );
   not U6255 ( n6009,n6007 );
   not U6256 ( n6010,n6007 );
   not U6257 ( n6013,n6218 );
   not U6258 ( n6012,n6218 );
   nand U6259 ( n6015,datao_reg_31_,n5936 );
   nand U6260 ( n6014,n5442,n6017 );
   nand U6261 ( n6019,datao_reg_30_,n5936 );
   nand U6262 ( n6018,n5442,n6020 );
   nand U6263 ( n6022,datao_reg_29_,n6016 );
   nand U6264 ( n6021,n5442,n6023 );
   nand U6265 ( n6025,datao_reg_28_,n5936 );
   nand U6266 ( n6024,n10807,n6026 );
   nand U6267 ( n6028,datao_reg_27_,n5936 );
   nand U6268 ( n6027,n10807,n6029 );
   nand U6269 ( n6031,datao_reg_26_,n5936 );
   nand U6270 ( n6030,n5442,n6032 );
   nand U6271 ( n6034,datao_reg_25_,n5936 );
   nand U6272 ( n6033,n5442,n6035 );
   nand U6273 ( n6037,datao_reg_24_,n5936 );
   nand U6274 ( n6036,n10807,n6038 );
   nand U6275 ( n6040,datao_reg_23_,n5936 );
   nand U6276 ( n6039,n10807,n6041 );
   nand U6277 ( n6043,datao_reg_22_,n5936 );
   nand U6278 ( n6042,n5442,n6044 );
   nand U6279 ( n6046,datao_reg_21_,n5936 );
   nand U6280 ( n6045,n5442,n6047 );
   nand U6281 ( n6049,datao_reg_20_,n5936 );
   nand U6282 ( n6048,n10807,n6050 );
   nand U6283 ( n6052,datao_reg_19_,n6016 );
   nand U6284 ( n6051,n10807,n6053 );
   nand U6285 ( n6055,datao_reg_18_,n6016 );
   nand U6286 ( n6054,n5442,n6056 );
   nand U6287 ( n6058,datao_reg_17_,n6016 );
   nand U6288 ( n6057,n5442,n6059 );
   nand U6289 ( n6061,datao_reg_16_,n6016 );
   nand U6290 ( n6060,n10807,n6062 );
   nand U6291 ( n6064,datao_reg_15_,n6016 );
   nand U6292 ( n6063,n10807,n6065 );
   nand U6293 ( n6067,datao_reg_14_,n6016 );
   nand U6294 ( n6066,n5442,n6068 );
   nand U6295 ( n6070,datao_reg_13_,n6016 );
   nand U6296 ( n6069,n5442,n6071 );
   nand U6297 ( n6073,datao_reg_12_,n6016 );
   nand U6298 ( n6072,n10807,n6074 );
   nand U6299 ( n6076,datao_reg_11_,n6016 );
   nand U6300 ( n6075,n10807,n6077 );
   nand U6301 ( n6079,datao_reg_10_,n6016 );
   nand U6302 ( n6078,n5442,n6080 );
   nand U6303 ( n6082,datao_reg_9_,n6016 );
   nand U6304 ( n6081,n5442,n6083 );
   nand U6305 ( n6085,datao_reg_8_,n6016 );
   nand U6306 ( n6084,n10807,n6086 );
   nand U6307 ( n6088,datao_reg_7_,n6016 );
   nand U6308 ( n6087,n10807,n6089 );
   nand U6309 ( n6091,datao_reg_6_,n6016 );
   nand U6310 ( n6090,n5442,n6092 );
   nand U6311 ( n6094,datao_reg_5_,n6016 );
   nand U6312 ( n6093,n5442,n6095 );
   nand U6313 ( n6097,datao_reg_4_,n6016 );
   nand U6314 ( n6096,n10807,n6098 );
   nand U6315 ( n6100,datao_reg_3_,n6016 );
   nand U6316 ( n6099,n10807,n6101 );
   nand U6317 ( n6103,datao_reg_2_,n6016 );
   nand U6318 ( n6102,n5442,n6104 );
   nand U6319 ( n6106,datao_reg_1_,n5936 );
   nand U6320 ( n6105,n10807,n6107 );
   nand U6321 ( n6109,datao_reg_0_,n6016 );
   nand U6322 ( n6108,n10807,n6110 );
   nand U6323 ( n6112,n5941,n6114 );
   nand U6324 ( n6111,reg1_reg_31_,n5933 );
   nand U6325 ( n6117,reg1_reg_30_,n5933 );
   nand U6326 ( n6116,n5941,n6118 );
   nand U6327 ( n6120,reg1_reg_29_,n5933 );
   nand U6328 ( n6119,n5941,n6121 );
   nand U6329 ( n6123,reg1_reg_28_,n6115 );
   nand U6330 ( n6122,n5941,n6124 );
   nand U6331 ( n6126,reg1_reg_27_,n5933 );
   nand U6332 ( n6125,n5941,n6127 );
   nand U6333 ( n6129,reg1_reg_26_,n5933 );
   nand U6334 ( n6128,n5941,n6130 );
   nand U6335 ( n6132,reg1_reg_25_,n5933 );
   nand U6336 ( n6131,n5941,n6133 );
   nand U6337 ( n6135,reg1_reg_24_,n6115 );
   nand U6338 ( n6134,n5941,n6136 );
   nand U6339 ( n6138,reg1_reg_23_,n5933 );
   nand U6340 ( n6137,n5941,n6139 );
   nand U6341 ( n6141,reg1_reg_22_,n5933 );
   nand U6342 ( n6140,n5941,n6142 );
   nand U6343 ( n6144,reg1_reg_21_,n5933 );
   nand U6344 ( n6143,n5941,n6145 );
   nand U6345 ( n6147,reg1_reg_20_,n5933 );
   nand U6346 ( n6146,n5941,n6148 );
   nand U6347 ( n6150,reg1_reg_19_,n5933 );
   nand U6348 ( n6149,n5941,n6151 );
   nand U6349 ( n6153,reg1_reg_18_,n6115 );
   nand U6350 ( n6152,n5941,n6154 );
   nand U6351 ( n6156,reg1_reg_17_,n6115 );
   nand U6352 ( n6155,n5941,n6157 );
   nand U6353 ( n6159,reg1_reg_16_,n5933 );
   nand U6354 ( n6158,n5941,n6160 );
   nand U6355 ( n6162,reg1_reg_15_,n6115 );
   nand U6356 ( n6161,n5941,n6163 );
   nand U6357 ( n6165,reg1_reg_14_,n6115 );
   nand U6358 ( n6164,n6113,n6166 );
   nand U6359 ( n6168,reg1_reg_13_,n6115 );
   nand U6360 ( n6167,n6113,n6169 );
   nand U6361 ( n6171,reg1_reg_12_,n6115 );
   nand U6362 ( n6170,n6113,n6172 );
   nand U6363 ( n6174,reg1_reg_11_,n6115 );
   nand U6364 ( n6173,n6113,n6175 );
   nand U6365 ( n6177,reg1_reg_10_,n6115 );
   nand U6366 ( n6176,n6113,n6178 );
   nand U6367 ( n6180,reg1_reg_9_,n6115 );
   nand U6368 ( n6179,n6113,n6181 );
   nand U6369 ( n6183,reg1_reg_8_,n6115 );
   nand U6370 ( n6182,n6113,n6184 );
   nand U6371 ( n6186,reg1_reg_7_,n6115 );
   nand U6372 ( n6185,n6113,n6187 );
   nand U6373 ( n6189,reg1_reg_6_,n6115 );
   nand U6374 ( n6188,n6113,n6190 );
   nand U6375 ( n6192,reg1_reg_5_,n6115 );
   nand U6376 ( n6191,n6113,n6193 );
   nand U6377 ( n6195,reg1_reg_4_,n6115 );
   nand U6378 ( n6194,n6113,n6196 );
   nand U6379 ( n6198,reg1_reg_3_,n6115 );
   nand U6380 ( n6197,n6113,n6199 );
   nand U6381 ( n6201,reg1_reg_2_,n6115 );
   nand U6382 ( n6200,n6113,n6202 );
   nand U6383 ( n6204,reg1_reg_1_,n6115 );
   nand U6384 ( n6203,n6113,n6205 );
   nand U6385 ( n6207,reg1_reg_0_,n5933 );
   nand U6386 ( n6206,n6113,n6208 );
   not U6387 ( n6113,n6115 );
   nand U6388 ( n6115,n6209,n6210 );
   nor U6389 ( n6209,n6211,n6212 );
   nand U6390 ( n6214,n5942,n6114 );
   nand U6391 ( n6114,n6216,n6217 );
   nand U6392 ( n6217,n6218,n6219 );
   nor U6393 ( n6216,n6220,n6221 );
   nor U6394 ( n6221,n6222,n6223 );
   nand U6395 ( n6213,reg0_reg_31_,n5934 );
   nand U6396 ( n6226,n5942,n6118 );
   nand U6397 ( n6118,n6227,n6228 );
   nand U6398 ( n6228,n6229,n6218 );
   nor U6399 ( n6227,n6220,n6230 );
   nor U6400 ( n6230,n6223,n6231 );
   nand U6401 ( n6225,reg0_reg_30_,n5934 );
   nand U6402 ( n6233,n5942,n6121 );
   nand U6403 ( n6121,n6234,n6235 );
   nor U6404 ( n6235,n6236,n6237 );
   nor U6405 ( n6237,n6223,n6238 );
   nor U6406 ( n6236,n6239,n6240 );
   nor U6407 ( n6234,n6241,n6242 );
   nor U6408 ( n6241,n6243,n6244 );
   nand U6409 ( n6232,reg0_reg_29_,n5934 );
   nand U6410 ( n6246,n5942,n6124 );
   nand U6411 ( n6124,n6247,n6248 );
   nor U6412 ( n6248,n6249,n6250 );
   nand U6413 ( n6250,n6251,n6252 );
   nand U6414 ( n6252,n6253,n5997 );
   nand U6415 ( n6251,n6255,n6256 );
   nor U6416 ( n6249,n6257,n5943 );
   nor U6417 ( n6247,n6259,n6260 );
   nor U6418 ( n6259,n6012,n6261 );
   nand U6419 ( n6245,reg0_reg_28_,n6224 );
   nand U6420 ( n6263,n5942,n6127 );
   nand U6421 ( n6127,n6264,n6265 );
   nor U6422 ( n6265,n6266,n6267 );
   nand U6423 ( n6267,n6268,n6269 );
   nand U6424 ( n6269,n6270,n5994 );
   nand U6425 ( n6268,n6271,n5997 );
   nor U6426 ( n6266,n6272,n5944 );
   nor U6427 ( n6264,n6273,n6274 );
   nor U6428 ( n6273,n6243,n6275 );
   nand U6429 ( n6262,reg0_reg_27_,n5934 );
   nand U6430 ( n6277,n5942,n6130 );
   nand U6431 ( n6130,n6278,n6279 );
   nor U6432 ( n6279,n6280,n6281 );
   nand U6433 ( n6281,n6282,n6283 );
   nand U6434 ( n6283,n6284,n5997 );
   nand U6435 ( n6282,n6285,n6255 );
   nor U6436 ( n6280,n6286,n5943 );
   nor U6437 ( n6278,n6287,n6288 );
   nor U6438 ( n6287,n6013,n6289 );
   nand U6439 ( n6276,reg0_reg_26_,n5934 );
   nand U6440 ( n6291,n5942,n6133 );
   nand U6441 ( n6133,n6292,n6293 );
   nor U6442 ( n6293,n6294,n6295 );
   nand U6443 ( n6295,n6296,n6297 );
   nand U6444 ( n6297,n6298,n5994 );
   nand U6445 ( n6296,n6299,n5997 );
   nor U6446 ( n6294,n6300,n5944 );
   nor U6447 ( n6292,n6301,n6302 );
   nor U6448 ( n6301,n6012,n6303 );
   nand U6449 ( n6290,reg0_reg_25_,n5934 );
   nand U6450 ( n6305,n5942,n6136 );
   nand U6451 ( n6136,n6306,n6307 );
   nor U6452 ( n6307,n6308,n6309 );
   nand U6453 ( n6309,n6310,n6311 );
   nand U6454 ( n6311,n6312,n5997 );
   nand U6455 ( n6310,n6255,n6313 );
   nor U6456 ( n6308,n6314,n5944 );
   nor U6457 ( n6306,n6315,n6316 );
   nor U6458 ( n6315,n6012,n6317 );
   nand U6459 ( n6304,reg0_reg_24_,n6224 );
   nand U6460 ( n6319,n5942,n6139 );
   nand U6461 ( n6139,n6320,n6321 );
   nor U6462 ( n6321,n6322,n6323 );
   nand U6463 ( n6323,n6324,n6325 );
   nand U6464 ( n6325,n6255,n6326 );
   nand U6465 ( n6324,n6327,n5997 );
   nor U6466 ( n6322,n6328,n6258 );
   nor U6467 ( n6320,n6329,n6330 );
   nor U6468 ( n6329,n6243,n6331 );
   nand U6469 ( n6318,reg0_reg_23_,n5934 );
   nand U6470 ( n6333,n5942,n6142 );
   nand U6471 ( n6142,n6334,n6335 );
   nor U6472 ( n6335,n6336,n6337 );
   nand U6473 ( n6337,n6338,n6339 );
   nand U6474 ( n6339,n6340,n6254 );
   nand U6475 ( n6338,n6341,n6255 );
   nor U6476 ( n6336,n6342,n5943 );
   nor U6477 ( n6334,n6343,n6344 );
   nor U6478 ( n6343,n6013,n6345 );
   nand U6479 ( n6332,reg0_reg_22_,n5934 );
   nand U6480 ( n6347,n5942,n6145 );
   nand U6481 ( n6145,n6348,n6349 );
   nor U6482 ( n6349,n6350,n6351 );
   nand U6483 ( n6351,n6352,n6353 );
   nand U6484 ( n6353,n6354,n5997 );
   nand U6485 ( n6352,n6355,n5994 );
   nor U6486 ( n6350,n6356,n5944 );
   nor U6487 ( n6348,n6357,n6358 );
   nor U6488 ( n6357,n6012,n6359 );
   nand U6489 ( n6346,reg0_reg_21_,n5934 );
   nand U6490 ( n6361,n5942,n6148 );
   nand U6491 ( n6148,n6362,n6363 );
   nor U6492 ( n6363,n6364,n6365 );
   nand U6493 ( n6365,n6366,n6367 );
   nand U6494 ( n6367,n6368,n5997 );
   nand U6495 ( n6366,n6369,n6255 );
   nor U6496 ( n6364,n6370,n6258 );
   nor U6497 ( n6362,n6371,n6372 );
   nor U6498 ( n6371,n6243,n6373 );
   nand U6499 ( n6360,reg0_reg_20_,n5934 );
   nand U6500 ( n6375,n5942,n6151 );
   nand U6501 ( n6151,n6376,n6377 );
   nor U6502 ( n6377,n6378,n6379 );
   nand U6503 ( n6379,n6380,n6381 );
   nand U6504 ( n6381,n6254,n6382 );
   nand U6505 ( n6380,n6255,n6383 );
   nor U6506 ( n6378,n6384,n5943 );
   nor U6507 ( n6376,n6385,n6386 );
   nor U6508 ( n6385,n6013,n6387 );
   nand U6509 ( n6374,reg0_reg_19_,n5934 );
   nand U6510 ( n6389,n5942,n6154 );
   nand U6511 ( n6154,n6390,n6391 );
   nor U6512 ( n6391,n6392,n6393 );
   nand U6513 ( n6393,n6394,n6395 );
   nand U6514 ( n6395,n6396,n5997 );
   nand U6515 ( n6394,n6397,n5994 );
   nor U6516 ( n6392,n6398,n5944 );
   nor U6517 ( n6390,n6399,n6400 );
   nor U6518 ( n6399,n6012,n6401 );
   nand U6519 ( n6388,reg0_reg_18_,n6224 );
   nand U6520 ( n6403,n5942,n6157 );
   nand U6521 ( n6157,n6404,n6405 );
   nor U6522 ( n6405,n6406,n6407 );
   nand U6523 ( n6407,n6408,n6409 );
   nand U6524 ( n6409,n6254,n6410 );
   nand U6525 ( n6408,n6411,n6255 );
   nor U6526 ( n6406,n6412,n6258 );
   nor U6527 ( n6404,n6413,n6414 );
   nor U6528 ( n6413,n6243,n6415 );
   nand U6529 ( n6402,reg0_reg_17_,n6224 );
   nand U6530 ( n6417,n5942,n6160 );
   nand U6531 ( n6160,n6418,n6419 );
   nor U6532 ( n6419,n6420,n6421 );
   nand U6533 ( n6421,n6422,n6423 );
   nand U6534 ( n6423,n6424,n5997 );
   nand U6535 ( n6422,n6425,n6255 );
   nor U6536 ( n6420,n6426,n5943 );
   nor U6537 ( n6418,n6427,n6428 );
   nor U6538 ( n6427,n6013,n6429 );
   nand U6539 ( n6416,reg0_reg_16_,n5934 );
   nand U6540 ( n6431,n5942,n6163 );
   nand U6541 ( n6163,n6432,n6433 );
   nor U6542 ( n6433,n6434,n6435 );
   nand U6543 ( n6435,n6436,n6437 );
   nand U6544 ( n6437,n6254,n6438 );
   nand U6545 ( n6436,n6255,n6439 );
   nor U6546 ( n6434,n6440,n5944 );
   nor U6547 ( n6432,n6441,n6442 );
   nor U6548 ( n6441,n6013,n6443 );
   nand U6549 ( n6430,reg0_reg_15_,n6224 );
   nand U6550 ( n6445,n6215,n6166 );
   nand U6551 ( n6166,n6446,n6447 );
   nor U6552 ( n6447,n6448,n6449 );
   nand U6553 ( n6449,n6450,n6451 );
   nand U6554 ( n6451,n6452,n6254 );
   nand U6555 ( n6450,n6453,n6255 );
   nor U6556 ( n6448,n6454,n6258 );
   nor U6557 ( n6446,n6455,n6456 );
   nor U6558 ( n6455,n6013,n6457 );
   nand U6559 ( n6444,reg0_reg_14_,n6224 );
   nand U6560 ( n6459,n6215,n6169 );
   nand U6561 ( n6169,n6460,n6461 );
   nor U6562 ( n6461,n6462,n6463 );
   nand U6563 ( n6463,n6464,n6465 );
   nand U6564 ( n6465,n6254,n6466 );
   nand U6565 ( n6464,n6467,n6255 );
   nor U6566 ( n6462,n6468,n6258 );
   nor U6567 ( n6460,n6469,n6470 );
   nor U6568 ( n6469,n6243,n6471 );
   nand U6569 ( n6458,reg0_reg_13_,n6224 );
   nand U6570 ( n6473,n6215,n6172 );
   nand U6571 ( n6172,n6474,n6475 );
   nor U6572 ( n6475,n6476,n6477 );
   nand U6573 ( n6477,n6478,n6479 );
   nand U6574 ( n6479,n6480,n5997 );
   nand U6575 ( n6478,n6481,n6255 );
   nor U6576 ( n6476,n6482,n6258 );
   nor U6577 ( n6474,n6483,n6484 );
   nor U6578 ( n6483,n6012,n6485 );
   nand U6579 ( n6472,reg0_reg_12_,n6224 );
   nand U6580 ( n6487,n6215,n6175 );
   nand U6581 ( n6175,n6488,n6489 );
   nor U6582 ( n6489,n6490,n6491 );
   nand U6583 ( n6491,n6492,n6493 );
   nand U6584 ( n6493,n6254,n6494 );
   nand U6585 ( n6492,n6495,n6255 );
   nor U6586 ( n6490,n6496,n6258 );
   nor U6587 ( n6488,n6497,n6498 );
   nor U6588 ( n6497,n6012,n6499 );
   nand U6589 ( n6486,reg0_reg_11_,n6224 );
   nand U6590 ( n6501,n6215,n6178 );
   nand U6591 ( n6178,n6502,n6503 );
   nor U6592 ( n6503,n6504,n6505 );
   nand U6593 ( n6505,n6506,n6507 );
   nand U6594 ( n6507,n6508,n5997 );
   nand U6595 ( n6506,n6509,n5994 );
   nor U6596 ( n6504,n6510,n5943 );
   nor U6597 ( n6502,n6511,n6512 );
   nor U6598 ( n6511,n6243,n6513 );
   nand U6599 ( n6500,reg0_reg_10_,n6224 );
   nand U6600 ( n6515,n6215,n6181 );
   nand U6601 ( n6181,n6516,n6517 );
   nor U6602 ( n6517,n6518,n6519 );
   nand U6603 ( n6519,n6520,n6521 );
   nand U6604 ( n6521,n6254,n6522 );
   nand U6605 ( n6520,n6523,n6255 );
   nor U6606 ( n6518,n6524,n5944 );
   nor U6607 ( n6516,n6525,n6526 );
   nor U6608 ( n6525,n6013,n6527 );
   nand U6609 ( n6514,reg0_reg_9_,n6224 );
   nand U6610 ( n6529,n6215,n6184 );
   nand U6611 ( n6184,n6530,n6531 );
   nor U6612 ( n6531,n6532,n6533 );
   nand U6613 ( n6533,n6534,n6535 );
   nand U6614 ( n6535,n6536,n5997 );
   nand U6615 ( n6534,n6537,n6255 );
   nor U6616 ( n6532,n6538,n6258 );
   nor U6617 ( n6530,n6539,n6540 );
   nor U6618 ( n6539,n6012,n6541 );
   nand U6619 ( n6528,reg0_reg_8_,n6224 );
   nand U6620 ( n6543,n6215,n6187 );
   nand U6621 ( n6187,n6544,n6545 );
   nor U6622 ( n6545,n6546,n6547 );
   nand U6623 ( n6547,n6548,n6549 );
   nand U6624 ( n6549,n6254,n6550 );
   nand U6625 ( n6548,n6551,n6255 );
   nor U6626 ( n6546,n6552,n5943 );
   nor U6627 ( n6544,n6553,n6554 );
   nor U6628 ( n6553,n6243,n6555 );
   nand U6629 ( n6542,reg0_reg_7_,n6224 );
   nand U6630 ( n6557,n6215,n6190 );
   nand U6631 ( n6190,n6558,n6559 );
   nor U6632 ( n6559,n6560,n6561 );
   nand U6633 ( n6561,n6562,n6563 );
   nand U6634 ( n6563,n6564,n5997 );
   nand U6635 ( n6562,n6565,n6255 );
   nor U6636 ( n6560,n6566,n5944 );
   nor U6637 ( n6558,n6567,n6568 );
   nor U6638 ( n6567,n6013,n6569 );
   nand U6639 ( n6556,reg0_reg_6_,n6224 );
   nand U6640 ( n6571,n6215,n6193 );
   nand U6641 ( n6193,n6572,n6573 );
   nor U6642 ( n6573,n6574,n6575 );
   nand U6643 ( n6575,n6576,n6577 );
   nand U6644 ( n6577,n6254,n6578 );
   nand U6645 ( n6576,n6579,n6255 );
   nor U6646 ( n6574,n6580,n6258 );
   nor U6647 ( n6572,n6581,n6582 );
   nor U6648 ( n6581,n6012,n6583 );
   nand U6649 ( n6570,reg0_reg_5_,n6224 );
   nand U6650 ( n6585,n6215,n6196 );
   nand U6651 ( n6196,n6586,n6587 );
   nor U6652 ( n6587,n6588,n6589 );
   nand U6653 ( n6589,n6590,n6591 );
   nand U6654 ( n6591,n6592,n5997 );
   nand U6655 ( n6590,n6593,n6255 );
   nor U6656 ( n6588,n6594,n5943 );
   nor U6657 ( n6586,n6595,n6596 );
   nor U6658 ( n6595,n6243,n6597 );
   nand U6659 ( n6584,reg0_reg_4_,n6224 );
   nand U6660 ( n6599,n6215,n6199 );
   nand U6661 ( n6199,n6600,n6601 );
   nor U6662 ( n6601,n6602,n6603 );
   nand U6663 ( n6603,n6604,n6605 );
   nand U6664 ( n6605,n6254,n6606 );
   nand U6665 ( n6604,n6607,n5994 );
   nor U6666 ( n6602,n6608,n5944 );
   nor U6667 ( n6600,n6609,n6610 );
   nor U6668 ( n6609,n6013,n6611 );
   nand U6669 ( n6598,reg0_reg_3_,n6224 );
   nand U6670 ( n6613,n6215,n6202 );
   nand U6671 ( n6202,n6614,n6615 );
   nor U6672 ( n6615,n6616,n6617 );
   nand U6673 ( n6617,n6618,n6619 );
   nand U6674 ( n6619,n6620,n5997 );
   nand U6675 ( n6618,n6621,n5994 );
   nor U6676 ( n6616,n6622,n6258 );
   nor U6677 ( n6614,n6623,n6624 );
   nor U6678 ( n6623,n6012,n6625 );
   nand U6679 ( n6612,reg0_reg_2_,n6224 );
   nand U6680 ( n6627,n6215,n6205 );
   nand U6681 ( n6205,n6628,n6629 );
   nor U6682 ( n6629,n6630,n6631 );
   nand U6683 ( n6631,n6632,n6633 );
   nand U6684 ( n6633,n6254,n6634 );
   nand U6685 ( n6632,n6255,n6635 );
   not U6686 ( n6255,n6240 );
   nor U6687 ( n6630,n6636,n5943 );
   nor U6688 ( n6628,n6637,n6638 );
   nor U6689 ( n6637,n6243,n6639 );
   nand U6690 ( n6626,reg0_reg_1_,n6224 );
   nand U6691 ( n6641,n6215,n6208 );
   nand U6692 ( n6208,n6642,n6643 );
   nor U6693 ( n6643,n6644,n6645 );
   nor U6694 ( n6645,n6646,n6647 );
   nor U6695 ( n6646,n6218,n6254 );
   nor U6696 ( n6642,n6648,n6649 );
   nor U6697 ( n6649,n6650,n5943 );
   nor U6698 ( n6648,n6240,n6651 );
   nand U6699 ( n6240,n6652,n6653 );
   not U6700 ( n6215,n6224 );
   nand U6701 ( n6640,reg0_reg_0_,n5934 );
   nand U6702 ( n6224,n6654,n6210 );
   nor U6703 ( n6654,n6655,n6211 );
   nand U6704 ( n6211,n6656,n6657 );
   not U6705 ( n6657,n6658 );
   nor U6706 ( n6656,n6659,n6660 );
   nor U6707 ( n6660,n6661,n6662 );
   or U6708 ( n6662,n6663,n6664 );
   nor U6709 ( n6661,n6665,n6666 );
   nor U6710 ( n6665,n6667,n6668 );
   nand U6711 ( n6670,d_reg_1_,n6671 );
   nand U6712 ( n6669,n5935,n6673 );
   nand U6713 ( n6675,d_reg_0_,n6671 );
   nand U6714 ( n6674,n5935,n6676 );
   nor U6715 ( n6678,n6679,n6680 );
   nand U6716 ( n6680,n6681,n6682 );
   or U6717 ( n6682,n6683,n6684 );
   or U6718 ( n6681,n6685,n6239 );
   xor U6719 ( n6239,n6686,n6687 );
   nor U6720 ( n6686,n6688,n6689 );
   nor U6721 ( n6688,n6690,n6691 );
   nor U6722 ( n6679,n6238,n6692 );
   xor U6723 ( n6238,n6693,n6694 );
   nor U6724 ( n6677,n6695,n6696 );
   nand U6725 ( n6696,n6697,n6698 );
   nand U6726 ( n6698,reg2_reg_29_,n6002 );
   nand U6727 ( n6697,n6700,n6242 );
   nand U6728 ( n6242,n6701,n6702 );
   nor U6729 ( n6702,n6703,n6704 );
   nor U6730 ( n6704,n6705,n6706 );
   nand U6731 ( n6706,n6707,n6708 );
   nand U6732 ( n6708,n6709,n6710 );
   nor U6733 ( n6709,n6711,n6712 );
   nor U6734 ( n6712,n6713,n6714 );
   nand U6735 ( n6707,n6715,n6687 );
   nor U6736 ( n6715,n6713,n6716 );
   nor U6737 ( n6716,n6711,n6717 );
   nor U6738 ( n6703,n6718,n6719 );
   xor U6739 ( n6719,n6720,n6710 );
   not U6740 ( n6710,n6687 );
   nand U6741 ( n6720,n6721,n6722 );
   nand U6742 ( n6722,n6723,n6724 );
   not U6743 ( n6724,n6690 );
   not U6744 ( n6721,n6689 );
   nor U6745 ( n6701,n6725,n6726 );
   nor U6746 ( n6726,n6727,n6728 );
   nor U6747 ( n6725,n6272,n6729 );
   nor U6748 ( n6695,n6244,n6730 );
   nand U6749 ( n6732,ir_reg_0_,n6733 );
   nand U6750 ( n6733,n6734,n5946 );
   nand U6751 ( n6731,datai_0_,n5973 );
   nand U6752 ( n6736,datai_1_,n5973 );
   nor U6753 ( n6735,n6737,n6738 );
   nor U6754 ( n6738,ir_reg_1_,n6739 );
   nand U6755 ( n6739,n6740,ir_reg_0_ );
   nor U6756 ( n6737,n6741,n6742 );
   nor U6757 ( n6741,n6743,n6744 );
   nor U6758 ( n6743,ir_reg_0_,n5948 );
   nand U6759 ( n6746,datai_2_,n5973 );
   nor U6760 ( n6745,n6747,n6748 );
   nor U6761 ( n6748,n6749,n6734 );
   nor U6762 ( n6747,n5948,n6750 );
   nand U6763 ( n6752,datai_3_,n5932 );
   nor U6764 ( n6751,n6753,n6754 );
   and U6765 ( n6754,ir_reg_3_,n5451 );
   nor U6766 ( n6753,n5947,n6755 );
   nand U6767 ( n6755,n6756,n6757 );
   nand U6768 ( n6759,datai_4_,n5975 );
   nor U6769 ( n6758,n6760,n6761 );
   nor U6770 ( n6761,ir_reg_4_,n6762 );
   nand U6771 ( n6762,n6740,n6757 );
   nor U6772 ( n6760,n6763,n6764 );
   nor U6773 ( n6763,n6765,n5451 );
   nor U6774 ( n6765,n6757,n5948 );
   nand U6775 ( n6767,datai_5_,n5932 );
   nor U6776 ( n6766,n6768,n6769 );
   nor U6777 ( n6769,n6770,n6734 );
   nor U6778 ( n6768,n5947,n6771 );
   nand U6779 ( n6773,datai_6_,n5932 );
   nor U6780 ( n6772,n6774,n6775 );
   nor U6781 ( n6775,ir_reg_6_,n6776 );
   nand U6782 ( n6776,n6740,n6777 );
   nor U6783 ( n6774,n6778,n6779 );
   nor U6784 ( n6778,n6780,n5451 );
   nor U6785 ( n6780,n6777,n5948 );
   nand U6786 ( n6782,datai_7_,n5973 );
   nor U6787 ( n6781,n6783,n6784 );
   nor U6788 ( n6784,n6785,n6734 );
   nor U6789 ( n6783,n5947,n6786 );
   nand U6790 ( n6788,datai_8_,n5975 );
   nor U6791 ( n6787,n6789,n6790 );
   nor U6792 ( n6790,ir_reg_8_,n6791 );
   nand U6793 ( n6791,n6740,n6792 );
   nor U6794 ( n6789,n6793,n6794 );
   nor U6795 ( n6793,n6795,n5451 );
   nor U6796 ( n6795,n6792,n5947 );
   nand U6797 ( n6797,datai_9_,n5975 );
   nor U6798 ( n6796,n6798,n6799 );
   nor U6799 ( n6799,n6800,n6734 );
   nor U6800 ( n6798,n5947,n6801 );
   nand U6801 ( n6803,datai_10_,n5932 );
   nor U6802 ( n6802,n6804,n6805 );
   nor U6803 ( n6805,ir_reg_10_,n6806 );
   nand U6804 ( n6806,n6740,n6807 );
   nor U6805 ( n6804,n6808,n6809 );
   not U6806 ( n6809,ir_reg_10_ );
   nor U6807 ( n6808,n6810,n6744 );
   nor U6808 ( n6810,n6807,n5946 );
   nand U6809 ( n6812,datai_11_,n5932 );
   nor U6810 ( n6811,n6813,n6814 );
   nor U6811 ( n6814,n6815,n6734 );
   nor U6812 ( n6813,n5946,n6816 );
   nand U6813 ( n6818,datai_12_,n5973 );
   nor U6814 ( n6817,n6819,n6820 );
   nor U6815 ( n6820,ir_reg_12_,n6821 );
   nand U6816 ( n6821,n6740,n6822 );
   nor U6817 ( n6819,n6823,n6824 );
   not U6818 ( n6824,ir_reg_12_ );
   nor U6819 ( n6823,n6825,n6744 );
   nor U6820 ( n6825,n6822,n5946 );
   nand U6821 ( n6827,datai_13_,n5975 );
   nor U6822 ( n6826,n6828,n6829 );
   nor U6823 ( n6829,n6830,n6734 );
   nor U6824 ( n6828,n5946,n6831 );
   nand U6825 ( n6833,datai_14_,n5932 );
   nor U6826 ( n6832,n6834,n6835 );
   nor U6827 ( n6835,ir_reg_14_,n6836 );
   nand U6828 ( n6836,n6740,n6837 );
   nor U6829 ( n6834,n6838,n6839 );
   not U6830 ( n6839,ir_reg_14_ );
   nor U6831 ( n6838,n6840,n6744 );
   nor U6832 ( n6840,n6837,n5947 );
   nand U6833 ( n6842,datai_15_,n5973 );
   nor U6834 ( n6841,n6843,n6844 );
   nor U6835 ( n6844,n6845,n6734 );
   nor U6836 ( n6843,n5946,n6846 );
   nand U6837 ( n6848,datai_16_,n5975 );
   nor U6838 ( n6847,n6849,n6850 );
   nor U6839 ( n6850,ir_reg_16_,n6851 );
   nand U6840 ( n6851,n6740,n6852 );
   nor U6841 ( n6849,n6853,n6854 );
   not U6842 ( n6854,ir_reg_16_ );
   nor U6843 ( n6853,n6855,n6744 );
   nor U6844 ( n6855,n6852,n5948 );
   nand U6845 ( n6857,datai_17_,n5975 );
   nor U6846 ( n6856,n6858,n6859 );
   nor U6847 ( n6859,n6860,n6734 );
   nor U6848 ( n6858,n5946,n6861 );
   nand U6849 ( n6863,datai_18_,n5975 );
   nor U6850 ( n6862,n6864,n6865 );
   nor U6851 ( n6865,ir_reg_18_,n6866 );
   nand U6852 ( n6866,n6740,n6867 );
   nor U6853 ( n6864,n6868,n6869 );
   not U6854 ( n6869,ir_reg_18_ );
   nor U6855 ( n6868,n6870,n6744 );
   nor U6856 ( n6870,n6867,n5946 );
   nand U6857 ( n6872,datai_19_,n5975 );
   nor U6858 ( n6871,n6873,n6874 );
   nor U6859 ( n6874,n6875,n6734 );
   nor U6860 ( n6873,n5948,n6876 );
   nand U6861 ( n6878,datai_20_,n5975 );
   nor U6862 ( n6877,n6879,n6880 );
   nor U6863 ( n6880,ir_reg_20_,n6881 );
   nand U6864 ( n6881,n6740,n6882 );
   nor U6865 ( n6879,n6883,n6884 );
   not U6866 ( n6884,ir_reg_20_ );
   nor U6867 ( n6883,n6885,n6744 );
   nor U6868 ( n6885,n6882,n5948 );
   nand U6869 ( n6887,datai_21_,n5932 );
   nor U6870 ( n6886,n6888,n6889 );
   nor U6871 ( n6889,n6890,n6734 );
   nor U6872 ( n6888,n5946,n6891 );
   nand U6873 ( n6893,datai_22_,n5932 );
   nor U6874 ( n6892,n6894,n6895 );
   nor U6875 ( n6895,ir_reg_22_,n6896 );
   nand U6876 ( n6896,n6740,n6897 );
   nor U6877 ( n6894,n6898,n6899 );
   not U6878 ( n6899,ir_reg_22_ );
   nor U6879 ( n6898,n6900,n5451 );
   nor U6880 ( n6900,n6897,n5946 );
   nand U6881 ( n6902,datai_23_,n5932 );
   nor U6882 ( n6901,n6903,n6904 );
   nor U6883 ( n6904,n6905,n6734 );
   nor U6884 ( n6903,n5947,n6906 );
   nand U6885 ( n6908,datai_24_,n5975 );
   nor U6886 ( n6907,n6909,n6910 );
   nor U6887 ( n6910,ir_reg_24_,n6911 );
   nand U6888 ( n6911,n6740,n6912 );
   nor U6889 ( n6909,n6913,n6914 );
   not U6890 ( n6914,ir_reg_24_ );
   nor U6891 ( n6913,n6915,n6744 );
   nor U6892 ( n6915,n6912,n5947 );
   nand U6893 ( n6917,datai_25_,n5975 );
   nor U6894 ( n6916,n6918,n6919 );
   nor U6895 ( n6919,n6920,n6734 );
   nor U6896 ( n6918,n5947,n6921 );
   nand U6897 ( n6923,datai_26_,n5973 );
   nor U6898 ( n6922,n6924,n6925 );
   and U6899 ( n6925,ir_reg_26_,n5451 );
   nor U6900 ( n6924,n5948,n6926 );
   nand U6901 ( n6926,n6927,n6928 );
   nand U6902 ( n6930,datai_27_,n5975 );
   nor U6903 ( n6929,n6931,n6932 );
   nor U6904 ( n6932,ir_reg_27_,n6933 );
   nand U6905 ( n6933,n6740,n6928 );
   nor U6906 ( n6931,n6934,n6935 );
   nor U6907 ( n6934,n6936,n6744 );
   nor U6908 ( n6936,n6928,n5947 );
   not U6909 ( n6928,n6937 );
   nand U6910 ( n6939,datai_28_,n5975 );
   nor U6911 ( n6938,n6940,n6941 );
   nor U6912 ( n6941,n6942,n5448 );
   nor U6913 ( n6940,n5948,n6943 );
   nand U6914 ( n6945,datai_29_,n5932 );
   nor U6915 ( n6944,n6946,n6947 );
   nor U6916 ( n6947,ir_reg_29_,n6948 );
   nand U6917 ( n6948,n6740,n6949 );
   nor U6918 ( n6946,n6950,n6951 );
   nor U6919 ( n6950,n6952,n6744 );
   nor U6920 ( n6952,n6949,n5946 );
   nand U6921 ( n6954,datai_30_,n5973 );
   nor U6922 ( n6953,n6955,n6956 );
   nor U6923 ( n6956,n6957,n6734 );
   not U6924 ( n6734,n6744 );
   nor U6925 ( n6955,n5948,n6958 );
   or U6926 ( n6960,n6961,n5947 );
   nor U6927 ( n6740,n6744,n5973 );
   nor U6928 ( n6744,n5975,ir_reg_31_ );
   nand U6929 ( n6959,datai_31_,n5932 );
   nor U6930 ( n10797,n6672,n6968 );
   nor U6931 ( n10798,n5935,n6970 );
   nor U6932 ( n10799,n6672,n6971 );
   nor U6933 ( n10800,n6672,n6972 );
   nor U6934 ( n10801,n5935,n6973 );
   nor U6935 ( n10802,n5935,n6974 );
   not U6936 ( n6671,n5935 );
   nor U6937 ( n10803,n5935,n6975 );
   nor U6938 ( n10804,n6672,n6976 );
   nor U6939 ( n10805,n5935,n6977 );
   nor U6940 ( n10806,n6672,n6978 );
   nor U6941 ( n6672,n6979,n6980 );
   nor U6942 ( n6982,n6983,n6984 );
   nand U6943 ( n6984,n6985,n6986 );
   nand U6944 ( n6986,n6987,n6988 );
   nand U6945 ( n6988,n6692,n6730 );
   nand U6946 ( n6985,n6989,n6107 );
   nor U6947 ( n6983,n6651,n6685 );
   not U6948 ( n6685,n6990 );
   nor U6949 ( n6981,n6991,n6992 );
   nand U6950 ( n6992,n6993,n6994 );
   nand U6951 ( n6994,reg2_reg_0_,n6699 );
   nand U6952 ( n6993,n6644,n5989 );
   nor U6953 ( n6644,n6651,n6995 );
   and U6954 ( n6995,n5999,n5986 );
   nor U6955 ( n6991,n6996,n6683 );
   nor U6956 ( n6998,n6999,n7000 );
   nand U6957 ( n7000,n7001,n7002 );
   nand U6958 ( n7002,n7003,n6634 );
   xor U6959 ( n6634,n6647,n6639 );
   nand U6960 ( n7001,n6990,n6635 );
   nor U6961 ( n6999,n6636,n7004 );
   nor U6962 ( n6997,n7005,n7006 );
   nand U6963 ( n7006,n7007,n7008 );
   nand U6964 ( n7008,n7009,reg3_reg_1_ );
   nand U6965 ( n7007,n7010,n7011 );
   nand U6966 ( n7005,n7012,n7013 );
   nand U6967 ( n7013,reg2_reg_1_,n6699 );
   nand U6968 ( n7012,n5989,n6638 );
   nand U6969 ( n6638,n7014,n7015 );
   nand U6970 ( n7015,n7016,n6110 );
   nor U6971 ( n7014,n7017,n7018 );
   and U6972 ( n7018,n7019,n6635 );
   xor U6973 ( n6635,n7020,n7021 );
   nor U6974 ( n7017,n5998,n7022 );
   xor U6975 ( n7022,n7023,n7021 );
   nor U6976 ( n7025,n7026,n7027 );
   nand U6977 ( n7027,n7028,n7029 );
   nand U6978 ( n7029,n6620,n7003 );
   nor U6979 ( n6620,n7030,n7031 );
   and U6980 ( n7031,n7032,n7033 );
   nand U6981 ( n7033,n6639,n6647 );
   nand U6982 ( n7028,n5978,n6621 );
   not U6983 ( n6621,n7034 );
   nor U6984 ( n7026,n6622,n7004 );
   nor U6985 ( n7024,n7035,n7036 );
   nand U6986 ( n7036,n7037,n7038 );
   nand U6987 ( n7038,n7009,reg3_reg_2_ );
   nand U6988 ( n7037,n7010,n7032 );
   nand U6989 ( n7035,n7039,n7040 );
   nand U6990 ( n7040,reg2_reg_2_,n6002 );
   nand U6991 ( n7039,n5989,n6624 );
   nand U6992 ( n6624,n7041,n7042 );
   nor U6993 ( n7042,n7043,n7044 );
   nor U6994 ( n7044,n7045,n7046 );
   nand U6995 ( n7046,n7047,n7048 );
   nand U6996 ( n7047,n7049,n7050 );
   not U6997 ( n7050,n7051 );
   nor U6998 ( n7043,n7052,n7053 );
   nand U6999 ( n7053,n7054,n7048 );
   nand U7000 ( n7048,n7055,n7051 );
   nand U7001 ( n7054,n7056,n7057 );
   nor U7002 ( n7052,n7058,n7059 );
   nor U7003 ( n7041,n7060,n7061 );
   nor U7004 ( n7061,n6650,n6729 );
   nor U7005 ( n7060,n6718,n7034 );
   nand U7006 ( n7034,n7062,n7063 );
   nand U7007 ( n7063,n7055,n7064 );
   nand U7008 ( n7062,n7049,n7065 );
   not U7009 ( n7065,n7064 );
   nor U7010 ( n7049,n7066,n7067 );
   nor U7011 ( n7069,n7070,n7071 );
   nand U7012 ( n7071,n7072,n7073 );
   nand U7013 ( n7073,n7003,n6606 );
   xor U7014 ( n6606,n7030,n6611 );
   nand U7015 ( n7072,n6990,n6607 );
   nor U7016 ( n7070,n6608,n6000 );
   nor U7017 ( n7068,n7074,n7075 );
   nand U7018 ( n7075,n7076,n7077 );
   nand U7019 ( n7077,n5976,n7078 );
   nand U7020 ( n7076,n5981,n7079 );
   nand U7021 ( n7074,n7080,n7081 );
   nand U7022 ( n7081,reg2_reg_3_,n6699 );
   nand U7023 ( n7080,n5989,n6610 );
   nand U7024 ( n6610,n7082,n7083 );
   nor U7025 ( n7083,n7084,n7085 );
   nor U7026 ( n7085,n7086,n7087 );
   nand U7027 ( n7087,n7088,n7089 );
   or U7028 ( n7089,n7090,n7056 );
   or U7029 ( n7088,n7091,n7092 );
   nor U7030 ( n7084,n7057,n7093 );
   nand U7031 ( n7093,n7091,n7094 );
   nor U7032 ( n7082,n7095,n7096 );
   nor U7033 ( n7096,n6636,n6729 );
   and U7034 ( n7095,n7019,n6607 );
   xor U7035 ( n6607,n7091,n7097 );
   not U7036 ( n7091,n7090 );
   nor U7037 ( n7099,n7100,n7101 );
   nand U7038 ( n7101,n7102,n7103 );
   nand U7039 ( n7103,n6592,n5977 );
   nor U7040 ( n6592,n7104,n7105 );
   and U7041 ( n7105,n7106,n7107 );
   nand U7042 ( n7107,n7030,n6611 );
   nand U7043 ( n7102,n5978,n6593 );
   not U7044 ( n6593,n7108 );
   nor U7045 ( n7100,n6594,n6000 );
   nor U7046 ( n7098,n7109,n7110 );
   nand U7047 ( n7110,n7111,n7112 );
   nand U7048 ( n7112,n7009,n7113 );
   nand U7049 ( n7111,n7010,n7106 );
   nand U7050 ( n7109,n7114,n7115 );
   nand U7051 ( n7115,reg2_reg_4_,n6002 );
   nand U7052 ( n7114,n5989,n6596 );
   nand U7053 ( n6596,n7116,n7117 );
   nand U7054 ( n7117,n7016,n6101 );
   nor U7055 ( n7116,n7118,n7119 );
   nor U7056 ( n7119,n6705,n7120 );
   nand U7057 ( n7120,n7121,n7122 );
   or U7058 ( n7122,n7123,n7124 );
   nand U7059 ( n7121,n7125,n7124 );
   and U7060 ( n7125,n7126,n7127 );
   nor U7061 ( n7118,n5986,n7108 );
   xor U7062 ( n7108,n7123,n7128 );
   nor U7063 ( n7130,n7131,n7132 );
   nand U7064 ( n7132,n7133,n7134 );
   nand U7065 ( n7134,n7003,n6578 );
   xor U7066 ( n6578,n7104,n6583 );
   nand U7067 ( n7133,n5978,n6579 );
   not U7068 ( n6579,n7135 );
   nor U7069 ( n7131,n6580,n7004 );
   nor U7070 ( n7129,n7136,n7137 );
   nand U7071 ( n7137,n7138,n7139 );
   nand U7072 ( n7139,n5976,n7140 );
   nand U7073 ( n7138,n5981,n7141 );
   nand U7074 ( n7136,n7142,n7143 );
   nand U7075 ( n7143,reg2_reg_5_,n6002 );
   nand U7076 ( n7142,n5989,n6582 );
   nand U7077 ( n6582,n7144,n7145 );
   nand U7078 ( n7145,n7016,n6098 );
   nor U7079 ( n7144,n7146,n7147 );
   nor U7080 ( n7147,n6705,n7148 );
   nand U7081 ( n7148,n7149,n7150 );
   nand U7082 ( n7150,n7151,n7152 );
   nor U7083 ( n7151,n7153,n7154 );
   or U7084 ( n7149,n7155,n7152 );
   nor U7085 ( n7146,n6718,n7135 );
   nand U7086 ( n7135,n7156,n7157 );
   nand U7087 ( n7157,n7158,n7159 );
   nand U7088 ( n7159,n7128,n7160 );
   nor U7089 ( n7158,n7161,n7162 );
   nand U7090 ( n7156,n7163,n7164 );
   nor U7091 ( n7163,n7165,n7166 );
   nor U7092 ( n7166,n7161,n7128 );
   nor U7093 ( n7168,n7169,n7170 );
   nand U7094 ( n7170,n7171,n7172 );
   nand U7095 ( n7172,n6564,n5977 );
   nor U7096 ( n6564,n7173,n7174 );
   and U7097 ( n7174,n7175,n7176 );
   nand U7098 ( n7176,n7104,n6583 );
   nand U7099 ( n7171,n5978,n6565 );
   nor U7100 ( n7169,n6566,n6000 );
   nor U7101 ( n7167,n7177,n7178 );
   nand U7102 ( n7178,n7179,n7180 );
   nand U7103 ( n7180,n5976,n7181 );
   nand U7104 ( n7179,n5981,n7175 );
   nand U7105 ( n7177,n7182,n7183 );
   nand U7106 ( n7183,reg2_reg_6_,n6699 );
   nand U7107 ( n7182,n5989,n6568 );
   nand U7108 ( n6568,n7184,n7185 );
   nor U7109 ( n7185,n7186,n7187 );
   nor U7110 ( n7187,n7188,n7086 );
   nor U7111 ( n7188,n7189,n7190 );
   nor U7112 ( n7190,n7191,n7192 );
   nand U7113 ( n7192,n7193,n7194 );
   nor U7114 ( n7189,n7195,n7193 );
   nand U7115 ( n7193,n7152,n7196 );
   nand U7116 ( n7152,n7127,n7197 );
   nand U7117 ( n7197,n7124,n7126 );
   nor U7118 ( n7186,n7198,n7199 );
   nand U7119 ( n7199,n7200,n7094 );
   nor U7120 ( n7184,n7201,n7202 );
   nor U7121 ( n7202,n6594,n6729 );
   and U7122 ( n7201,n7019,n6565 );
   xor U7123 ( n6565,n7200,n7203 );
   nor U7124 ( n7205,n7206,n7207 );
   nand U7125 ( n7207,n7208,n7209 );
   nand U7126 ( n7209,n7003,n6550 );
   xor U7127 ( n6550,n6555,n7173 );
   nand U7128 ( n7208,n6990,n6551 );
   not U7129 ( n6551,n7210 );
   nor U7130 ( n7206,n6552,n7004 );
   nor U7131 ( n7204,n7211,n7212 );
   nand U7132 ( n7212,n7213,n7214 );
   nand U7133 ( n7214,n5976,n7215 );
   nand U7134 ( n7213,n5981,n7216 );
   nand U7135 ( n7211,n7217,n7218 );
   nand U7136 ( n7218,reg2_reg_7_,n6699 );
   nand U7137 ( n7217,n5989,n6554 );
   nand U7138 ( n6554,n7219,n7220 );
   nor U7139 ( n7220,n7221,n7222 );
   nor U7140 ( n7222,n7045,n7223 );
   nand U7141 ( n7223,n7224,n7225 );
   nand U7142 ( n7225,n7226,n7227 );
   nor U7143 ( n7226,n7228,n7229 );
   or U7144 ( n7224,n7227,n7230 );
   nor U7145 ( n7221,n7231,n7232 );
   nand U7146 ( n7232,n7233,n7234 );
   or U7147 ( n7234,n7235,n7228 );
   not U7148 ( n7233,n7236 );
   nor U7149 ( n7231,n7230,n7227 );
   nor U7150 ( n7219,n7237,n7238 );
   nor U7151 ( n7238,n6580,n6729 );
   nor U7152 ( n7237,n5986,n7210 );
   nand U7153 ( n7210,n7239,n7240 );
   nand U7154 ( n7240,n7241,n7230 );
   nor U7155 ( n7241,n7242,n7243 );
   nand U7156 ( n7239,n7244,n7245 );
   not U7157 ( n7245,n7230 );
   nor U7158 ( n7244,n7246,n7247 );
   nor U7159 ( n7247,n7242,n7203 );
   nor U7160 ( n7249,n7250,n7251 );
   nand U7161 ( n7251,n7252,n7253 );
   nand U7162 ( n7253,n6536,n5977 );
   nor U7163 ( n6536,n7254,n7255 );
   and U7164 ( n7255,n7256,n7257 );
   nand U7165 ( n7257,n7173,n6555 );
   nand U7166 ( n7252,n6990,n6537 );
   nor U7167 ( n7250,n6538,n6000 );
   nor U7168 ( n7248,n7258,n7259 );
   nand U7169 ( n7259,n7260,n7261 );
   nand U7170 ( n7261,n7009,n7262 );
   nand U7171 ( n7260,n7010,n7256 );
   nand U7172 ( n7258,n7263,n7264 );
   nand U7173 ( n7264,reg2_reg_8_,n6002 );
   nand U7174 ( n7263,n5989,n6540 );
   nand U7175 ( n6540,n7265,n7266 );
   nor U7176 ( n7266,n7267,n7268 );
   nor U7177 ( n7268,n7086,n7269 );
   nand U7178 ( n7269,n7270,n7271 );
   nand U7179 ( n7271,n7272,n7235 );
   nand U7180 ( n7270,n7273,n7274 );
   nand U7181 ( n7273,n7235,n7275 );
   nand U7182 ( n7235,n7227,n7276 );
   nand U7183 ( n7227,n7277,n7278 );
   nand U7184 ( n7278,n7124,n7279 );
   not U7185 ( n7124,n7280 );
   nor U7186 ( n7277,n7281,n7282 );
   and U7187 ( n7282,n7194,n7191 );
   not U7188 ( n7281,n7283 );
   nor U7189 ( n7086,n7058,n7284 );
   not U7190 ( n7284,n7285 );
   nor U7191 ( n7267,n7274,n7286 );
   nand U7192 ( n7286,n7228,n7094 );
   nand U7193 ( n7094,n7285,n7287 );
   not U7194 ( n7274,n7272 );
   nor U7195 ( n7265,n7288,n7289 );
   nor U7196 ( n7289,n6566,n6729 );
   and U7197 ( n7288,n7019,n6537 );
   xor U7198 ( n6537,n7290,n7272 );
   nor U7199 ( n7292,n7293,n7294 );
   nand U7200 ( n7294,n7295,n7296 );
   nand U7201 ( n7296,n7003,n6522 );
   xor U7202 ( n6522,n7254,n6527 );
   nand U7203 ( n7295,n6990,n6523 );
   nor U7204 ( n7293,n6524,n7004 );
   nor U7205 ( n7291,n7297,n7298 );
   nand U7206 ( n7298,n7299,n7300 );
   or U7207 ( n7300,n6683,n7301 );
   nand U7208 ( n7299,n7010,n7302 );
   nand U7209 ( n7297,n7303,n7304 );
   nand U7210 ( n7304,reg2_reg_9_,n6699 );
   nand U7211 ( n7303,n5989,n6526 );
   nand U7212 ( n6526,n7305,n7306 );
   nand U7213 ( n7306,n7016,n6086 );
   nor U7214 ( n7305,n7307,n7308 );
   nor U7215 ( n7308,n5999,n7309 );
   nand U7216 ( n7309,n7310,n7311 );
   nand U7217 ( n7311,n7312,n7313 );
   nor U7218 ( n7312,n7314,n7315 );
   nand U7219 ( n7310,n7316,n7317 );
   and U7220 ( n7307,n7019,n6523 );
   xor U7221 ( n6523,n7318,n7316 );
   nor U7222 ( n7320,n7321,n7322 );
   nand U7223 ( n7322,n7323,n7324 );
   nand U7224 ( n7324,n6508,n5977 );
   nor U7225 ( n6508,n7325,n7326 );
   and U7226 ( n7326,n7327,n7328 );
   nand U7227 ( n7328,n7254,n6527 );
   nand U7228 ( n7323,n6990,n6509 );
   not U7229 ( n6509,n7329 );
   nor U7230 ( n7321,n6510,n6000 );
   nor U7231 ( n7319,n7330,n7331 );
   nand U7232 ( n7331,n7332,n7333 );
   nand U7233 ( n7333,n7009,n7334 );
   nand U7234 ( n7332,n7010,n7327 );
   nand U7235 ( n7330,n7335,n7336 );
   nand U7236 ( n7336,reg2_reg_10_,n6002 );
   nand U7237 ( n7335,n5989,n6512 );
   nand U7238 ( n6512,n7337,n7338 );
   nand U7239 ( n7338,n7016,n6083 );
   nor U7240 ( n7337,n7339,n7340 );
   nor U7241 ( n7340,n6705,n7341 );
   nand U7242 ( n7341,n7342,n7343 );
   nand U7243 ( n7343,n7344,n7345 );
   nor U7244 ( n7344,n7346,n7347 );
   nand U7245 ( n7342,n7348,n7349 );
   nor U7246 ( n7339,n6718,n7329 );
   nand U7247 ( n7329,n7350,n7351 );
   nand U7248 ( n7351,n7352,n7353 );
   nand U7249 ( n7353,n7354,n7318 );
   nor U7250 ( n7352,n7355,n7348 );
   nand U7251 ( n7350,n7356,n7357 );
   not U7252 ( n7357,n7358 );
   nor U7253 ( n7356,n7359,n7360 );
   nor U7254 ( n7360,n7355,n7318 );
   nand U7255 ( n7318,n7361,n7362 );
   nand U7256 ( n7362,n7290,n7363 );
   not U7257 ( n7363,n7364 );
   nand U7258 ( n7290,n7365,n7366 );
   nand U7259 ( n7366,n7243,n7367 );
   not U7260 ( n7361,n7368 );
   nor U7261 ( n7370,n7371,n7372 );
   nand U7262 ( n7372,n7373,n7374 );
   nand U7263 ( n7374,n7003,n6494 );
   xor U7264 ( n6494,n6499,n7325 );
   nand U7265 ( n7373,n6990,n6495 );
   not U7266 ( n6495,n7375 );
   nor U7267 ( n7371,n6496,n7004 );
   nor U7268 ( n7369,n7376,n7377 );
   nand U7269 ( n7377,n7378,n7379 );
   nand U7270 ( n7379,n7009,n7380 );
   nand U7271 ( n7378,n7010,n7381 );
   nand U7272 ( n7376,n7382,n7383 );
   nand U7273 ( n7383,reg2_reg_11_,n6699 );
   nand U7274 ( n7382,n5989,n6498 );
   nand U7275 ( n6498,n7384,n7385 );
   nand U7276 ( n7385,n7016,n6080 );
   nor U7277 ( n7384,n7386,n7387 );
   nor U7278 ( n7387,n5986,n7375 );
   xor U7279 ( n7375,n7388,n7389 );
   nor U7280 ( n7386,n5998,n7390 );
   nor U7281 ( n7390,n7391,n7392 );
   nor U7282 ( n7392,n7388,n7393 );
   nand U7283 ( n7393,n7394,n7395 );
   nand U7284 ( n7394,n7349,n7396 );
   nor U7285 ( n7391,n7397,n7398 );
   nand U7286 ( n7398,n7399,n7396 );
   nand U7287 ( n7399,n7395,n7345 );
   not U7288 ( n7345,n7349 );
   nor U7289 ( n7349,n7400,n7315 );
   nand U7290 ( n7397,n7401,n7402 );
   nor U7291 ( n7404,n7405,n7406 );
   nand U7292 ( n7406,n7407,n7408 );
   nand U7293 ( n7408,n6480,n5977 );
   nor U7294 ( n6480,n7409,n7410 );
   and U7295 ( n7410,n7411,n7412 );
   nand U7296 ( n7412,n7325,n6499 );
   nand U7297 ( n7407,n6990,n6481 );
   nor U7298 ( n7405,n6482,n6000 );
   nor U7299 ( n7403,n7413,n7414 );
   nand U7300 ( n7414,n7415,n7416 );
   nand U7301 ( n7416,n7009,n7417 );
   nand U7302 ( n7415,n7010,n7411 );
   nand U7303 ( n7413,n7418,n7419 );
   nand U7304 ( n7419,reg2_reg_12_,n6699 );
   nand U7305 ( n7418,n5989,n6484 );
   nand U7306 ( n6484,n7420,n7421 );
   nand U7307 ( n7421,n7016,n6077 );
   nor U7308 ( n7420,n7422,n7423 );
   nor U7309 ( n7423,n5999,n7424 );
   xor U7310 ( n7424,n7425,n7426 );
   nand U7311 ( n7426,n7427,n7428 );
   and U7312 ( n7422,n7019,n6481 );
   xor U7313 ( n6481,n7425,n7429 );
   nor U7314 ( n7431,n7432,n7433 );
   nand U7315 ( n7433,n7434,n7435 );
   nand U7316 ( n7435,n7003,n6466 );
   xor U7317 ( n6466,n7409,n6471 );
   nand U7318 ( n7434,n6990,n6467 );
   not U7319 ( n6467,n7436 );
   nor U7320 ( n7432,n6468,n7004 );
   nor U7321 ( n7430,n7437,n7438 );
   nand U7322 ( n7438,n7439,n7440 );
   nand U7323 ( n7440,n7009,n7441 );
   nand U7324 ( n7439,n7010,n7442 );
   nand U7325 ( n7437,n7443,n7444 );
   nand U7326 ( n7444,reg2_reg_13_,n6002 );
   nand U7327 ( n7443,n5989,n6470 );
   nand U7328 ( n6470,n7445,n7446 );
   nand U7329 ( n7446,n7016,n6074 );
   nor U7330 ( n7445,n7447,n7448 );
   nor U7331 ( n7448,n6718,n7436 );
   nand U7332 ( n7436,n7449,n7450 );
   nand U7333 ( n7450,n7451,n7452 );
   nor U7334 ( n7451,n7453,n7454 );
   nor U7335 ( n7454,n7455,n7429 );
   nand U7336 ( n7449,n7456,n7457 );
   nand U7337 ( n7457,n7458,n7429 );
   nand U7338 ( n7429,n7459,n7460 );
   nand U7339 ( n7459,n7381,n6077 );
   nor U7340 ( n7456,n7455,n7461 );
   nor U7341 ( n7447,n6705,n7462 );
   xor U7342 ( n7462,n7463,n7461 );
   not U7343 ( n7461,n7464 );
   nor U7344 ( n7466,n7467,n7468 );
   nand U7345 ( n7468,n7469,n7470 );
   nand U7346 ( n7470,n6452,n5977 );
   nor U7347 ( n6452,n7471,n7472 );
   and U7348 ( n7472,n7473,n7474 );
   nand U7349 ( n7474,n7409,n6471 );
   nand U7350 ( n7469,n6990,n6453 );
   nor U7351 ( n7467,n6454,n6000 );
   nor U7352 ( n7465,n7475,n7476 );
   nand U7353 ( n7476,n7477,n7478 );
   or U7354 ( n7478,n6683,n7479 );
   nand U7355 ( n7477,n7010,n7473 );
   nand U7356 ( n7475,n7480,n7481 );
   nand U7357 ( n7481,reg2_reg_14_,n6699 );
   nand U7358 ( n7480,n6700,n6456 );
   nand U7359 ( n6456,n7482,n7483 );
   nand U7360 ( n7483,n7016,n6071 );
   nor U7361 ( n7482,n7484,n7485 );
   and U7362 ( n7485,n7019,n6453 );
   xor U7363 ( n6453,n7486,n7487 );
   nor U7364 ( n7486,n7488,n7489 );
   nor U7365 ( n7484,n5998,n7490 );
   nand U7366 ( n7490,n7491,n7492 );
   nand U7367 ( n7492,n7493,n7494 );
   nor U7368 ( n7493,n7495,n7496 );
   or U7369 ( n7491,n7487,n7494 );
   nor U7370 ( n7498,n7499,n7500 );
   nand U7371 ( n7500,n7501,n7502 );
   nand U7372 ( n7502,n7003,n6438 );
   xor U7373 ( n6438,n6443,n7471 );
   nand U7374 ( n7501,n5978,n6439 );
   not U7375 ( n6439,n7503 );
   nor U7376 ( n7499,n6440,n7004 );
   nor U7377 ( n7497,n7504,n7505 );
   nand U7378 ( n7505,n7506,n7507 );
   nand U7379 ( n7507,n7009,n7508 );
   nand U7380 ( n7506,n7010,n7509 );
   nand U7381 ( n7504,n7510,n7511 );
   nand U7382 ( n7511,reg2_reg_15_,n6002 );
   nand U7383 ( n7510,n6700,n6442 );
   nand U7384 ( n6442,n7512,n7513 );
   nor U7385 ( n7513,n7514,n7515 );
   nor U7386 ( n7515,n7516,n7503 );
   xor U7387 ( n7503,n7517,n7518 );
   and U7388 ( n7516,n7519,n7520 );
   nor U7389 ( n7514,n7285,n7521 );
   nor U7390 ( n7285,n7522,n7523 );
   nor U7391 ( n7512,n7524,n7525 );
   nor U7392 ( n7525,n6468,n6729 );
   nor U7393 ( n7524,n7287,n7521 );
   nand U7394 ( n7521,n7526,n7527 );
   nand U7395 ( n7527,n7528,n7529 );
   and U7396 ( n7528,n7530,n7531 );
   nand U7397 ( n7526,n7517,n7532 );
   not U7398 ( n7517,n7533 );
   nor U7399 ( n7535,n7536,n7537 );
   nand U7400 ( n7537,n7538,n7539 );
   nand U7401 ( n7539,n6424,n5977 );
   nor U7402 ( n6424,n7540,n7541 );
   and U7403 ( n7541,n7542,n7543 );
   nand U7404 ( n7543,n7471,n6443 );
   nand U7405 ( n7538,n6990,n6425 );
   not U7406 ( n6425,n7544 );
   nor U7407 ( n7536,n6426,n6000 );
   nor U7408 ( n7534,n7545,n7546 );
   nand U7409 ( n7546,n7547,n7548 );
   nand U7410 ( n7548,n7009,n7549 );
   nand U7411 ( n7547,n5981,n7542 );
   nand U7412 ( n7545,n7550,n7551 );
   nand U7413 ( n7551,reg2_reg_16_,n6002 );
   nand U7414 ( n7550,n6700,n6428 );
   nand U7415 ( n6428,n7552,n7553 );
   nand U7416 ( n7553,n7016,n6065 );
   nor U7417 ( n7552,n7554,n7555 );
   nor U7418 ( n7555,n5998,n7556 );
   nor U7419 ( n7556,n7557,n7558 );
   nor U7420 ( n7558,n7559,n7560 );
   nand U7421 ( n7560,n7561,n7531 );
   nand U7422 ( n7561,n7532,n7530 );
   not U7423 ( n7532,n7529 );
   nor U7424 ( n7557,n7562,n7563 );
   nand U7425 ( n7563,n7564,n7565 );
   nand U7426 ( n7564,n7531,n7529 );
   nand U7427 ( n7529,n7566,n7567 );
   nand U7428 ( n7567,n7494,n7568 );
   nor U7429 ( n7554,n5986,n7544 );
   xor U7430 ( n7544,n7559,n7569 );
   nor U7431 ( n7571,n7572,n7573 );
   nand U7432 ( n7573,n7574,n7575 );
   nand U7433 ( n7575,n7003,n6410 );
   xor U7434 ( n6410,n7540,n6415 );
   nand U7435 ( n7574,n6990,n6411 );
   not U7436 ( n6411,n7576 );
   nor U7437 ( n7572,n6412,n7004 );
   nor U7438 ( n7570,n7577,n7578 );
   nand U7439 ( n7578,n7579,n7580 );
   nand U7440 ( n7580,n7009,n7581 );
   nand U7441 ( n7579,n7010,n7582 );
   nand U7442 ( n7577,n7583,n7584 );
   nand U7443 ( n7584,reg2_reg_17_,n6002 );
   nand U7444 ( n7583,n6700,n6414 );
   nand U7445 ( n6414,n7585,n7586 );
   nand U7446 ( n7586,n7016,n6062 );
   nor U7447 ( n7585,n7587,n7588 );
   nor U7448 ( n7588,n5999,n7589 );
   xor U7449 ( n7589,n7590,n7591 );
   nor U7450 ( n7590,n7592,n7593 );
   not U7451 ( n7593,n7594 );
   nor U7452 ( n7587,n6718,n7576 );
   nand U7453 ( n7576,n7595,n7596 );
   nand U7454 ( n7596,n7597,n7598 );
   nand U7455 ( n7598,n7569,n7599 );
   and U7456 ( n7597,n7600,n7591 );
   nand U7457 ( n7595,n7601,n7602 );
   nor U7458 ( n7601,n7603,n7604 );
   nor U7459 ( n7604,n7605,n7569 );
   nor U7460 ( n7603,n6426,n6415 );
   nor U7461 ( n7607,n7608,n7609 );
   nand U7462 ( n7609,n7610,n7611 );
   nand U7463 ( n7611,n6396,n5977 );
   nor U7464 ( n6396,n7612,n7613 );
   and U7465 ( n7613,n7614,n7615 );
   nand U7466 ( n7615,n7540,n6415 );
   nand U7467 ( n7610,n6990,n6397 );
   not U7468 ( n6397,n7616 );
   nor U7469 ( n7608,n6398,n6000 );
   nor U7470 ( n7606,n7617,n7618 );
   nand U7471 ( n7618,n7619,n7620 );
   or U7472 ( n7620,n6683,n7621 );
   nand U7473 ( n7619,n7010,n7614 );
   nand U7474 ( n7617,n7622,n7623 );
   nand U7475 ( n7623,reg2_reg_18_,n6699 );
   nand U7476 ( n7622,n6700,n6400 );
   nand U7477 ( n6400,n7624,n7625 );
   nand U7478 ( n7625,n7016,n6059 );
   nor U7479 ( n7624,n7626,n7627 );
   nor U7480 ( n7627,n5986,n7616 );
   xor U7481 ( n7616,n7628,n7629 );
   nor U7482 ( n7626,n6705,n7630 );
   xor U7483 ( n7630,n7628,n7631 );
   nor U7484 ( n7633,n7634,n7635 );
   nand U7485 ( n7635,n7636,n7637 );
   nand U7486 ( n7637,n7003,n6382 );
   xor U7487 ( n6382,n6387,n7612 );
   nand U7488 ( n7636,n6990,n6383 );
   nor U7489 ( n7634,n6384,n7004 );
   nor U7490 ( n7632,n7638,n7639 );
   nand U7491 ( n7639,n7640,n7641 );
   nand U7492 ( n7641,n5976,n7642 );
   nand U7493 ( n7640,n7010,n7643 );
   nand U7494 ( n7638,n7644,n7645 );
   nand U7495 ( n7645,reg2_reg_19_,n6699 );
   nand U7496 ( n7644,n6700,n6386 );
   nand U7497 ( n6386,n7646,n7647 );
   nand U7498 ( n7647,n7016,n6056 );
   nor U7499 ( n7646,n7648,n7649 );
   and U7500 ( n7649,n7019,n6383 );
   xor U7501 ( n6383,n7650,n7651 );
   nor U7502 ( n7648,n5999,n7652 );
   xor U7503 ( n7652,n7650,n7653 );
   nor U7504 ( n7655,n7656,n7657 );
   nand U7505 ( n7657,n7658,n7659 );
   nand U7506 ( n7659,n6368,n5977 );
   nor U7507 ( n6368,n7660,n7661 );
   and U7508 ( n7661,n7662,n7663 );
   nand U7509 ( n7663,n7612,n6387 );
   nand U7510 ( n7658,n6990,n6369 );
   not U7511 ( n6369,n7664 );
   nor U7512 ( n7656,n6370,n7004 );
   nor U7513 ( n7654,n7665,n7666 );
   nand U7514 ( n7666,n7667,n7668 );
   nand U7515 ( n7668,n7009,n7669 );
   nand U7516 ( n7667,n7010,n7662 );
   nand U7517 ( n7665,n7670,n7671 );
   nand U7518 ( n7671,reg2_reg_20_,n6002 );
   nand U7519 ( n7670,n6700,n6372 );
   nand U7520 ( n6372,n7672,n7673 );
   nand U7521 ( n7673,n7016,n6053 );
   nor U7522 ( n7672,n7674,n7675 );
   nor U7523 ( n7675,n5998,n7676 );
   xor U7524 ( n7676,n7677,n7678 );
   nand U7525 ( n7678,n7679,n7680 );
   or U7526 ( n7680,n7681,n7682 );
   nor U7527 ( n7674,n5986,n7664 );
   nand U7528 ( n7664,n7683,n7684 );
   nand U7529 ( n7684,n7685,n7686 );
   nor U7530 ( n7685,n7687,n7688 );
   nor U7531 ( n7688,n7651,n7689 );
   nand U7532 ( n7683,n7690,n7691 );
   nand U7533 ( n7691,n7651,n7692 );
   nor U7534 ( n7690,n7689,n7677 );
   not U7535 ( n7677,n7693 );
   nor U7536 ( n7695,n7696,n7697 );
   nand U7537 ( n7697,n7698,n7699 );
   nand U7538 ( n7699,n7003,n6354 );
   xor U7539 ( n6354,n7660,n6359 );
   nand U7540 ( n7698,n5978,n6355 );
   not U7541 ( n6355,n7700 );
   nor U7542 ( n7696,n6356,n6000 );
   nor U7543 ( n7694,n7701,n7702 );
   nand U7544 ( n7702,n7703,n7704 );
   nand U7545 ( n7704,n7009,n7705 );
   nand U7546 ( n7703,n5981,n7706 );
   nand U7547 ( n7701,n7707,n7708 );
   nand U7548 ( n7708,reg2_reg_21_,n6699 );
   nand U7549 ( n7707,n6700,n6358 );
   nand U7550 ( n6358,n7709,n7710 );
   nor U7551 ( n7710,n7711,n7712 );
   nor U7552 ( n7712,n6705,n7713 );
   nand U7553 ( n7713,n7714,n7715 );
   nand U7554 ( n7715,n7716,n7717 );
   and U7555 ( n7716,n7718,n7719 );
   or U7556 ( n7714,n7720,n7717 );
   nor U7557 ( n7711,n7519,n7700 );
   nor U7558 ( n7709,n7721,n7722 );
   nor U7559 ( n7722,n6384,n6729 );
   nor U7560 ( n7721,n7520,n7700 );
   xor U7561 ( n7700,n7723,n7720 );
   nand U7562 ( n7723,n7724,n7725 );
   nand U7563 ( n7725,n7651,n7686 );
   not U7564 ( n7686,n7726 );
   and U7565 ( n7651,n7727,n7728 );
   nand U7566 ( n7728,n7629,n7729 );
   and U7567 ( n7629,n7730,n7731 );
   nor U7568 ( n7733,n7734,n7735 );
   nand U7569 ( n7735,n7736,n7737 );
   nand U7570 ( n7737,n6340,n5977 );
   nor U7571 ( n6340,n7738,n7739 );
   and U7572 ( n7739,n7740,n7741 );
   nand U7573 ( n7741,n7660,n6359 );
   nand U7574 ( n7736,n5978,n6341 );
   nor U7575 ( n7734,n6342,n7004 );
   nor U7576 ( n7732,n7742,n7743 );
   nand U7577 ( n7743,n7744,n7745 );
   or U7578 ( n7745,n6683,n7746 );
   nand U7579 ( n7744,n5981,n7740 );
   nand U7580 ( n7742,n7747,n7748 );
   nand U7581 ( n7748,reg2_reg_22_,n6699 );
   nand U7582 ( n7747,n6700,n6344 );
   nand U7583 ( n6344,n7749,n7750 );
   nor U7584 ( n7750,n7751,n7752 );
   nand U7585 ( n7752,n7753,n7754 );
   nand U7586 ( n7754,n7755,n7756 );
   nand U7587 ( n7756,n7287,n7045 );
   nor U7588 ( n7755,n7757,n7758 );
   nor U7589 ( n7758,n7759,n7760 );
   and U7590 ( n7757,n7761,n7762 );
   nand U7591 ( n7753,n7763,n7764 );
   nor U7592 ( n7751,n7765,n7766 );
   nor U7593 ( n7766,n7767,n7768 );
   nor U7594 ( n7768,n7769,n7759 );
   nor U7595 ( n7767,n7759,n7770 );
   nor U7596 ( n7749,n7771,n7772 );
   nor U7597 ( n7772,n6370,n6729 );
   and U7598 ( n7771,n7019,n6341 );
   xor U7599 ( n6341,n7765,n7773 );
   nand U7600 ( n7773,n7774,n7775 );
   not U7601 ( n7765,n7760 );
   nor U7602 ( n7777,n7778,n7779 );
   nand U7603 ( n7779,n7780,n7781 );
   nand U7604 ( n7781,n5978,n6326 );
   xor U7605 ( n6326,n7782,n7783 );
   nand U7606 ( n7780,n7003,n6327 );
   xor U7607 ( n6327,n6331,n7738 );
   nor U7608 ( n7778,n6328,n6000 );
   nor U7609 ( n7776,n7784,n7785 );
   nand U7610 ( n7785,n7786,n7787 );
   nand U7611 ( n7787,n7009,n7788 );
   nand U7612 ( n7786,n7010,n7789 );
   nand U7613 ( n7784,n7790,n7791 );
   nand U7614 ( n7791,reg2_reg_23_,n6002 );
   nand U7615 ( n7790,n6700,n6330 );
   nand U7616 ( n6330,n7792,n7793 );
   nor U7617 ( n7793,n7794,n7795 );
   nor U7618 ( n7795,n7796,n7797 );
   nand U7619 ( n7797,n7019,n7798 );
   not U7620 ( n7796,n7782 );
   nor U7621 ( n7794,n7799,n7782 );
   nor U7622 ( n7799,n7800,n7801 );
   nand U7623 ( n7801,n7802,n7803 );
   nand U7624 ( n7803,n7764,n7804 );
   nand U7625 ( n7764,n7805,n7806 );
   nand U7626 ( n7806,n7807,n7759 );
   nand U7627 ( n7805,n7523,n7759 );
   nand U7628 ( n7802,n7808,n7019 );
   nand U7629 ( n7800,n7809,n7810 );
   nand U7630 ( n7810,n7811,n7812 );
   nand U7631 ( n7812,n7813,n7770 );
   nand U7632 ( n7809,n7814,n7762 );
   nand U7633 ( n7762,n7815,n7816 );
   nand U7634 ( n7816,n7817,n7717 );
   nand U7635 ( n7815,n7818,n7804 );
   nor U7636 ( n7792,n7819,n7820 );
   nor U7637 ( n7820,n6356,n6729 );
   nor U7638 ( n7819,n7821,n7822 );
   nand U7639 ( n7822,n7823,n7824 );
   nand U7640 ( n7823,n7825,n7826 );
   or U7641 ( n7826,n7770,n7759 );
   nor U7642 ( n7825,n7827,n7828 );
   nor U7643 ( n7828,n5998,n7804 );
   nor U7644 ( n7827,n7813,n7759 );
   nand U7645 ( n7759,n7719,n7829 );
   nand U7646 ( n7829,n7717,n7718 );
   nand U7647 ( n7717,n7830,n7831 );
   nand U7648 ( n7831,n7832,n7653 );
   not U7649 ( n7830,n7833 );
   nor U7650 ( n7813,n7834,n7835 );
   nor U7651 ( n7837,n7838,n7839 );
   nand U7652 ( n7839,n7840,n7841 );
   nand U7653 ( n7841,n6312,n5977 );
   nor U7654 ( n6312,n7842,n7843 );
   and U7655 ( n7843,n7844,n7845 );
   nand U7656 ( n7845,n7738,n6331 );
   nand U7657 ( n7840,n5978,n6313 );
   xor U7658 ( n6313,n7846,n7847 );
   nor U7659 ( n7838,n6314,n7004 );
   nor U7660 ( n7836,n7848,n7849 );
   nand U7661 ( n7849,n7850,n7851 );
   nand U7662 ( n7851,n7009,n7852 );
   nand U7663 ( n7850,n5981,n7844 );
   nand U7664 ( n7848,n7853,n7854 );
   nand U7665 ( n7854,reg2_reg_24_,n6699 );
   nand U7666 ( n7853,n6700,n6316 );
   nand U7667 ( n6316,n7855,n7856 );
   nand U7668 ( n7856,n5992,n6041 );
   nor U7669 ( n7855,n7857,n7858 );
   nor U7670 ( n7858,n5999,n7859 );
   xor U7671 ( n7859,n7860,n7861 );
   nand U7672 ( n7861,n7862,n7863 );
   nor U7673 ( n7857,n5986,n7864 );
   xor U7674 ( n7864,n7846,n7865 );
   nor U7675 ( n7867,n7868,n7869 );
   nand U7676 ( n7869,n7870,n7871 );
   nand U7677 ( n7871,n5978,n6298 );
   xor U7678 ( n6298,n7872,n7873 );
   nand U7679 ( n7870,n7003,n6299 );
   xor U7680 ( n6299,n7842,n6303 );
   nor U7681 ( n7868,n6300,n6000 );
   nor U7682 ( n7866,n7874,n7875 );
   nand U7683 ( n7875,n7876,n7877 );
   or U7684 ( n7877,n6683,n7878 );
   not U7685 ( n6683,n7009 );
   nand U7686 ( n7876,n5981,n7879 );
   nand U7687 ( n7874,n7880,n7881 );
   nand U7688 ( n7881,reg2_reg_25_,n6002 );
   nand U7689 ( n7880,n6700,n6302 );
   nand U7690 ( n6302,n7882,n7883 );
   nand U7691 ( n7883,n7016,n6038 );
   nor U7692 ( n7882,n7884,n7885 );
   nor U7693 ( n7885,n7886,n7887 );
   nor U7694 ( n7886,n7888,n7889 );
   nor U7695 ( n7889,n5986,n7890 );
   nor U7696 ( n7888,n5999,n7891 );
   nor U7697 ( n7884,n7873,n7892 );
   nor U7698 ( n7892,n7893,n7894 );
   nor U7699 ( n7894,n6718,n7895 );
   nor U7700 ( n7893,n7896,n5998 );
   not U7701 ( n7873,n7887 );
   nor U7702 ( n7898,n7899,n7900 );
   nand U7703 ( n7900,n7901,n7902 );
   nand U7704 ( n7902,n6284,n7003 );
   nor U7705 ( n6284,n7903,n7904 );
   and U7706 ( n7904,n7905,n7906 );
   nand U7707 ( n7906,n7842,n6303 );
   nand U7708 ( n7901,n5978,n6285 );
   and U7709 ( n6285,n7907,n7908 );
   nand U7710 ( n7908,n7909,n7910 );
   nand U7711 ( n7910,n7911,n7872 );
   not U7712 ( n7872,n7912 );
   nand U7713 ( n7907,n7913,n7914 );
   nand U7714 ( n7914,n7912,n7915 );
   nor U7715 ( n7912,n7916,n7917 );
   not U7716 ( n7913,n7918 );
   nor U7717 ( n7899,n6286,n7004 );
   nor U7718 ( n7897,n7919,n7920 );
   nand U7719 ( n7920,n7921,n7922 );
   nand U7720 ( n7922,n7009,n7923 );
   nand U7721 ( n7921,n5981,n7905 );
   nand U7722 ( n7919,n7924,n7925 );
   nand U7723 ( n7925,reg2_reg_26_,n6002 );
   nand U7724 ( n7924,n6700,n6288 );
   nand U7725 ( n6288,n7926,n7927 );
   nor U7726 ( n7927,n7928,n7929 );
   nor U7727 ( n7929,n7236,n7930 );
   nand U7728 ( n7930,n7931,n7932 );
   nand U7729 ( n7931,n7933,n7934 );
   nor U7730 ( n7928,n7935,n7936 );
   nand U7731 ( n7936,n7019,n7937 );
   nand U7732 ( n7937,n7909,n7938 );
   nand U7733 ( n7938,n7890,n7911 );
   nor U7734 ( n7909,n7939,n7940 );
   nor U7735 ( n7935,n7941,n7918 );
   nand U7736 ( n7918,n7942,n7943 );
   nor U7737 ( n7941,n7939,n7890 );
   not U7738 ( n7890,n7895 );
   nand U7739 ( n7895,n7944,n7945 );
   nand U7740 ( n7945,n7946,n7947 );
   not U7741 ( n7944,n7948 );
   nor U7742 ( n7926,n7949,n7950 );
   nor U7743 ( n7950,n6314,n6729 );
   nor U7744 ( n7949,n7045,n7951 );
   nand U7745 ( n7951,n7952,n7932 );
   nand U7746 ( n7932,n7940,n7953 );
   not U7747 ( n7940,n7954 );
   nand U7748 ( n7952,n7955,n7956 );
   not U7749 ( n7956,n7953 );
   nor U7750 ( n7955,n7957,n7958 );
   nor U7751 ( n7960,n7961,n7962 );
   nand U7752 ( n7962,n7963,n7964 );
   nand U7753 ( n7964,n5978,n6270 );
   xor U7754 ( n6270,n7965,n7966 );
   nand U7755 ( n7963,n7003,n6271 );
   xor U7756 ( n6271,n6275,n7903 );
   nor U7757 ( n7961,n6272,n6000 );
   nor U7758 ( n7959,n7967,n7968 );
   nand U7759 ( n7968,n7969,n7970 );
   nand U7760 ( n7970,n5976,n7971 );
   nand U7761 ( n7969,n5981,n7972 );
   nand U7762 ( n7967,n7973,n7974 );
   nand U7763 ( n7974,reg2_reg_27_,n6699 );
   nand U7764 ( n7973,n6700,n6274 );
   nand U7765 ( n6274,n7975,n7976 );
   nor U7766 ( n7976,n7977,n7978 );
   nor U7767 ( n7978,n7965,n7979 );
   nor U7768 ( n7979,n7980,n7981 );
   nor U7769 ( n7981,n6718,n7982 );
   nor U7770 ( n7980,n7983,n7984 );
   nand U7771 ( n7984,n7985,n7934 );
   nor U7772 ( n7977,n7986,n7987 );
   nor U7773 ( n7986,n7988,n7989 );
   nand U7774 ( n7989,n7990,n7991 );
   nand U7775 ( n7991,n7982,n7019 );
   and U7776 ( n7982,n7992,n7993 );
   or U7777 ( n7990,n7985,n7983 );
   nor U7778 ( n7983,n7807,n7058 );
   nor U7779 ( n7988,n7236,n7934 );
   nor U7780 ( n7236,n7807,n7834 );
   nor U7781 ( n7975,n7994,n7995 );
   nor U7782 ( n7995,n6300,n6729 );
   not U7783 ( n6729,n7016 );
   nor U7784 ( n7994,n7996,n7997 );
   nor U7785 ( n7997,n7998,n7999 );
   nor U7786 ( n7999,n8000,n7769 );
   nor U7787 ( n8000,n8001,n7933 );
   nor U7788 ( n8001,n7965,n7957 );
   nor U7789 ( n7998,n8002,n7045 );
   nor U7790 ( n8002,n7933,n8003 );
   xor U7791 ( n8003,n7987,n7957 );
   nor U7792 ( n7996,n7965,n7985 );
   not U7793 ( n7985,n7933 );
   nor U7794 ( n8005,n8006,n8007 );
   nand U7795 ( n8007,n8008,n8009 );
   nand U7796 ( n8009,n6253,n5977 );
   nor U7797 ( n6253,n6693,n8010 );
   and U7798 ( n8010,n8011,n8012 );
   nand U7799 ( n8012,n7903,n6275 );
   nand U7800 ( n8008,n6990,n6256 );
   xor U7801 ( n6256,n6691,n8013 );
   and U7802 ( n6691,n8014,n8015 );
   or U7803 ( n8015,n7966,n8016 );
   nand U7804 ( n7966,n7992,n8017 );
   nand U7805 ( n8017,n7916,n7942 );
   not U7806 ( n7942,n8018 );
   nor U7807 ( n7916,n7847,n7948 );
   nand U7808 ( n7847,n8019,n8020 );
   nand U7809 ( n8020,n8021,n7783 );
   nand U7810 ( n7783,n8022,n8023 );
   nand U7811 ( n8023,n8024,n7774 );
   and U7812 ( n8024,n7775,n8025 );
   nor U7813 ( n7992,n8026,n8027 );
   not U7814 ( n8027,n8028 );
   nor U7815 ( n6990,n8029,n6002 );
   nor U7816 ( n8006,n6257,n6000 );
   not U7817 ( n7004,n6989 );
   nor U7818 ( n6989,n6699,n5944 );
   nor U7819 ( n8004,n8030,n8031 );
   nand U7820 ( n8031,n8032,n8033 );
   nand U7821 ( n8033,n5976,n8034 );
   nor U7822 ( n7009,n6002,n8035 );
   nand U7823 ( n8032,n5981,n8011 );
   nand U7824 ( n8030,n8036,n8037 );
   nand U7825 ( n8037,reg2_reg_28_,n6002 );
   nand U7826 ( n8036,n6700,n6260 );
   nand U7827 ( n6260,n8038,n8039 );
   nand U7828 ( n8039,n7016,n6029 );
   nor U7829 ( n7016,n8040,n8041 );
   nor U7830 ( n8038,n8042,n8043 );
   nor U7831 ( n8043,n8044,n8045 );
   nor U7832 ( n8044,n8046,n8047 );
   nor U7833 ( n8047,n5998,n6714 );
   not U7834 ( n6714,n6717 );
   nor U7835 ( n8046,n5986,n8048 );
   nor U7836 ( n8042,n8013,n8049 );
   nor U7837 ( n8049,n8050,n8051 );
   nor U7838 ( n8051,n6717,n6705 );
   nor U7839 ( n6705,n7834,n7522 );
   nand U7840 ( n7522,n7770,n7045 );
   nand U7841 ( n7834,n7769,n7287 );
   nor U7842 ( n6717,n8052,n8053 );
   and U7843 ( n8052,n8054,n8055 );
   nor U7844 ( n8054,n7957,n7933 );
   nor U7845 ( n7933,n7953,n7958 );
   nand U7846 ( n7953,n8056,n8057 );
   or U7847 ( n8056,n8058,n7896 );
   not U7848 ( n7896,n7891 );
   nand U7849 ( n7891,n8059,n8060 );
   nand U7850 ( n8059,n8061,n7863 );
   nand U7851 ( n7863,n8062,n8063 );
   nor U7852 ( n8063,n8064,n8065 );
   and U7853 ( n8062,n7653,n7832 );
   not U7854 ( n7653,n7681 );
   nand U7855 ( n7681,n8066,n8067 );
   nand U7856 ( n8067,n6412,n8068 );
   nand U7857 ( n8068,n6401,n7631 );
   or U7858 ( n8066,n7631,n6401 );
   nand U7859 ( n7631,n8069,n8070 );
   nand U7860 ( n8070,n8071,n8072 );
   nand U7861 ( n8072,n8073,n7594 );
   nand U7862 ( n7594,n8074,n7565 );
   nand U7863 ( n8074,n8075,n8076 );
   nand U7864 ( n8076,n8077,n7495 );
   not U7865 ( n8075,n7562 );
   nand U7866 ( n7562,n7530,n8078 );
   nand U7867 ( n8069,n7592,n8071 );
   not U7868 ( n8071,n8079 );
   and U7869 ( n7592,n8080,n8077 );
   not U7870 ( n8077,n8081 );
   and U7871 ( n8080,n7568,n7494 );
   nand U7872 ( n7494,n8082,n8083 );
   nand U7873 ( n8083,n7463,n8084 );
   nor U7874 ( n7463,n8085,n8086 );
   and U7875 ( n8085,n8087,n8088 );
   and U7876 ( n8087,n7427,n7428 );
   nand U7877 ( n7428,n8089,n7400 );
   nor U7878 ( n7400,n7317,n7314 );
   not U7879 ( n7317,n7313 );
   nand U7880 ( n7313,n8090,n8091 );
   nor U7881 ( n8091,n8092,n8093 );
   nor U7882 ( n8093,n7280,n8094 );
   nand U7883 ( n8094,n7279,n8095 );
   nand U7884 ( n7280,n8096,n8097 );
   nand U7885 ( n8096,n7092,n8098 );
   nor U7886 ( n8092,n8099,n8100 );
   nand U7887 ( n8100,n8101,n7194 );
   or U7888 ( n8101,n7191,n8102 );
   or U7889 ( n7191,n7154,n8103 );
   not U7890 ( n8099,n8095 );
   nor U7891 ( n8090,n8104,n8105 );
   nor U7892 ( n8105,n6552,n7256 );
   nor U7893 ( n8104,n8106,n7275 );
   not U7894 ( n7275,n7228 );
   and U7895 ( n8089,n7401,n7395 );
   nand U7896 ( n7427,n8107,n7401 );
   nand U7897 ( n8107,n8108,n8109 );
   nand U7898 ( n8109,n7315,n7395 );
   and U7899 ( n8108,n7402,n7396 );
   not U7900 ( n7396,n7346 );
   and U7901 ( n8061,n7862,n8110 );
   nand U7902 ( n7862,n8111,n7824 );
   not U7903 ( n7824,n8064 );
   nand U7904 ( n8111,n8112,n8113 );
   nand U7905 ( n8113,n7817,n7833 );
   nand U7906 ( n7833,n8114,n8115 );
   nand U7907 ( n8115,n8116,n8117 );
   nor U7908 ( n8050,n6723,n5986 );
   not U7909 ( n6718,n7019 );
   nand U7910 ( n7019,n7520,n7519 );
   nor U7911 ( n7520,n8118,n8119 );
   not U7912 ( n8119,n8120 );
   not U7913 ( n6723,n8048 );
   nand U7914 ( n8048,n8121,n8122 );
   nor U7915 ( n8122,n8123,n8016 );
   and U7916 ( n8123,n8014,n8026 );
   nor U7917 ( n8026,n8018,n7947 );
   not U7918 ( n7947,n7917 );
   not U7919 ( n8014,n8124 );
   nor U7920 ( n8121,n8125,n8126 );
   nor U7921 ( n8126,n8124,n7993 );
   nand U7922 ( n7993,n8127,n7865 );
   not U7923 ( n7865,n7946 );
   nand U7924 ( n7946,n8019,n8128 );
   nand U7925 ( n8128,n7808,n8021 );
   not U7926 ( n7808,n7798 );
   nand U7927 ( n7798,n8129,n8130 );
   nand U7928 ( n8130,n8022,n8131 );
   nand U7929 ( n8131,n8025,n7775 );
   nand U7930 ( n7775,n8132,n8133 );
   nand U7931 ( n8132,n8134,n7724 );
   and U7932 ( n7724,n8135,n8136 );
   nand U7933 ( n8136,n7689,n8137 );
   nor U7934 ( n8134,n8138,n8139 );
   nor U7935 ( n8139,n6370,n6359 );
   nor U7936 ( n8138,n8140,n7726 );
   nor U7937 ( n8140,n8141,n8142 );
   nor U7938 ( n8142,n6401,n7731 );
   nor U7939 ( n8141,n6412,n8143 );
   and U7940 ( n8143,n7731,n6401 );
   nand U7941 ( n7731,n8144,n8145 );
   nand U7942 ( n8145,n8146,n7600 );
   nand U7943 ( n8129,n8147,n8022 );
   not U7944 ( n8147,n7774 );
   nand U7945 ( n7774,n8148,n8149 );
   and U7946 ( n8149,n7727,n8133 );
   nor U7947 ( n8148,n7726,n7730 );
   nand U7948 ( n7730,n7602,n7569 );
   nand U7949 ( n7569,n8150,n8151 );
   nand U7950 ( n8151,n8152,n6065 );
   nand U7951 ( n8152,n6443,n7518 );
   or U7952 ( n8150,n7518,n6443 );
   nand U7953 ( n7518,n8153,n8154 );
   nand U7954 ( n8153,n8155,n8156 );
   not U7955 ( n8156,n7489 );
   nand U7956 ( n7489,n8157,n8158 );
   nand U7957 ( n8158,n8159,n8160 );
   nand U7958 ( n8159,n8161,n8162 );
   nand U7959 ( n8162,n8163,n7452 );
   not U7960 ( n7452,n8164 );
   nor U7961 ( n8163,n6510,n6499 );
   nor U7962 ( n8155,n7488,n8165 );
   nor U7963 ( n8165,n6468,n6457 );
   nor U7964 ( n7488,n8164,n7460 );
   nand U7965 ( n7460,n7389,n8166 );
   nand U7966 ( n8166,n6510,n6499 );
   nand U7967 ( n7389,n8167,n8168 );
   nand U7968 ( n8168,n7355,n8169 );
   nor U7969 ( n8167,n7359,n8170 );
   nor U7970 ( n8170,n8171,n7358 );
   nand U7971 ( n7358,n8169,n7354 );
   nor U7972 ( n8171,n8172,n7368 );
   nor U7973 ( n8172,n7364,n8173 );
   nor U7974 ( n8173,n8174,n8175 );
   not U7975 ( n8175,n7365 );
   nand U7976 ( n7365,n7367,n8176 );
   nand U7977 ( n8176,n8177,n8178 );
   not U7978 ( n8178,n7242 );
   and U7979 ( n8174,n7367,n7243 );
   and U7980 ( n7243,n8179,n7203 );
   nand U7981 ( n7203,n8180,n8181 );
   nand U7982 ( n8181,n7164,n7128 );
   nand U7983 ( n7128,n8182,n8183 );
   nand U7984 ( n8183,n7097,n8184 );
   nand U7985 ( n7097,n8185,n8186 );
   nand U7986 ( n8186,n7064,n8187 );
   nand U7987 ( n7064,n8188,n8189 );
   nand U7988 ( n8188,n8190,n8191 );
   and U7989 ( n7164,n7160,n8192 );
   nand U7990 ( n8192,n6594,n6583 );
   nor U7991 ( n8180,n7165,n8193 );
   nor U7992 ( n8193,n8194,n8195 );
   not U7993 ( n8179,n7246 );
   nand U7994 ( n8164,n8160,n7458 );
   and U7995 ( n7602,n7599,n8144 );
   nand U7996 ( n7726,n7692,n8137 );
   nor U7997 ( n8127,n7948,n8018 );
   nand U7998 ( n8018,n8196,n7911 );
   nor U7999 ( n8125,n8124,n8028 );
   nand U8000 ( n8028,n8196,n8197 );
   nand U8001 ( n8197,n7943,n7915 );
   nor U8002 ( n8199,n8200,n8201 );
   nor U8003 ( n8201,n6231,n6692 );
   nand U8004 ( n6231,n8202,n8203 );
   nand U8005 ( n8203,n6229,n8204 );
   nor U8006 ( n8198,n8205,n8206 );
   and U8007 ( n8206,n6002,reg2_reg_30_ );
   nor U8008 ( n8205,n8207,n6730 );
   nor U8009 ( n8209,n8200,n8210 );
   nor U8010 ( n8210,n6222,n6692 );
   not U8011 ( n6692,n7003 );
   nor U8012 ( n7003,n8211,n6699 );
   xor U8013 ( n6222,n8202,n8212 );
   or U8014 ( n8202,n8204,n6229 );
   nand U8015 ( n8204,n6693,n6244 );
   and U8016 ( n6693,n8213,n7903 );
   and U8017 ( n7903,n8214,n7842 );
   and U8018 ( n7842,n8215,n7738 );
   and U8019 ( n7738,n8216,n7660 );
   and U8020 ( n7660,n8217,n7612 );
   and U8021 ( n7612,n8218,n7540 );
   and U8022 ( n7540,n8219,n7471 );
   and U8023 ( n7471,n8220,n7409 );
   and U8024 ( n7409,n8221,n7325 );
   and U8025 ( n7325,n8222,n7254 );
   and U8026 ( n7254,n8223,n7173 );
   and U8027 ( n7173,n8224,n7104 );
   and U8028 ( n7104,n8225,n7030 );
   and U8029 ( n7030,n8226,n6639 );
   nor U8030 ( n8226,n7032,n6987 );
   nor U8031 ( n8225,n7106,n7079 );
   nor U8032 ( n8224,n7141,n7175 );
   nor U8033 ( n8223,n7216,n7256 );
   nor U8034 ( n8222,n7327,n7302 );
   nor U8035 ( n8221,n7411,n7381 );
   nor U8036 ( n8220,n7442,n7473 );
   nor U8037 ( n8219,n7542,n7509 );
   nor U8038 ( n8218,n7582,n7614 );
   nor U8039 ( n8217,n7662,n7643 );
   nor U8040 ( n8216,n7706,n7740 );
   nor U8041 ( n8215,n7844,n7789 );
   nor U8042 ( n8214,n7905,n7879 );
   nor U8043 ( n8213,n7972,n8011 );
   and U8044 ( n8200,n6220,n5989 );
   not U8045 ( n6700,n6002 );
   nor U8046 ( n6220,n6728,n8227 );
   and U8047 ( n6728,n8228,n8229 );
   or U8048 ( n8229,n5943,b_reg );
   nand U8049 ( n6258,n6666,n8040 );
   nand U8050 ( n8228,n5966,n6666 );
   nor U8051 ( n8208,n8230,n8231 );
   and U8052 ( n8231,n6699,reg2_reg_31_ );
   nor U8053 ( n8230,n8212,n6730 );
   not U8054 ( n6730,n7010 );
   nor U8055 ( n7010,n6699,n6013 );
   not U8056 ( n6243,n6218 );
   nand U8057 ( n6699,n6210,n8232 );
   nand U8058 ( n8232,n8035,n8233 );
   nand U8059 ( n8233,n8234,n8235 );
   nor U8060 ( n8235,n6655,n8236 );
   not U8061 ( n6655,n6212 );
   nor U8062 ( n8234,n6658,n8237 );
   nor U8063 ( n8239,n8240,n8241 );
   nand U8064 ( n8241,n8242,n8243 );
   nand U8065 ( n8243,n8244,n5450 );
   xor U8066 ( n8244,n8246,n8247 );
   xor U8067 ( n8246,reg2_reg_19_,n8248 );
   nand U8068 ( n8248,n8249,n8250 );
   nand U8069 ( n8250,n8251,n8252 );
   or U8070 ( n8251,n8253,n8254 );
   nand U8071 ( n8249,n8254,n8253 );
   nand U8072 ( n8242,n8255,n6001 );
   xor U8073 ( n8255,n6653,n8257 );
   xor U8074 ( n8257,n8258,n8259 );
   nand U8075 ( n8258,n8260,n8261 );
   nand U8076 ( n8261,n8262,n8263 );
   or U8077 ( n8262,n8264,n8253 );
   nand U8078 ( n8260,n8264,n8253 );
   nor U8079 ( n8240,n8247,n8265 );
   nor U8080 ( n8238,n8266,n8267 );
   and U8081 ( n8266,addr_reg_19_,n8268 );
   nand U8082 ( n8270,n8271,n8272 );
   nand U8083 ( n8272,addr_reg_18_,n8268 );
   nand U8084 ( n8271,reg3_reg_18_,n5975 );
   nand U8085 ( n8269,n8273,n8274 );
   nand U8086 ( n8274,n8275,n8276 );
   nand U8087 ( n8276,n8277,n8278 );
   nand U8088 ( n8278,n8279,n8256 );
   xor U8089 ( n8279,n8264,reg1_reg_18_ );
   nor U8090 ( n8277,n8280,n8281 );
   nor U8091 ( n8281,n8282,n8283 );
   not U8092 ( n8275,n8253 );
   nand U8093 ( n8273,n8284,n8253 );
   nand U8094 ( n8284,n8285,n8286 );
   nand U8095 ( n8286,n8245,n8283 );
   xor U8096 ( n8283,n8254,n8252 );
   nand U8097 ( n8254,n8287,n8288 );
   nand U8098 ( n8288,n8289,n8290 );
   or U8099 ( n8289,n8291,n8292 );
   nand U8100 ( n8287,n8292,n8291 );
   nand U8101 ( n8285,n6001,n8293 );
   xor U8102 ( n8293,n8263,n8264 );
   nand U8103 ( n8264,n8294,n8295 );
   nand U8104 ( n8295,n8296,n8297 );
   or U8105 ( n8296,n8298,n8292 );
   nand U8106 ( n8294,n8292,n8298 );
   nand U8107 ( n8300,n8301,n8302 );
   nand U8108 ( n8302,addr_reg_17_,n8268 );
   nand U8109 ( n8301,reg3_reg_17_,n5973 );
   nand U8110 ( n8299,n8303,n8304 );
   nand U8111 ( n8304,n8292,n8305 );
   nand U8112 ( n8305,n8306,n8307 );
   nand U8113 ( n8307,n8245,n8308 );
   nand U8114 ( n8306,n6001,n8309 );
   xor U8115 ( n8309,n8298,n8297 );
   nand U8116 ( n8303,n8310,n8311 );
   nand U8117 ( n8311,n8312,n8313 );
   nand U8118 ( n8313,n8314,n6001 );
   xor U8119 ( n8314,reg1_reg_17_,n8298 );
   nand U8120 ( n8298,n8315,n8316 );
   nand U8121 ( n8316,n8317,n8318 );
   nand U8122 ( n8317,n8319,n8320 );
   or U8123 ( n8315,n8320,n8319 );
   nor U8124 ( n8312,n8280,n8321 );
   nor U8125 ( n8321,n8282,n8308 );
   xor U8126 ( n8308,n8291,n8290 );
   nand U8127 ( n8291,n8322,n8323 );
   nand U8128 ( n8323,n8324,n8325 );
   or U8129 ( n8324,n8326,n8327 );
   nand U8130 ( n8322,n8327,n8326 );
   not U8131 ( n8310,n8292 );
   nand U8132 ( n8329,n8330,n8331 );
   nand U8133 ( n8331,addr_reg_16_,n8268 );
   nand U8134 ( n8330,reg3_reg_16_,n5975 );
   nand U8135 ( n8328,n8332,n8333 );
   nand U8136 ( n8333,n8319,n8334 );
   nand U8137 ( n8334,n8335,n8336 );
   nand U8138 ( n8336,n8256,n8337 );
   xor U8139 ( n8337,n8320,n8318 );
   nor U8140 ( n8335,n8280,n8338 );
   nor U8141 ( n8338,n8282,n8339 );
   not U8142 ( n8319,n8326 );
   nand U8143 ( n8332,n8340,n8326 );
   nand U8144 ( n8340,n8341,n8342 );
   nand U8145 ( n8342,n8245,n8339 );
   xor U8146 ( n8339,n8327,n8325 );
   nand U8147 ( n8327,n8343,n8344 );
   nand U8148 ( n8344,n8345,n8346 );
   or U8149 ( n8345,n8347,n8348 );
   nand U8150 ( n8343,n8348,n8347 );
   nand U8151 ( n8341,n8349,n6001 );
   xor U8152 ( n8349,reg1_reg_16_,n8320 );
   nand U8153 ( n8320,n8350,n8351 );
   nand U8154 ( n8351,reg1_reg_15_,n8352 );
   or U8155 ( n8352,n8353,n8354 );
   nand U8156 ( n8350,n8354,n8353 );
   nand U8157 ( n8356,n8357,n8358 );
   nand U8158 ( n8358,addr_reg_15_,n8268 );
   nand U8159 ( n8357,reg3_reg_15_,n5973 );
   nand U8160 ( n8355,n8359,n8360 );
   nand U8161 ( n8360,n8348,n8361 );
   nand U8162 ( n8361,n8362,n8363 );
   nand U8163 ( n8363,n8245,n8364 );
   nand U8164 ( n8362,n8365,n8256 );
   xor U8165 ( n8365,reg1_reg_15_,n8353 );
   nand U8166 ( n8359,n8354,n8366 );
   nand U8167 ( n8366,n8367,n8368 );
   nand U8168 ( n8368,n8256,n8369 );
   xor U8169 ( n8369,n8353,n8370 );
   nand U8170 ( n8353,n8371,n8372 );
   nand U8171 ( n8372,reg1_reg_14_,n8373 );
   or U8172 ( n8373,n8374,n8375 );
   nand U8173 ( n8371,n8375,n8374 );
   nor U8174 ( n8367,n8280,n8376 );
   nor U8175 ( n8376,n8282,n8364 );
   xor U8176 ( n8364,n8347,n8346 );
   nand U8177 ( n8347,n8377,n8378 );
   nand U8178 ( n8378,n8379,n8380 );
   or U8179 ( n8379,n8381,n8382 );
   nand U8180 ( n8377,n8382,n8381 );
   not U8181 ( n8354,n8348 );
   nand U8182 ( n8384,n8385,n8386 );
   nand U8183 ( n8386,addr_reg_14_,n8268 );
   nand U8184 ( n8385,reg3_reg_14_,n5932 );
   nand U8185 ( n8383,n8387,n8388 );
   nand U8186 ( n8388,n8375,n8389 );
   nand U8187 ( n8389,n8390,n8391 );
   nand U8188 ( n8391,n8256,n8392 );
   xor U8189 ( n8392,n8374,n8393 );
   nor U8190 ( n8390,n8280,n8394 );
   nor U8191 ( n8394,n5980,n8395 );
   not U8192 ( n8375,n8381 );
   nand U8193 ( n8387,n8396,n8381 );
   nand U8194 ( n8396,n8397,n8398 );
   nand U8195 ( n8398,n8245,n8395 );
   xor U8196 ( n8395,n8382,n8380 );
   nand U8197 ( n8382,n8399,n8400 );
   nand U8198 ( n8400,n8401,n8402 );
   or U8199 ( n8401,n8403,n8404 );
   nand U8200 ( n8399,n8404,n8403 );
   nand U8201 ( n8397,n8405,n8256 );
   xor U8202 ( n8405,reg1_reg_14_,n8374 );
   nand U8203 ( n8374,n8406,n8407 );
   nand U8204 ( n8407,reg1_reg_13_,n8408 );
   or U8205 ( n8408,n8409,n8410 );
   nand U8206 ( n8406,n8410,n8409 );
   nand U8207 ( n8412,n8413,n8414 );
   nand U8208 ( n8414,addr_reg_13_,n5449 );
   nand U8209 ( n8413,reg3_reg_13_,n5932 );
   nand U8210 ( n8411,n8415,n8416 );
   nand U8211 ( n8416,n8404,n8417 );
   nand U8212 ( n8417,n8418,n8419 );
   nand U8213 ( n8419,n8245,n8420 );
   nand U8214 ( n8418,n8421,n8256 );
   xor U8215 ( n8421,reg1_reg_13_,n8409 );
   nand U8216 ( n8415,n8410,n8422 );
   nand U8217 ( n8422,n8423,n8424 );
   nand U8218 ( n8424,n6001,n8425 );
   xor U8219 ( n8425,n8409,n8426 );
   nand U8220 ( n8409,n8427,n8428 );
   nand U8221 ( n8428,reg1_reg_12_,n8429 );
   nand U8222 ( n8429,n8430,n8431 );
   or U8223 ( n8427,n8431,n8430 );
   nor U8224 ( n8423,n8280,n8432 );
   nor U8225 ( n8432,n8282,n8420 );
   xor U8226 ( n8420,n8403,n8402 );
   nand U8227 ( n8403,n8433,n8434 );
   nand U8228 ( n8434,n8435,n8436 );
   or U8229 ( n8435,n8430,n8437 );
   nand U8230 ( n8433,n8437,n8430 );
   not U8231 ( n8410,n8404 );
   nand U8232 ( n8439,n8440,n8441 );
   nand U8233 ( n8441,addr_reg_12_,n8268 );
   nand U8234 ( n8440,reg3_reg_12_,n5932 );
   nand U8235 ( n8438,n8442,n8443 );
   nand U8236 ( n8443,n8444,n8445 );
   nand U8237 ( n8445,n8446,n8447 );
   nand U8238 ( n8447,n8448,n6001 );
   xor U8239 ( n8448,reg1_reg_12_,n8431 );
   nor U8240 ( n8446,n8280,n8449 );
   nor U8241 ( n8449,n5980,n8450 );
   not U8242 ( n8444,n8430 );
   nand U8243 ( n8442,n8451,n8430 );
   nand U8244 ( n8451,n8452,n8453 );
   nand U8245 ( n8453,n8245,n8450 );
   xor U8246 ( n8450,n8437,n8436 );
   nand U8247 ( n8437,n8454,n8455 );
   nand U8248 ( n8455,n8456,n8457 );
   or U8249 ( n8456,n8458,n8459 );
   nand U8250 ( n8454,n8459,n8458 );
   nand U8251 ( n8452,n8256,n8460 );
   xor U8252 ( n8460,n8431,n8461 );
   nand U8253 ( n8431,n8462,n8463 );
   nand U8254 ( n8463,n8464,n8465 );
   nand U8255 ( n8464,n8466,n8467 );
   or U8256 ( n8462,n8467,n8466 );
   nand U8257 ( n8469,n8470,n8471 );
   nand U8258 ( n8471,addr_reg_11_,n8268 );
   nand U8259 ( n8470,reg3_reg_11_,n5973 );
   nand U8260 ( n8468,n8472,n8473 );
   nand U8261 ( n8473,n8459,n8474 );
   nand U8262 ( n8474,n8475,n8476 );
   nand U8263 ( n8476,n5450,n8477 );
   nand U8264 ( n8475,n8478,n8256 );
   xor U8265 ( n8478,reg1_reg_11_,n8467 );
   nand U8266 ( n8472,n8466,n8479 );
   nand U8267 ( n8479,n8480,n8481 );
   nand U8268 ( n8481,n6001,n8482 );
   xor U8269 ( n8482,n8467,n8465 );
   nand U8270 ( n8467,n8483,n8484 );
   nand U8271 ( n8484,reg1_reg_10_,n8485 );
   or U8272 ( n8485,n8486,n8487 );
   nand U8273 ( n8483,n8487,n8486 );
   nor U8274 ( n8480,n5988,n8488 );
   nor U8275 ( n8488,n8282,n8477 );
   xor U8276 ( n8477,n8458,n8457 );
   nand U8277 ( n8458,n8489,n8490 );
   nand U8278 ( n8490,n8491,n8492 );
   or U8279 ( n8491,n8493,n8494 );
   nand U8280 ( n8489,n8494,n8493 );
   not U8281 ( n8466,n8459 );
   nand U8282 ( n8496,n8497,n8498 );
   nand U8283 ( n8498,addr_reg_10_,n8268 );
   nand U8284 ( n8497,reg3_reg_10_,n5932 );
   nand U8285 ( n8495,n8499,n8500 );
   nand U8286 ( n8500,n8487,n8501 );
   nand U8287 ( n8501,n8502,n8503 );
   nand U8288 ( n8503,n6001,n8504 );
   xor U8289 ( n8504,n8486,n8505 );
   nor U8290 ( n8502,n8280,n8506 );
   nor U8291 ( n8506,n5980,n8507 );
   not U8292 ( n8487,n8493 );
   nand U8293 ( n8499,n8508,n8493 );
   nand U8294 ( n8508,n8509,n8510 );
   nand U8295 ( n8510,n8245,n8507 );
   xor U8296 ( n8507,n8494,n8492 );
   nand U8297 ( n8494,n8511,n8512 );
   nand U8298 ( n8512,n8513,n8514 );
   or U8299 ( n8513,n8515,n8516 );
   nand U8300 ( n8511,n8516,n8515 );
   nand U8301 ( n8509,n8517,n6001 );
   xor U8302 ( n8517,reg1_reg_10_,n8486 );
   nand U8303 ( n8486,n8518,n8519 );
   nand U8304 ( n8519,reg1_reg_9_,n8520 );
   or U8305 ( n8520,n8521,n8522 );
   nand U8306 ( n8518,n8522,n8521 );
   nand U8307 ( n8524,n8525,n8526 );
   nand U8308 ( n8526,addr_reg_9_,n5449 );
   nand U8309 ( n8525,reg3_reg_9_,n5973 );
   nand U8310 ( n8523,n8527,n8528 );
   nand U8311 ( n8528,n8516,n8529 );
   nand U8312 ( n8529,n8530,n8531 );
   nand U8313 ( n8531,n8245,n8532 );
   nand U8314 ( n8530,n8533,n8256 );
   xor U8315 ( n8533,reg1_reg_9_,n8521 );
   nand U8316 ( n8527,n8522,n8534 );
   nand U8317 ( n8534,n8535,n8536 );
   nand U8318 ( n8536,n8256,n8537 );
   xor U8319 ( n8537,n8521,n8538 );
   nand U8320 ( n8521,n8539,n8540 );
   nand U8321 ( n8540,reg1_reg_8_,n8541 );
   or U8322 ( n8541,n8542,n8543 );
   nand U8323 ( n8539,n8543,n8542 );
   nor U8324 ( n8535,n5988,n8544 );
   nor U8325 ( n8544,n5980,n8532 );
   xor U8326 ( n8532,n8515,n8514 );
   nand U8327 ( n8515,n8545,n8546 );
   nand U8328 ( n8546,n8547,n8548 );
   or U8329 ( n8547,n8549,n8550 );
   nand U8330 ( n8545,n8550,n8549 );
   not U8331 ( n8522,n8516 );
   nand U8332 ( n8552,n8553,n8554 );
   nand U8333 ( n8554,addr_reg_8_,n8268 );
   nand U8334 ( n8553,reg3_reg_8_,n5975 );
   nand U8335 ( n8551,n8555,n8556 );
   nand U8336 ( n8556,n8543,n8557 );
   nand U8337 ( n8557,n8558,n8559 );
   nand U8338 ( n8559,n8256,n8560 );
   xor U8339 ( n8560,n8542,n8561 );
   nor U8340 ( n8558,n5988,n8562 );
   nor U8341 ( n8562,n8282,n8563 );
   not U8342 ( n8543,n8549 );
   nand U8343 ( n8555,n8564,n8549 );
   nand U8344 ( n8564,n8565,n8566 );
   nand U8345 ( n8566,n8245,n8563 );
   xor U8346 ( n8563,n8550,n8548 );
   nand U8347 ( n8550,n8567,n8568 );
   nand U8348 ( n8568,n8569,n8570 );
   or U8349 ( n8569,n8571,n8572 );
   nand U8350 ( n8567,n8572,n8571 );
   nand U8351 ( n8565,n8573,n6001 );
   xor U8352 ( n8573,reg1_reg_8_,n8542 );
   nand U8353 ( n8542,n8574,n8575 );
   nand U8354 ( n8575,reg1_reg_7_,n8576 );
   nand U8355 ( n8576,n8572,n8577 );
   or U8356 ( n8574,n8577,n8572 );
   nand U8357 ( n8579,n8580,n8581 );
   nand U8358 ( n8581,addr_reg_7_,n8268 );
   nand U8359 ( n8580,reg3_reg_7_,n5973 );
   nand U8360 ( n8578,n8582,n8583 );
   nand U8361 ( n8583,n8572,n8584 );
   nand U8362 ( n8584,n8585,n8586 );
   nand U8363 ( n8586,n8245,n8587 );
   nand U8364 ( n8585,n8256,n8588 );
   xor U8365 ( n8588,n8577,n8589 );
   nand U8366 ( n8582,n8590,n8591 );
   nand U8367 ( n8591,n8592,n8593 );
   nand U8368 ( n8593,n8594,n8256 );
   xor U8369 ( n8594,reg1_reg_7_,n8577 );
   nand U8370 ( n8577,n8595,n8596 );
   nand U8371 ( n8596,n8597,n8598 );
   nand U8372 ( n8597,n8599,n8600 );
   or U8373 ( n8595,n8600,n8599 );
   nor U8374 ( n8592,n5988,n8601 );
   nor U8375 ( n8601,n5980,n8587 );
   xor U8376 ( n8587,n8571,n8570 );
   nand U8377 ( n8571,n8602,n8603 );
   nand U8378 ( n8603,n8604,n8605 );
   or U8379 ( n8604,n8606,n8607 );
   nand U8380 ( n8602,n8607,n8606 );
   not U8381 ( n8590,n8572 );
   nand U8382 ( n8609,n8610,n8611 );
   nand U8383 ( n8611,addr_reg_6_,n8268 );
   nand U8384 ( n8610,reg3_reg_6_,n5975 );
   nand U8385 ( n8608,n8612,n8613 );
   nand U8386 ( n8613,n8599,n8614 );
   nand U8387 ( n8614,n8615,n8616 );
   nand U8388 ( n8616,n6001,n8617 );
   xor U8389 ( n8617,n8600,n8598 );
   nor U8390 ( n8615,n5988,n8618 );
   nor U8391 ( n8618,n5980,n8619 );
   not U8392 ( n8599,n8606 );
   nand U8393 ( n8612,n8620,n8606 );
   nand U8394 ( n8620,n8621,n8622 );
   nand U8395 ( n8622,n8245,n8619 );
   xor U8396 ( n8619,n8607,n8605 );
   nand U8397 ( n8607,n8623,n8624 );
   nand U8398 ( n8624,n8625,n8626 );
   or U8399 ( n8625,n8627,n8628 );
   nand U8400 ( n8623,n8628,n8627 );
   nand U8401 ( n8621,n8629,n8256 );
   xor U8402 ( n8629,reg1_reg_6_,n8600 );
   nand U8403 ( n8600,n8630,n8631 );
   nand U8404 ( n8631,reg1_reg_5_,n8632 );
   or U8405 ( n8632,n8633,n8634 );
   nand U8406 ( n8630,n8634,n8633 );
   nand U8407 ( n8636,n8637,n8638 );
   nand U8408 ( n8638,addr_reg_5_,n5449 );
   nand U8409 ( n8637,reg3_reg_5_,n5973 );
   nand U8410 ( n8635,n8639,n8640 );
   nand U8411 ( n8640,n8628,n8641 );
   nand U8412 ( n8641,n8642,n8643 );
   nand U8413 ( n8643,n8245,n8644 );
   nand U8414 ( n8642,n8645,n6001 );
   xor U8415 ( n8645,reg1_reg_5_,n8633 );
   nand U8416 ( n8639,n8634,n8646 );
   nand U8417 ( n8646,n8647,n8648 );
   nand U8418 ( n8648,n6001,n8649 );
   xor U8419 ( n8649,n8633,n8650 );
   nand U8420 ( n8633,n8651,n8652 );
   nand U8421 ( n8652,reg1_reg_4_,n8653 );
   or U8422 ( n8653,n8654,n8655 );
   nand U8423 ( n8651,n8655,n8654 );
   nor U8424 ( n8647,n5988,n8656 );
   nor U8425 ( n8656,n8282,n8644 );
   xor U8426 ( n8644,n8627,n8626 );
   nand U8427 ( n8627,n8657,n8658 );
   nand U8428 ( n8658,n8659,n8660 );
   or U8429 ( n8659,n8661,n8662 );
   nand U8430 ( n8657,n8662,n8661 );
   not U8431 ( n8634,n8628 );
   and U8432 ( n8664,n8665,n8666 );
   nand U8433 ( n8665,addr_reg_4_,n8268 );
   nor U8434 ( n8663,n8667,n8668 );
   nand U8435 ( n8668,n8669,n8670 );
   nand U8436 ( n8670,n8655,n8671 );
   nand U8437 ( n8671,n8672,n8673 );
   nand U8438 ( n8673,n8256,n8674 );
   xor U8439 ( n8674,n8654,n8675 );
   nor U8440 ( n8672,n5988,n8676 );
   nor U8441 ( n8676,n5980,n8677 );
   not U8442 ( n8655,n8661 );
   nand U8443 ( n8669,n8678,n8661 );
   nand U8444 ( n8678,n8679,n8680 );
   nand U8445 ( n8680,n8245,n8677 );
   xor U8446 ( n8677,n8662,n8660 );
   nand U8447 ( n8662,n8681,n8682 );
   nand U8448 ( n8682,n8683,n8684 );
   or U8449 ( n8683,n8685,n8686 );
   nand U8450 ( n8681,n8686,n8685 );
   nand U8451 ( n8679,n8687,n8256 );
   xor U8452 ( n8687,reg1_reg_4_,n8654 );
   nand U8453 ( n8654,n8688,n8689 );
   nand U8454 ( n8689,n8690,n8691 );
   nand U8455 ( n8693,n8694,n8695 );
   nand U8456 ( n8695,addr_reg_3_,n8268 );
   nand U8457 ( n8692,n8696,n8697 );
   nand U8458 ( n8697,n8690,n8698 );
   nand U8459 ( n8698,n8699,n8700 );
   nand U8460 ( n8700,n6001,n8701 );
   nand U8461 ( n8701,n8688,n8691 );
   nor U8462 ( n8699,n5988,n8702 );
   nor U8463 ( n8702,n5980,n8703 );
   nand U8464 ( n8696,n8686,n8704 );
   nand U8465 ( n8704,n8705,n8706 );
   nand U8466 ( n8706,n8707,n6001 );
   and U8467 ( n8707,n8688,n8691 );
   nand U8468 ( n8691,n8708,n8709 );
   nand U8469 ( n8709,n8710,n8711 );
   nor U8470 ( n8708,reg1_reg_3_,n8712 );
   nor U8471 ( n8712,n8713,n8714 );
   nand U8472 ( n8688,n8715,reg1_reg_3_ );
   nor U8473 ( n8715,n8716,n8713 );
   nor U8474 ( n8713,n8710,n8711 );
   nor U8475 ( n8716,reg1_reg_2_,n8717 );
   nor U8476 ( n8717,n8718,n8719 );
   nand U8477 ( n8705,n8245,n8703 );
   xor U8478 ( n8703,n8685,n8684 );
   nand U8479 ( n8685,n8720,n8721 );
   nand U8480 ( n8721,n8722,n8723 );
   or U8481 ( n8722,n8724,n8718 );
   nand U8482 ( n8720,n8718,n8724 );
   and U8483 ( n8726,n8727,n8666 );
   nand U8484 ( n8666,n10807,n8728 );
   nand U8485 ( n8728,n8729,n8730 );
   nand U8486 ( n8730,n8731,n8732 );
   nor U8487 ( n8731,n8733,n8734 );
   nand U8488 ( n8729,n8735,n8736 );
   nand U8489 ( n8736,n8732,n8737 );
   nand U8490 ( n8737,n8734,n8738 );
   nand U8491 ( n8735,n8739,n8740 );
   nand U8492 ( n8739,n8732,reg2_reg_0_ );
   not U8493 ( n10807,n6016 );
   nand U8494 ( n8727,addr_reg_2_,n8268 );
   nor U8495 ( n8725,n8741,n8742 );
   nand U8496 ( n8742,n8743,n8744 );
   nand U8497 ( n8744,n8718,n8745 );
   nand U8498 ( n8745,n8746,n8747 );
   nand U8499 ( n8747,n8245,n8748 );
   nand U8500 ( n8746,n6001,n8749 );
   xor U8501 ( n8749,n8710,reg1_reg_2_ );
   nand U8502 ( n8743,n8711,n8750 );
   nand U8503 ( n8750,n8751,n8752 );
   nand U8504 ( n8752,n8753,n6001 );
   xor U8505 ( n8753,n8714,n8710 );
   not U8506 ( n8710,n8719 );
   nand U8507 ( n8719,n8754,n8755 );
   nand U8508 ( n8755,n8756,n8757 );
   nand U8509 ( n8756,n8758,n8759 );
   nand U8510 ( n8754,n8760,n8761 );
   nor U8511 ( n8751,n5988,n8762 );
   nor U8512 ( n8762,n5980,n8748 );
   xor U8513 ( n8748,n8724,n8723 );
   nand U8514 ( n8724,n8763,n8764 );
   nand U8515 ( n8764,n8765,n8766 );
   or U8516 ( n8765,n8738,n8760 );
   nand U8517 ( n8763,n8760,n8738 );
   not U8518 ( n8711,n8718 );
   nor U8519 ( n8741,state_reg,n8767 );
   nor U8520 ( n8769,n8770,n8771 );
   nor U8521 ( n8771,n8772,n8759 );
   nor U8522 ( n8772,n8773,n8774 );
   nand U8523 ( n8774,n8775,n8776 );
   nand U8524 ( n8776,n8777,n8757 );
   and U8525 ( n8777,n8758,n6001 );
   nand U8526 ( n8775,n8778,reg1_reg_1_ );
   nand U8527 ( n8773,n8779,n8780 );
   nand U8528 ( n8780,n8781,n8766 );
   nand U8529 ( n8779,n8782,reg2_reg_1_ );
   nor U8530 ( n8770,n8783,n8760 );
   nor U8531 ( n8783,n8784,n8785 );
   nand U8532 ( n8785,n8786,n8265 );
   not U8533 ( n8265,n8280 );
   nor U8534 ( n8786,n8787,n8788 );
   nor U8535 ( n8788,n8757,n8789 );
   nand U8536 ( n8789,n8256,n8758 );
   nor U8537 ( n8787,reg1_reg_1_,n8790 );
   nand U8538 ( n8784,n8791,n8792 );
   nand U8539 ( n8792,n8782,n8766 );
   nand U8540 ( n8791,n8781,reg2_reg_1_ );
   nor U8541 ( n8781,n8738,n5980 );
   nor U8542 ( n8768,n8793,n8794 );
   nor U8543 ( n8794,state_reg,n8795 );
   and U8544 ( n8793,addr_reg_1_,n8268 );
   nor U8545 ( n8797,n8798,n8799 );
   nand U8546 ( n8799,n8800,n8801 );
   nand U8547 ( n8801,n8782,reg2_reg_0_ );
   not U8548 ( n8782,n8802 );
   nand U8549 ( n8800,n8778,reg1_reg_0_ );
   not U8550 ( n8778,n8790 );
   nor U8551 ( n8798,n8803,n8740 );
   nor U8552 ( n8803,n8280,n8804 );
   nand U8553 ( n8804,n8802,n8790 );
   nand U8554 ( n8790,n8256,n8761 );
   not U8555 ( n8761,n8758 );
   nor U8556 ( n8758,n8740,n8805 );
   nor U8557 ( n8256,n8734,n8806 );
   nand U8558 ( n8802,n8245,n8738 );
   nand U8559 ( n8738,ir_reg_0_,reg2_reg_0_ );
   not U8560 ( n8245,n5980 );
   nand U8561 ( n8282,n8807,n8732 );
   and U8562 ( n8807,n8808,n8734 );
   nor U8563 ( n8280,n8732,n8806 );
   not U8564 ( n8806,n8808 );
   nand U8565 ( n8808,n8809,n8810 );
   nand U8566 ( n8810,n8811,n8812 );
   nor U8567 ( n8811,n5973,n8268 );
   nand U8568 ( n8809,n8813,n6210 );
   nor U8569 ( n8813,n8268,n8814 );
   nor U8570 ( n8814,n8815,n8816 );
   nand U8571 ( n8816,n8817,n8818 );
   and U8572 ( n8818,n8029,n8819 );
   nor U8573 ( n8817,n6254,n7814 );
   not U8574 ( n7814,n8820 );
   nand U8575 ( n8815,n8821,n8822 );
   nor U8576 ( n8822,n7523,n6218 );
   not U8577 ( n7523,n7769 );
   nor U8578 ( n8821,n8118,n8823 );
   nor U8579 ( n8796,n8824,n8825 );
   nor U8580 ( n8825,state_reg,n6996 );
   and U8581 ( n8824,addr_reg_0_,n8268 );
   nor U8582 ( n8268,n8826,n5939 );
   nand U8583 ( n8828,n8829,state_reg );
   nand U8584 ( n8829,n8830,n8831 );
   nand U8585 ( n8831,n8832,n5970 );
   nor U8586 ( n8832,n8833,n8247 );
   nand U8587 ( n8830,n8812,n8834 );
   nand U8588 ( n8834,n8835,n8836 );
   nor U8589 ( n8836,n8837,n8838 );
   nor U8590 ( n8838,n8029,n8833 );
   nor U8591 ( n8837,n8035,n8839 );
   nand U8592 ( n8839,n8840,n8841 );
   nor U8593 ( n8835,n8842,n8843 );
   nand U8594 ( n8843,n8844,n8845 );
   nand U8595 ( n8845,n7835,n8846 );
   nand U8596 ( n8844,n8847,n8848 );
   not U8597 ( n8848,n8846 );
   nand U8598 ( n8846,n8849,n8850 );
   nor U8599 ( n8850,n8851,n8852 );
   nand U8600 ( n8852,n8853,n8854 );
   nand U8601 ( n8853,n8855,n8856 );
   nor U8602 ( n8856,n8857,n7958 );
   nor U8603 ( n8857,n8058,n8858 );
   nor U8604 ( n8858,n8859,n8860 );
   nor U8605 ( n8860,n8861,n8862 );
   nor U8606 ( n8859,n8863,n8864 );
   nand U8607 ( n8864,n8865,n8866 );
   nor U8608 ( n8866,n8867,n8868 );
   nand U8609 ( n8868,n8869,n8870 );
   nand U8610 ( n8870,n8871,n8872 );
   nor U8611 ( n8871,n7566,n8081 );
   nand U8612 ( n8869,n7346,n8873 );
   nor U8613 ( n8867,n8874,n8875 );
   nor U8614 ( n8874,n8876,n8877 );
   nand U8615 ( n8877,n8878,n7402 );
   nand U8616 ( n8878,n8879,n8880 );
   nor U8617 ( n8879,n8881,n8882 );
   nor U8618 ( n8865,n8883,n8884 );
   not U8619 ( n8884,n8112 );
   nor U8620 ( n8112,n7821,n8885 );
   and U8621 ( n8885,n7818,n7804 );
   nand U8622 ( n7821,n7761,n8886 );
   and U8623 ( n8883,n8887,n8872 );
   nand U8624 ( n8863,n8888,n8889 );
   nor U8625 ( n8889,n8890,n8891 );
   nand U8626 ( n8891,n8110,n8892 );
   nand U8627 ( n8892,n8893,n8873 );
   nor U8628 ( n8893,n8894,n8882 );
   nand U8629 ( n8882,n8895,n8095 );
   nor U8630 ( n8095,n7229,n8106 );
   nor U8631 ( n8895,n7314,n7347 );
   nor U8632 ( n8894,n8896,n8897 );
   nand U8633 ( n8897,n8898,n8899 );
   nand U8634 ( n8899,n8900,n7279 );
   not U8635 ( n7279,n8881 );
   nand U8636 ( n8881,n8901,n7196 );
   not U8637 ( n7196,n7153 );
   and U8638 ( n8901,n7126,n7194 );
   nor U8639 ( n8900,n8902,n7092 );
   nor U8640 ( n7092,n7066,n7056 );
   nor U8641 ( n7056,n7051,n7067 );
   nand U8642 ( n7051,n8903,n8904 );
   nand U8643 ( n8904,n7023,n8905 );
   nand U8644 ( n8903,n6650,n7011 );
   nand U8645 ( n8898,n7154,n7194 );
   nand U8646 ( n8896,n8906,n7283 );
   nand U8647 ( n7283,n8102,n7194 );
   nor U8648 ( n8102,n7127,n7153 );
   nor U8649 ( n8890,n8907,n8908 );
   nand U8650 ( n8908,n8873,n7395 );
   not U8651 ( n8873,n8875 );
   nand U8652 ( n8875,n8909,n8910 );
   nor U8653 ( n8910,n8081,n8911 );
   nand U8654 ( n8911,n8912,n7568 );
   or U8655 ( n8912,n7401,n8876 );
   nand U8656 ( n8081,n7531,n7565 );
   nor U8657 ( n8909,n8913,n8914 );
   nand U8658 ( n8907,n8915,n8916 );
   nor U8659 ( n8888,n8917,n8918 );
   nand U8660 ( n8918,n8919,n8920 );
   nand U8661 ( n8920,n8921,n8922 );
   and U8662 ( n8921,n7565,n8872 );
   not U8663 ( n8872,n8913 );
   nand U8664 ( n8919,n8923,n7817 );
   nor U8665 ( n8917,n8913,n8073 );
   nand U8666 ( n8913,n8924,n7832 );
   nor U8667 ( n7832,n8925,n7682 );
   nor U8668 ( n8924,n8065,n8926 );
   and U8669 ( n8855,n8057,n8927 );
   nor U8670 ( n8851,n8928,n8929 );
   nand U8671 ( n8928,n6017,n8930 );
   nor U8672 ( n8849,n8931,n8932 );
   nand U8673 ( n8932,n8933,n8934 );
   nand U8674 ( n8934,n8935,n8936 );
   and U8675 ( n8935,n8930,n8937 );
   nand U8676 ( n8933,n8927,n8938 );
   nand U8677 ( n8938,n8055,n7934 );
   nor U8678 ( n8927,n8939,n8940 );
   or U8679 ( n8939,n8053,n6713 );
   nor U8680 ( n8931,n8941,n8940 );
   nand U8681 ( n8940,n8942,n8937 );
   nand U8682 ( n8937,n6229,n8943 );
   nand U8683 ( n8943,n6020,n6017 );
   nor U8684 ( n8942,n8944,n8945 );
   nor U8685 ( n8847,n6667,n7287 );
   not U8686 ( n7287,n7058 );
   nand U8687 ( n8842,n8946,n8947 );
   nand U8688 ( n8947,n8247,n8948 );
   nand U8689 ( n8948,n8949,n8950 );
   nand U8690 ( n8950,n8951,n6664 );
   nor U8691 ( n8949,n8952,n8953 );
   nor U8692 ( n8953,n8041,n8954 );
   xor U8693 ( n8954,n8955,n8956 );
   and U8694 ( n8955,n8840,n8841 );
   nand U8695 ( n8841,n8957,n8958 );
   nand U8696 ( n8958,n8959,n8960 );
   nor U8697 ( n8957,n8961,n8962 );
   nor U8698 ( n8962,n8963,n8964 );
   nor U8699 ( n8961,n8965,n8966 );
   nand U8700 ( n8966,n8967,n8968 );
   nand U8701 ( n8968,n8969,n8970 );
   nand U8702 ( n8970,n8971,n8972 );
   nor U8703 ( n8969,n8973,n8974 );
   nor U8704 ( n8974,n8975,n8976 );
   nand U8705 ( n8976,n8977,n8978 );
   nand U8706 ( n8978,n8011,n6272 );
   nand U8707 ( n8977,n8979,n8980 );
   nand U8708 ( n8975,n8981,n8941 );
   nand U8709 ( n8981,n8982,n8983 );
   or U8710 ( n8983,n8980,n8979 );
   and U8711 ( n8979,n8984,n8985 );
   nand U8712 ( n8985,n5970,n7972 );
   nand U8713 ( n8984,n5951,n6029 );
   nand U8714 ( n8980,n8986,n8987 );
   nand U8715 ( n8987,n5970,n6029 );
   nand U8716 ( n8986,n7972,n5951 );
   nor U8717 ( n8982,n8988,n8989 );
   nor U8718 ( n8989,n8990,n8991 );
   nand U8719 ( n8991,n8992,n8993 );
   nand U8720 ( n8993,n8994,n8995 );
   nand U8721 ( n8995,n8996,n8997 );
   nor U8722 ( n8994,n8998,n8999 );
   nor U8723 ( n8999,n9000,n9001 );
   nand U8724 ( n9001,n9002,n9003 );
   nand U8725 ( n9003,n9004,n9005 );
   nand U8726 ( n9005,n9006,n9007 );
   nor U8727 ( n9004,n9008,n9009 );
   nor U8728 ( n9009,n7763,n9010 );
   nand U8729 ( n9010,n9011,n9012 );
   nand U8730 ( n9012,n9013,n9014 );
   nand U8731 ( n9014,n9015,n9016 );
   nor U8732 ( n9013,n9017,n9018 );
   nor U8733 ( n9018,n9019,n9020 );
   nand U8734 ( n9020,n9021,n9022 );
   nand U8735 ( n9022,n9023,n9024 );
   nand U8736 ( n9024,n9025,n9026 );
   nor U8737 ( n9023,n9027,n9028 );
   nor U8738 ( n9028,n9029,n9030 );
   nand U8739 ( n9030,n9031,n9032 );
   nand U8740 ( n9032,n9033,n9034 );
   nand U8741 ( n9034,n9035,n9036 );
   nor U8742 ( n9033,n9037,n9038 );
   nor U8743 ( n9038,n9039,n9040 );
   nand U8744 ( n9040,n9041,n9042 );
   nand U8745 ( n9042,n9043,n9044 );
   nor U8746 ( n9044,n9045,n9046 );
   nor U8747 ( n9046,n7496,n9047 );
   nand U8748 ( n9047,n9048,n9049 );
   nor U8749 ( n9049,n9050,n9051 );
   nand U8750 ( n9051,n7566,n9052 );
   nand U8751 ( n9052,n9053,n9054 );
   not U8752 ( n9054,n9055 );
   nor U8753 ( n9053,n9056,n9057 );
   not U8754 ( n9056,n9058 );
   nor U8755 ( n9050,n9059,n9060 );
   nand U8756 ( n9060,n9061,n9062 );
   nor U8757 ( n9048,n9063,n9064 );
   nor U8758 ( n9064,n9065,n9066 );
   nor U8759 ( n9063,n9067,n9068 );
   nand U8760 ( n9068,n9061,n9069 );
   nand U8761 ( n9069,n9070,n9059 );
   nand U8762 ( n9059,n9071,n9072 );
   nand U8763 ( n9072,n5969,n7381 );
   nand U8764 ( n9071,n5951,n6077 );
   not U8765 ( n9070,n9062 );
   nand U8766 ( n9062,n9073,n9074 );
   nand U8767 ( n9074,n5968,n6077 );
   nand U8768 ( n9073,n7381,n5950 );
   and U8769 ( n9061,n9058,n9075 );
   nand U8770 ( n9075,n9057,n9055 );
   nand U8771 ( n9055,n9076,n9077 );
   nand U8772 ( n9077,n5968,n7411 );
   nand U8773 ( n9076,n5951,n6074 );
   and U8774 ( n9057,n9078,n9079 );
   nand U8775 ( n9079,n5971,n6074 );
   nand U8776 ( n9078,n7411,n8819 );
   nand U8777 ( n9058,n9065,n9066 );
   nand U8778 ( n9066,n9080,n9081 );
   nand U8779 ( n9081,n8819,n6071 );
   nand U8780 ( n9080,n5971,n7442 );
   and U8781 ( n9065,n9082,n9083 );
   nand U8782 ( n9083,n5970,n6071 );
   nand U8783 ( n9082,n7442,n5950 );
   nand U8784 ( n9067,n9084,n9085 );
   nand U8785 ( n9085,n9086,n9087 );
   or U8786 ( n9087,n9088,n9089 );
   nor U8787 ( n9086,n9090,n9091 );
   nor U8788 ( n9091,n5949,n6513 );
   nor U8789 ( n9090,n6524,n5967 );
   nand U8790 ( n9084,n9089,n9088 );
   nand U8791 ( n9088,n9093,n9094 );
   nand U8792 ( n9094,n5971,n7327 );
   nand U8793 ( n9093,n5950,n6080 );
   nand U8794 ( n9089,n9095,n9096 );
   nand U8795 ( n9096,n9097,n9098 );
   nand U8796 ( n9098,n9099,n9100 );
   nand U8797 ( n9097,n9101,n9102 );
   nand U8798 ( n9102,n8819,n6083 );
   nand U8799 ( n9101,n5969,n7302 );
   or U8800 ( n9095,n9100,n9099 );
   and U8801 ( n9099,n9103,n9104 );
   nand U8802 ( n9104,n9105,n9106 );
   nand U8803 ( n9103,n9107,n9108 );
   nor U8804 ( n9108,n9109,n9110 );
   nor U8805 ( n9110,n9111,n9112 );
   nand U8806 ( n9112,n9113,n9114 );
   nand U8807 ( n9114,n9115,n9116 );
   not U8808 ( n9115,n9117 );
   nand U8809 ( n9113,n9118,n9119 );
   nand U8810 ( n9111,n9120,n9121 );
   nand U8811 ( n9121,n9122,n9123 );
   or U8812 ( n9123,n9119,n9118 );
   nand U8813 ( n9118,n9124,n9125 );
   nand U8814 ( n9125,n9126,n9127 );
   nand U8815 ( n9127,n9128,n9129 );
   nand U8816 ( n9126,n9130,n9131 );
   nand U8817 ( n9131,n5951,n6101 );
   nand U8818 ( n9130,n5969,n7079 );
   or U8819 ( n9124,n9129,n9128 );
   and U8820 ( n9128,n9132,n9133 );
   nand U8821 ( n9133,n9134,n9135 );
   nand U8822 ( n9135,n9136,n9137 );
   nor U8823 ( n9134,n9138,n9139 );
   nor U8824 ( n9139,n9140,n9141 );
   nand U8825 ( n9141,n9142,n9143 );
   nor U8826 ( n9138,n9144,n9145 );
   nand U8827 ( n9145,n9146,n9147 );
   nand U8828 ( n9147,n5950,n6110 );
   or U8829 ( n9146,n9137,n9136 );
   and U8830 ( n9136,n9148,n9149 );
   nand U8831 ( n9149,n5970,n7011 );
   nand U8832 ( n9148,n8819,n6107 );
   nand U8833 ( n9137,n9150,n9151 );
   nand U8834 ( n9151,n5970,n6107 );
   nand U8835 ( n9150,n7011,n5951 );
   nand U8836 ( n9144,n9152,n9153 );
   nand U8837 ( n9152,n5968,n6987 );
   nand U8838 ( n9132,n9154,n9155 );
   nand U8839 ( n9155,n9156,n9142 );
   nand U8840 ( n9142,n9157,n6104 );
   not U8841 ( n9156,n9140 );
   nand U8842 ( n9140,n9158,n9159 );
   nand U8843 ( n9159,n5968,n7032 );
   nand U8844 ( n9158,n9160,n6104 );
   not U8845 ( n9154,n9143 );
   nand U8846 ( n9143,n9161,n9162 );
   nand U8847 ( n9162,n5970,n6104 );
   nand U8848 ( n9161,n7032,n8819 );
   nand U8849 ( n9129,n9163,n9164 );
   nand U8850 ( n9164,n5971,n6101 );
   nand U8851 ( n9163,n7079,n5950 );
   nand U8852 ( n9119,n9165,n9166 );
   nand U8853 ( n9166,n5971,n7106 );
   nand U8854 ( n9165,n5950,n6098 );
   nor U8855 ( n9122,n9167,n9168 );
   nor U8856 ( n9168,n9092,n6597 );
   nor U8857 ( n9167,n6608,n5967 );
   nor U8858 ( n9120,n9169,n9170 );
   not U8859 ( n9169,n9171 );
   nor U8860 ( n9109,n9172,n9173 );
   nand U8861 ( n9173,n9174,n9175 );
   nor U8862 ( n9172,n6555,n5967 );
   nor U8863 ( n9107,n9176,n9177 );
   nor U8864 ( n9177,n9105,n9106 );
   nand U8865 ( n9106,n9178,n9179 );
   nand U8866 ( n9179,n5969,n7256 );
   nand U8867 ( n9178,n8819,n6086 );
   and U8868 ( n9105,n9180,n9181 );
   nand U8869 ( n9181,n5969,n6086 );
   nand U8870 ( n9180,n7256,n8819 );
   nor U8871 ( n9176,n9170,n9182 );
   nor U8872 ( n9182,n9183,n9184 );
   nor U8873 ( n9184,n9185,n9186 );
   nor U8874 ( n9183,n9187,n9116 );
   nand U8875 ( n9116,n9188,n9189 );
   nand U8876 ( n9189,n9157,n6095 );
   and U8877 ( n9188,n9190,n9191 );
   nand U8878 ( n9191,n5969,n7141 );
   nand U8879 ( n9190,n9160,n6095 );
   nand U8880 ( n9187,n9117,n9171 );
   nand U8881 ( n9171,n9185,n9186 );
   nand U8882 ( n9186,n9192,n9193 );
   nand U8883 ( n9193,n5971,n7175 );
   nand U8884 ( n9192,n8819,n6092 );
   and U8885 ( n9185,n9194,n9195 );
   nand U8886 ( n9195,n5968,n6092 );
   nand U8887 ( n9194,n7175,n5951 );
   nand U8888 ( n9117,n9196,n9197 );
   nand U8889 ( n9197,n5970,n6095 );
   nand U8890 ( n9196,n7141,n8819 );
   nor U8891 ( n9170,n9175,n9198 );
   and U8892 ( n9198,n6555,n9174 );
   nand U8893 ( n9174,n8819,n6089 );
   nand U8894 ( n9175,n9199,n9200 );
   nand U8895 ( n9200,n5969,n6089 );
   nand U8896 ( n9199,n7216,n5950 );
   nand U8897 ( n9100,n9201,n9202 );
   nand U8898 ( n9202,n5969,n6083 );
   nand U8899 ( n9201,n7302,n8819 );
   nor U8900 ( n9045,n5951,n7568 );
   nor U8901 ( n9043,n9203,n9204 );
   nor U8902 ( n9204,n5969,n7566 );
   nor U8903 ( n9203,n9205,n9206 );
   nand U8904 ( n9041,n9205,n9206 );
   nand U8905 ( n9206,n9207,n9208 );
   nand U8906 ( n9208,n5970,n6065 );
   nand U8907 ( n9207,n7509,n5950 );
   and U8908 ( n9205,n9209,n9210 );
   nand U8909 ( n9210,n5968,n7509 );
   nand U8910 ( n9209,n5950,n6065 );
   nand U8911 ( n9039,n8078,n7565 );
   nor U8912 ( n9037,n9211,n9212 );
   nand U8913 ( n9212,n7599,n9213 );
   nand U8914 ( n9213,n5968,n6062 );
   nor U8915 ( n9211,n9092,n6429 );
   xor U8916 ( n9031,n7614,n6412 );
   nor U8917 ( n9029,n9035,n9036 );
   nand U8918 ( n9036,n9214,n9215 );
   nand U8919 ( n9215,n5969,n7582 );
   nand U8920 ( n9214,n5950,n6059 );
   and U8921 ( n9035,n9216,n9217 );
   nand U8922 ( n9217,n5971,n6059 );
   nand U8923 ( n9216,n7582,n5951 );
   nor U8924 ( n9027,n9218,n9219 );
   nand U8925 ( n9219,n7727,n9220 );
   nand U8926 ( n9220,n5968,n6056 );
   nor U8927 ( n9218,n9092,n6401 );
   or U8928 ( n9021,n9026,n9025 );
   and U8929 ( n9025,n9221,n9222 );
   nand U8930 ( n9222,n5968,n6053 );
   nand U8931 ( n9221,n7643,n5951 );
   nand U8932 ( n9026,n9223,n9224 );
   nand U8933 ( n9224,n5970,n7643 );
   nand U8934 ( n9223,n5950,n6053 );
   nand U8935 ( n9019,n8117,n8114 );
   nor U8936 ( n9017,n9225,n9226 );
   nand U8937 ( n9226,n8137,n9227 );
   nand U8938 ( n9227,n5970,n6050 );
   nor U8939 ( n9225,n9092,n6373 );
   or U8940 ( n9011,n9016,n9015 );
   and U8941 ( n9015,n9228,n9229 );
   nand U8942 ( n9229,n5969,n6047 );
   nand U8943 ( n9228,n7706,n8819 );
   nand U8944 ( n9016,n9230,n9231 );
   nand U8945 ( n9231,n5971,n7706 );
   nand U8946 ( n9230,n5951,n6047 );
   nand U8947 ( n7763,n7761,n7804 );
   not U8948 ( n7761,n7811 );
   nor U8949 ( n9008,n9232,n9233 );
   nand U8950 ( n9233,n8022,n9234 );
   nand U8951 ( n9234,n5968,n6044 );
   nor U8952 ( n9232,n9092,n6345 );
   or U8953 ( n9002,n9007,n9006 );
   and U8954 ( n9006,n9235,n9236 );
   nand U8955 ( n9236,n5971,n6041 );
   nand U8956 ( n9235,n7789,n5951 );
   nand U8957 ( n9007,n9237,n9238 );
   nand U8958 ( n9238,n5971,n7789 );
   nand U8959 ( n9237,n5950,n6041 );
   nand U8960 ( n9000,n8110,n8060 );
   not U8961 ( n8060,n9239 );
   not U8962 ( n8110,n8861 );
   nor U8963 ( n8998,n9240,n9241 );
   nand U8964 ( n9241,n9242,n9243 );
   nand U8965 ( n9243,n5968,n6038 );
   nand U8966 ( n9242,n6328,n6317 );
   nor U8967 ( n9240,n9092,n6317 );
   or U8968 ( n8992,n8997,n8996 );
   and U8969 ( n8996,n9244,n9245 );
   nand U8970 ( n9245,n5970,n6035 );
   nand U8971 ( n9244,n7879,n5950 );
   nand U8972 ( n8997,n9246,n9247 );
   nand U8973 ( n9247,n5971,n7879 );
   nand U8974 ( n9246,n5951,n6035 );
   nand U8975 ( n8990,n9248,n7934 );
   not U8976 ( n7934,n7957 );
   nor U8977 ( n8988,n9249,n9250 );
   nand U8978 ( n9250,n8196,n9251 );
   nand U8979 ( n9251,n5969,n6032 );
   nor U8980 ( n9249,n9092,n6289 );
   nor U8981 ( n8973,n9252,n9253 );
   nand U8982 ( n9253,n9254,n9255 );
   nand U8983 ( n9255,n5969,n6026 );
   nand U8984 ( n9254,n6272,n6261 );
   nor U8985 ( n9252,n9092,n6261 );
   or U8986 ( n8967,n8960,n8959 );
   and U8987 ( n8959,n9256,n9257 );
   nand U8988 ( n9257,n6229,n5951 );
   nand U8989 ( n9256,n5970,n6020 );
   nand U8990 ( n8960,n9258,n9259 );
   nand U8991 ( n9259,n9260,n6020 );
   nand U8992 ( n9260,n6667,n9261 );
   nand U8993 ( n9261,n9157,n6017 );
   nand U8994 ( n9258,n5968,n6229 );
   nor U8995 ( n8965,n8971,n8972 );
   nand U8996 ( n8972,n9262,n9263 );
   nand U8997 ( n9263,n5968,n6694 );
   nand U8998 ( n9262,n5951,n6023 );
   and U8999 ( n8971,n9264,n9265 );
   nand U9000 ( n9265,n6694,n5950 );
   nand U9001 ( n9264,n5971,n6023 );
   nand U9002 ( n8840,n8963,n8964 );
   nand U9003 ( n8964,n9266,n9267 );
   nand U9004 ( n9267,n5969,n6219 );
   nand U9005 ( n9266,n8819,n6017 );
   and U9006 ( n8963,n9268,n9269 );
   nand U9007 ( n9269,n6219,n5950 );
   nand U9008 ( n9268,n5971,n6017 );
   nor U9009 ( n8952,n6666,n9271 );
   nand U9010 ( n9271,n8833,n8956 );
   nand U9011 ( n8833,n9272,n9273 );
   nor U9012 ( n9273,n9274,n9275 );
   nand U9013 ( n9275,n9276,n8930 );
   not U9014 ( n8930,n8944 );
   nand U9015 ( n9276,n9277,n9278 );
   nor U9016 ( n9278,n9279,n9280 );
   nand U9017 ( n9280,n7127,n8905 );
   nand U9018 ( n8905,n6639,n6107 );
   nand U9019 ( n9279,n9281,n7057 );
   not U9020 ( n7057,n7066 );
   nor U9021 ( n9281,n7811,n8880 );
   nor U9022 ( n9277,n9282,n9283 );
   nand U9023 ( n9283,n9284,n9285 );
   nand U9024 ( n9282,n9286,n9287 );
   nor U9025 ( n9286,n9288,n9289 );
   nor U9026 ( n9289,n9290,n6987 );
   not U9027 ( n6987,n6647 );
   nor U9028 ( n9288,n7023,n6668 );
   nor U9029 ( n7023,n6110,n6647 );
   nor U9030 ( n9274,n9291,n9292 );
   nand U9031 ( n9292,n9284,n9293 );
   nand U9032 ( n9293,n9294,n9295 );
   nor U9033 ( n9295,n9296,n9297 );
   nand U9034 ( n9297,n9298,n9299 );
   nand U9035 ( n9299,n9300,n9301 );
   nand U9036 ( n9301,n7401,n9302 );
   nand U9037 ( n9302,n9303,n9304 );
   not U9038 ( n9304,n9305 );
   nand U9039 ( n9303,n7395,n9306 );
   nand U9040 ( n9306,n9307,n9308 );
   nor U9041 ( n9308,n7228,n7346 );
   nor U9042 ( n9307,n8915,n7194 );
   nand U9043 ( n7194,n7175,n6580 );
   not U9044 ( n7395,n7347 );
   nor U9045 ( n7347,n6080,n6513 );
   nand U9046 ( n7401,n6510,n7381 );
   nand U9047 ( n9298,n7153,n9309 );
   nor U9048 ( n7153,n6095,n6583 );
   nand U9049 ( n9296,n9310,n9311 );
   nand U9050 ( n9311,n9312,n7719 );
   not U9051 ( n7719,n7818 );
   nand U9052 ( n9312,n8117,n9313 );
   nand U9053 ( n9313,n9314,n8114 );
   not U9054 ( n8114,n8923 );
   nand U9055 ( n9314,n9315,n9316 );
   not U9056 ( n9316,n8926 );
   nand U9057 ( n8926,n9317,n9318 );
   nand U9058 ( n9318,n9319,n7614 );
   nor U9059 ( n9319,n8116,n6056 );
   nand U9060 ( n9317,n8079,n9320 );
   nor U9061 ( n8079,n6059,n6415 );
   nor U9062 ( n9315,n7682,n9321 );
   nor U9063 ( n9321,n7565,n9322 );
   nand U9064 ( n9322,n9320,n8073 );
   not U9065 ( n8073,n9323 );
   nand U9066 ( n7565,n7542,n6440 );
   nor U9067 ( n7682,n6053,n6387 );
   not U9068 ( n8117,n8925 );
   nor U9069 ( n8925,n6373,n6050 );
   nand U9070 ( n9310,n9324,n9325 );
   nand U9071 ( n9325,n7531,n9326 );
   nand U9072 ( n9326,n9327,n7530 );
   not U9073 ( n7530,n8922 );
   nand U9074 ( n9327,n7568,n9328 );
   nand U9075 ( n9328,n8914,n7566 );
   not U9076 ( n7566,n7495 );
   nand U9077 ( n8914,n8084,n9329 );
   nand U9078 ( n9329,n8086,n8082 );
   nand U9079 ( n8084,n7442,n6482 );
   not U9080 ( n7568,n7496 );
   nor U9081 ( n7496,n6457,n6068 );
   nand U9082 ( n7531,n6454,n7509 );
   not U9083 ( n9324,n9330 );
   nor U9084 ( n9294,n9331,n9332 );
   nand U9085 ( n9332,n7817,n9333 );
   nand U9086 ( n9333,n9287,n9334 );
   nand U9087 ( n9334,n7126,n9335 );
   nand U9088 ( n9335,n9336,n7127 );
   nand U9089 ( n7127,n6597,n6098 );
   nand U9090 ( n9336,n8097,n9337 );
   nand U9091 ( n9337,n9338,n8098 );
   not U9092 ( n8098,n8880 );
   nor U9093 ( n8880,n7079,n6622 );
   nand U9094 ( n9338,n9339,n9340 );
   nand U9095 ( n9340,n9341,n6650 );
   nor U9096 ( n9341,n7066,n6639 );
   nor U9097 ( n7066,n7032,n6636 );
   not U9098 ( n9339,n7067 );
   nor U9099 ( n7067,n6625,n6104 );
   not U9100 ( n8097,n8902 );
   nor U9101 ( n8902,n6611,n6101 );
   nand U9102 ( n7126,n6608,n7106 );
   and U9103 ( n9287,n9309,n7198 );
   not U9104 ( n7198,n7154 );
   nor U9105 ( n7154,n7141,n6594 );
   and U9106 ( n9309,n9342,n8906 );
   nor U9107 ( n8906,n8103,n7228 );
   nor U9108 ( n7228,n7216,n6566 );
   nor U9109 ( n8103,n7175,n6580 );
   nor U9110 ( n9342,n9343,n8915 );
   not U9111 ( n7817,n8065 );
   nand U9112 ( n8065,n7718,n7804 );
   nand U9113 ( n7804,n7740,n6356 );
   nand U9114 ( n7718,n7706,n6370 );
   not U9115 ( n9331,n8862 );
   not U9116 ( n9284,n9344 );
   nor U9117 ( n9272,n9345,n9346 );
   nand U9118 ( n9346,n9347,n9348 );
   nand U9119 ( n9348,n9349,n9350 );
   nand U9120 ( n9350,n9351,n9352 );
   nand U9121 ( n9352,n8053,n8941 );
   nor U9122 ( n8053,n6275,n6029 );
   not U9123 ( n9351,n6713 );
   nor U9124 ( n6713,n6026,n6261 );
   nand U9125 ( n9347,n9353,n8854 );
   nand U9126 ( n9353,n9354,n9355 );
   nand U9127 ( n9355,n6727,n9356 );
   or U9128 ( n9356,n6229,n8945 );
   nand U9129 ( n9354,n8945,n6229 );
   nor U9130 ( n9345,n9357,n9344 );
   nand U9131 ( n9344,n9358,n9349 );
   nor U9132 ( n9349,n9359,n8936 );
   and U9133 ( n9358,n8941,n8055 );
   nand U9134 ( n8055,n6275,n6029 );
   not U9135 ( n8941,n6711 );
   nor U9136 ( n6711,n8011,n6272 );
   nor U9137 ( n9357,n9360,n9361 );
   nand U9138 ( n9361,n9362,n9248 );
   not U9139 ( n9248,n7958 );
   nor U9140 ( n7958,n6289,n6032 );
   nand U9141 ( n9362,n9363,n9364 );
   not U9142 ( n9364,n9291 );
   nand U9143 ( n9291,n9285,n9365 );
   nand U9144 ( n9365,n8862,n7811 );
   nor U9145 ( n7811,n6356,n7740 );
   nor U9146 ( n8862,n9239,n8064 );
   nor U9147 ( n8064,n6041,n6331 );
   and U9148 ( n9285,n9366,n9367 );
   nor U9149 ( n9367,n7957,n8058 );
   nor U9150 ( n8058,n6314,n7879 );
   nor U9151 ( n9366,n8861,n9368 );
   nor U9152 ( n9368,n9239,n8886 );
   nand U9153 ( n8886,n6331,n6041 );
   nor U9154 ( n9239,n6317,n6038 );
   nor U9155 ( n8861,n6328,n7844 );
   nor U9156 ( n9363,n9369,n9343 );
   nand U9157 ( n9343,n9370,n9300 );
   and U9158 ( n9300,n9371,n9372 );
   nor U9159 ( n9372,n7495,n8922 );
   nor U9160 ( n8922,n7509,n6454 );
   nor U9161 ( n7495,n7473,n6468 );
   nor U9162 ( n9371,n8876,n9330 );
   nand U9163 ( n9330,n9373,n9374 );
   nor U9164 ( n9374,n8923,n7818 );
   nor U9165 ( n7818,n6370,n7706 );
   nor U9166 ( n8923,n7662,n6384 );
   nor U9167 ( n9373,n9323,n8887 );
   nand U9168 ( n8887,n9320,n8078 );
   nand U9169 ( n8078,n6429,n6062 );
   and U9170 ( n9320,n7679,n9375 );
   nand U9171 ( n9375,n6401,n6056 );
   not U9172 ( n7679,n8116 );
   nor U9173 ( n8116,n7643,n6398 );
   nor U9174 ( n9323,n7582,n6426 );
   nand U9175 ( n8876,n8082,n8088 );
   nand U9176 ( n8088,n6485,n6074 );
   nand U9177 ( n8082,n6471,n6071 );
   nor U9178 ( n9370,n9305,n7346 );
   nor U9179 ( n7346,n7327,n6524 );
   nor U9180 ( n9305,n7402,n8086 );
   nor U9181 ( n8086,n6485,n6074 );
   nand U9182 ( n7402,n6499,n6077 );
   nor U9183 ( n9369,n9376,n9377 );
   nand U9184 ( n9377,n9378,n8916 );
   not U9185 ( n8916,n7314 );
   nor U9186 ( n7314,n6527,n6083 );
   nand U9187 ( n9378,n8106,n9379 );
   nor U9188 ( n8106,n6541,n6086 );
   nor U9189 ( n9376,n8915,n7276 );
   not U9190 ( n7276,n7229 );
   nor U9191 ( n7229,n6555,n6089 );
   nand U9192 ( n8915,n9380,n9379 );
   not U9193 ( n9379,n7315 );
   nor U9194 ( n7315,n7302,n6538 );
   nand U9195 ( n9380,n6541,n6086 );
   nor U9196 ( n9360,n7957,n8057 );
   nand U9197 ( n8057,n7879,n6314 );
   nor U9198 ( n7957,n6300,n7905 );
   nand U9199 ( n8946,n9381,n6653 );
   nor U9200 ( n9381,n8951,n9382 );
   and U9201 ( n8951,n9383,n9384 );
   nor U9202 ( n9384,n9385,n9386 );
   nand U9203 ( n9386,n9387,n9388 );
   nor U9204 ( n9388,n9389,n9390 );
   or U9205 ( n9390,n7628,n7650 );
   nor U9206 ( n7650,n7689,n9391 );
   not U9207 ( n9391,n7692 );
   nand U9208 ( n7692,n6398,n6387 );
   nor U9209 ( n7689,n6387,n6398 );
   and U9210 ( n7628,n7727,n7729 );
   nand U9211 ( n7729,n7614,n6056 );
   nand U9212 ( n7727,n6401,n6412 );
   nand U9213 ( n9389,n7693,n7720 );
   nand U9214 ( n7720,n8133,n9392 );
   nand U9215 ( n9392,n7706,n6047 );
   nand U9216 ( n8133,n6370,n6359 );
   not U9217 ( n6370,n6047 );
   nand U9218 ( n7693,n8135,n8137 );
   nand U9219 ( n8137,n6384,n6373 );
   not U9220 ( n8135,n7687 );
   nor U9221 ( n7687,n6373,n6384 );
   nor U9222 ( n9387,n9393,n9394 );
   nand U9223 ( n9394,n7464,n7487 );
   nand U9224 ( n7487,n8154,n9395 );
   nand U9225 ( n9395,n7473,n6068 );
   nand U9226 ( n8154,n6468,n6457 );
   nand U9227 ( n7464,n8160,n8157 );
   not U9228 ( n8157,n7453 );
   nor U9229 ( n7453,n6471,n6482 );
   nand U9230 ( n8160,n6482,n6471 );
   nand U9231 ( n9393,n7559,n7591 );
   nand U9232 ( n7591,n8144,n8146 );
   nand U9233 ( n8146,n7582,n6059 );
   nand U9234 ( n8144,n6426,n6415 );
   nand U9235 ( n7559,n7600,n7599 );
   nand U9236 ( n7599,n6429,n6440 );
   not U9237 ( n7600,n7605 );
   nor U9238 ( n7605,n6429,n6440 );
   nand U9239 ( n9385,n9396,n9397 );
   nor U9240 ( n9397,n9398,n9399 );
   nand U9241 ( n9399,n7954,n8045 );
   not U9242 ( n8045,n8013 );
   nor U9243 ( n8013,n6690,n6689 );
   nor U9244 ( n6689,n6026,n8011 );
   not U9245 ( n8011,n6261 );
   nor U9246 ( n6690,n6261,n6272 );
   nand U9247 ( n7954,n8196,n7943 );
   nand U9248 ( n7943,n7905,n6032 );
   nand U9249 ( n8196,n6300,n6289 );
   nand U9250 ( n9398,n9400,n7987 );
   not U9251 ( n7987,n7965 );
   nor U9252 ( n7965,n8016,n8124 );
   nor U9253 ( n8124,n6029,n7972 );
   nor U9254 ( n8016,n6275,n6286 );
   not U9255 ( n6286,n6029 );
   nor U9256 ( n9400,n8944,n7055 );
   and U9257 ( n7055,n8185,n8187 );
   nand U9258 ( n8187,n6636,n6625 );
   nand U9259 ( n8185,n7032,n6104 );
   nor U9260 ( n8944,n6219,n8227 );
   nor U9261 ( n9396,n9401,n9402 );
   nand U9262 ( n9402,n7760,n7782 );
   nand U9263 ( n7782,n8019,n8021 );
   nand U9264 ( n8021,n7789,n6041 );
   nand U9265 ( n8019,n6342,n6331 );
   nand U9266 ( n7760,n8025,n8022 );
   nand U9267 ( n8022,n6356,n6345 );
   nand U9268 ( n8025,n7740,n6044 );
   nand U9269 ( n9401,n7846,n7887 );
   nand U9270 ( n7887,n7915,n7911 );
   nand U9271 ( n7911,n6314,n6303 );
   not U9272 ( n7915,n7939 );
   nor U9273 ( n7939,n6303,n6314 );
   not U9274 ( n7846,n7860 );
   nor U9275 ( n7860,n7948,n7917 );
   nor U9276 ( n7917,n6317,n6328 );
   nor U9277 ( n7948,n6038,n7844 );
   nor U9278 ( n9383,n9403,n9404 );
   nand U9279 ( n9404,n9405,n9406 );
   nor U9280 ( n9406,n9407,n9408 );
   nand U9281 ( n9408,n9409,n6651 );
   nand U9282 ( n6651,n9153,n7020 );
   not U9283 ( n7020,n8190 );
   nor U9284 ( n8190,n6647,n9290 );
   nand U9285 ( n9153,n9290,n6647 );
   nand U9286 ( n9409,n6727,n6229 );
   not U9287 ( n6229,n8207 );
   not U9288 ( n6727,n6020 );
   nand U9289 ( n9407,n7021,n7090 );
   nand U9290 ( n7090,n8184,n8182 );
   nand U9291 ( n8182,n7079,n6101 );
   nand U9292 ( n8184,n6622,n6611 );
   nand U9293 ( n7021,n8189,n8191 );
   nand U9294 ( n8191,n6650,n6639 );
   nand U9295 ( n8189,n7011,n6107 );
   nor U9296 ( n9405,n9410,n9411 );
   nand U9297 ( n9411,n7388,n9412 );
   not U9298 ( n9412,n9359 );
   nand U9299 ( n9359,n8854,n8929 );
   nand U9300 ( n8929,n8207,n6020 );
   nand U9301 ( n6020,n9413,n9414 );
   nand U9302 ( n9414,reg2_reg_30_,n9415 );
   nor U9303 ( n9413,n9416,n9417 );
   nor U9304 ( n9417,n5958,n9418 );
   not U9305 ( n9418,reg0_reg_30_ );
   nor U9306 ( n9416,n5953,n9419 );
   not U9307 ( n9419,reg1_reg_30_ );
   nand U9308 ( n8207,datai_30_,n5962 );
   nand U9309 ( n8854,n8227,n6219 );
   not U9310 ( n6219,n8212 );
   nand U9311 ( n8212,datai_31_,n5962 );
   not U9312 ( n8227,n6017 );
   nand U9313 ( n6017,n9420,n9421 );
   nand U9314 ( n9421,reg2_reg_31_,n9415 );
   nor U9315 ( n9420,n9422,n9423 );
   nor U9316 ( n9423,n5959,n9424 );
   not U9317 ( n9424,reg0_reg_31_ );
   nor U9318 ( n9422,n5954,n9425 );
   not U9319 ( n9425,reg1_reg_31_ );
   xor U9320 ( n7388,n6077,n6499 );
   nand U9321 ( n9410,n7533,n6687 );
   nor U9322 ( n6687,n8945,n8936 );
   nor U9323 ( n8936,n6694,n6257 );
   not U9324 ( n6257,n6023 );
   not U9325 ( n6694,n6244 );
   nor U9326 ( n8945,n6023,n6244 );
   nand U9327 ( n6244,datai_29_,n5962 );
   xor U9328 ( n7533,n6454,n7509 );
   nand U9329 ( n9403,n9426,n9427 );
   nor U9330 ( n9427,n9428,n9429 );
   or U9331 ( n9429,n7272,n7316 );
   nor U9332 ( n7316,n7355,n9430 );
   not U9333 ( n9430,n7354 );
   nand U9334 ( n7354,n6538,n6527 );
   nor U9335 ( n7355,n6527,n6538 );
   nor U9336 ( n7272,n7364,n7368 );
   nor U9337 ( n7368,n6541,n6552 );
   nor U9338 ( n7364,n6086,n7256 );
   or U9339 ( n9428,n7348,n7425 );
   and U9340 ( n7425,n8161,n7458 );
   nand U9341 ( n7458,n6496,n6485 );
   not U9342 ( n8161,n7455 );
   nor U9343 ( n7455,n6485,n6496 );
   nor U9344 ( n7348,n7359,n9431 );
   not U9345 ( n9431,n8169 );
   nand U9346 ( n8169,n6524,n6513 );
   nor U9347 ( n7359,n6513,n6524 );
   not U9348 ( n6524,n6080 );
   nor U9349 ( n9426,n9432,n9433 );
   nand U9350 ( n9433,n7123,n7155 );
   not U9351 ( n7155,n7162 );
   nor U9352 ( n7162,n7165,n8194 );
   nor U9353 ( n8194,n6095,n7141 );
   nor U9354 ( n7165,n6583,n6594 );
   nand U9355 ( n7123,n8195,n7160 );
   nand U9356 ( n7160,n6608,n6597 );
   not U9357 ( n8195,n7161 );
   nor U9358 ( n7161,n6597,n6608 );
   nand U9359 ( n9432,n7195,n7230 );
   nand U9360 ( n7230,n7367,n8177 );
   nand U9361 ( n8177,n7216,n6089 );
   nand U9362 ( n7367,n6566,n6555 );
   not U9363 ( n6566,n6089 );
   not U9364 ( n7195,n7200 );
   nor U9365 ( n7200,n7242,n7246 );
   nor U9366 ( n7246,n6092,n7175 );
   nor U9367 ( n7242,n6569,n6580 );
   nand U9368 ( n8827,b_reg,n9434 );
   nand U9369 ( n9434,n9435,n9436 );
   nor U9370 ( n9436,n9437,n9438 );
   nor U9371 ( n9438,n9160,n9270 );
   nor U9372 ( n9437,n9439,n8812 );
   nor U9373 ( n9439,n9440,n9441 );
   nand U9374 ( n9441,n8732,n8823 );
   nand U9375 ( n9440,n6667,n8734 );
   nor U9376 ( n9435,n5973,n8826 );
   nor U9377 ( n9443,n9444,n9445 );
   nand U9378 ( n9445,n9446,n9447 );
   or U9379 ( n9447,n9448,n9449 );
   xor U9380 ( n9448,n9450,n9451 );
   xor U9381 ( n9451,n9452,n9453 );
   nand U9382 ( n9446,n9454,n6068 );
   nor U9383 ( n9444,n6443,n9455 );
   nor U9384 ( n9442,n9456,n9457 );
   nand U9385 ( n9457,n9458,n9459 );
   nand U9386 ( n9459,n7508,n9460 );
   nand U9387 ( n9458,n9461,n6062 );
   nor U9388 ( n9456,state_reg,n9462 );
   nor U9389 ( n9464,n9465,n9466 );
   nand U9390 ( n9466,n9467,n9468 );
   nand U9391 ( n9468,n9469,n5984 );
   nor U9392 ( n9469,n9471,n9472 );
   nor U9393 ( n9472,n9473,n9474 );
   nand U9394 ( n9474,n9475,n9476 );
   nand U9395 ( n9475,n9477,n9478 );
   nand U9396 ( n9477,n9479,n9480 );
   nor U9397 ( n9473,n9481,n9482 );
   nor U9398 ( n9471,n9483,n9484 );
   nand U9399 ( n9484,n9485,n9486 );
   nand U9400 ( n9485,n9487,n9476 );
   not U9401 ( n9483,n9488 );
   nand U9402 ( n9467,n9461,n6029 );
   nor U9403 ( n9465,n6314,n9489 );
   nor U9404 ( n9463,n9490,n9491 );
   nand U9405 ( n9491,n9492,n9493 );
   nand U9406 ( n9493,n9494,n7905 );
   nand U9407 ( n9492,n7923,n9495 );
   not U9408 ( n7923,n9496 );
   and U9409 ( n9490,n5973,reg3_reg_26_ );
   nor U9410 ( n9498,n9499,n9500 );
   nand U9411 ( n9500,n9501,n9502 );
   nand U9412 ( n9502,n9503,n5984 );
   nor U9413 ( n9503,n9504,n9505 );
   nor U9414 ( n9505,n9506,n9507 );
   nand U9415 ( n9507,n9508,n9509 );
   nor U9416 ( n9504,n9510,n9511 );
   xor U9417 ( n9511,n9512,n9513 );
   nand U9418 ( n9501,n9494,n7175 );
   nor U9419 ( n9499,n6594,n9489 );
   nor U9420 ( n9497,n9514,n9515 );
   nand U9421 ( n9515,n9516,n9517 );
   nand U9422 ( n9517,n5993,n6089 );
   nand U9423 ( n9516,n7181,n9460 );
   and U9424 ( n9514,n5932,reg3_reg_6_ );
   nor U9425 ( n9519,n9520,n9521 );
   nand U9426 ( n9521,n9522,n9523 );
   or U9427 ( n9523,n9524,n9449 );
   xor U9428 ( n9524,n9525,n9526 );
   xor U9429 ( n9525,n9527,n9528 );
   nand U9430 ( n9522,n9494,n7614 );
   nor U9431 ( n9520,n9529,n7621 );
   nor U9432 ( n9518,n9530,n9531 );
   nand U9433 ( n9531,n9532,n9533 );
   nand U9434 ( n9533,n9454,n6059 );
   nand U9435 ( n9532,n5993,n6053 );
   nor U9436 ( n9530,state_reg,n9534 );
   nor U9437 ( n9536,n9537,n9538 );
   nand U9438 ( n9538,n9539,n9540 );
   nand U9439 ( n9540,n9470,n9541 );
   nand U9440 ( n9541,n9542,n9543 );
   nand U9441 ( n9543,n9544,n9545 );
   nor U9442 ( n9542,n9546,n9547 );
   nor U9443 ( n9547,n9548,n9549 );
   xor U9444 ( n9549,n9550,n9545 );
   not U9445 ( n9548,n9551 );
   nor U9446 ( n9546,n9551,n9552 );
   nand U9447 ( n9552,n9553,n9550 );
   nand U9448 ( n9539,reg3_reg_2_,n9554 );
   nor U9449 ( n9537,n6650,n9489 );
   nor U9450 ( n9535,n9555,n9556 );
   nor U9451 ( n9556,n6622,n9557 );
   nor U9452 ( n9555,n6625,n9455 );
   nor U9453 ( n9559,n9560,n9561 );
   nand U9454 ( n9561,n9562,n9563 );
   nand U9455 ( n9563,n9564,n9470 );
   nor U9456 ( n9564,n9565,n9566 );
   nor U9457 ( n9566,n9567,n9568 );
   xor U9458 ( n9568,n9569,n9570 );
   nor U9459 ( n9565,n9571,n9572 );
   nor U9460 ( n9572,n9573,n9574 );
   nand U9461 ( n9562,n5983,n6080 );
   nor U9462 ( n9560,n6499,n5985 );
   nor U9463 ( n9558,n9575,n9576 );
   nand U9464 ( n9576,n9577,n9578 );
   nand U9465 ( n9578,n7380,n9460 );
   nand U9466 ( n9577,n5993,n6074 );
   nor U9467 ( n9575,state_reg,n9579 );
   nor U9468 ( n9581,n9582,n9583 );
   nand U9469 ( n9583,n9584,n9585 );
   nand U9470 ( n9585,n9470,n9586 );
   xor U9471 ( n9586,n9587,n9588 );
   xor U9472 ( n9588,n9589,n9590 );
   nand U9473 ( n9584,n9494,n7740 );
   nor U9474 ( n9582,n9591,n7746 );
   nor U9475 ( n9580,n9592,n9593 );
   nand U9476 ( n9593,n9594,n9595 );
   nand U9477 ( n9595,n5983,n6047 );
   nand U9478 ( n9594,n5993,n6041 );
   nor U9479 ( n9592,state_reg,n9596 );
   nor U9480 ( n9598,n9599,n9600 );
   nand U9481 ( n9600,n9601,n9602 );
   nand U9482 ( n9602,n9603,n9470 );
   nor U9483 ( n9603,n9604,n9605 );
   nor U9484 ( n9605,n9606,n9607 );
   nand U9485 ( n9607,n9608,n9609 );
   nand U9486 ( n9608,n9610,n9611 );
   nor U9487 ( n9606,n9612,n9613 );
   nor U9488 ( n9604,n9614,n9615 );
   nand U9489 ( n9615,n9616,n9617 );
   nand U9490 ( n9616,n9618,n9609 );
   nand U9491 ( n9601,n5993,n6068 );
   nor U9492 ( n9599,n6496,n9489 );
   nor U9493 ( n9597,n9619,n9620 );
   nand U9494 ( n9620,n9621,n9622 );
   nand U9495 ( n9622,n9494,n7442 );
   nand U9496 ( n9621,n7441,n9460 );
   nor U9497 ( n9619,state_reg,n9623 );
   nor U9498 ( n9625,n9626,n9627 );
   nand U9499 ( n9627,n9628,n9629 );
   nand U9500 ( n9629,n9470,n9630 );
   nand U9501 ( n9630,n9631,n9632 );
   nand U9502 ( n9632,n9633,n9634 );
   nor U9503 ( n9631,n9635,n9636 );
   nor U9504 ( n9636,n9637,n9638 );
   xor U9505 ( n9638,n9634,n9639 );
   nor U9506 ( n9635,n9640,n9641 );
   nand U9507 ( n9641,n9642,n9639 );
   nand U9508 ( n9628,n5983,n6053 );
   nor U9509 ( n9626,n6373,n9455 );
   nor U9510 ( n9624,n9643,n9644 );
   nand U9511 ( n9644,n9645,n9646 );
   nand U9512 ( n9646,n7669,n9495 );
   not U9513 ( n7669,n9647 );
   nand U9514 ( n9645,n9461,n6047 );
   nor U9515 ( n9643,state_reg,n9648 );
   nor U9516 ( n9650,n9651,n9652 );
   nor U9517 ( n9652,n8733,n9449 );
   xor U9518 ( n8733,n9653,n9654 );
   xor U9519 ( n9653,n9655,n6008 );
   and U9520 ( n9651,n9554,reg3_reg_0_ );
   nor U9521 ( n9649,n9656,n9657 );
   nor U9522 ( n9657,n6650,n9557 );
   nor U9523 ( n9656,n6647,n9455 );
   nor U9524 ( n9659,n9660,n9661 );
   nand U9525 ( n9661,n9662,n9663 );
   or U9526 ( n9663,n9664,n9449 );
   xor U9527 ( n9664,n9665,n9666 );
   xor U9528 ( n9665,n9667,n9668 );
   nand U9529 ( n9662,n9494,n7302 );
   nor U9530 ( n9660,n9529,n7301 );
   nor U9531 ( n9658,n9669,n9670 );
   nand U9532 ( n9670,n9671,n9672 );
   nand U9533 ( n9672,n9461,n6080 );
   nand U9534 ( n9671,n9454,n6086 );
   and U9535 ( n9669,n5975,reg3_reg_9_ );
   nor U9536 ( n9674,n9675,n9676 );
   nand U9537 ( n9676,n9677,n9678 );
   nand U9538 ( n9678,n9679,n9470 );
   xor U9539 ( n9679,n9680,n9681 );
   xor U9540 ( n9680,n9682,n9683 );
   nand U9541 ( n9677,n9454,n6101 );
   nor U9542 ( n9675,n6597,n5985 );
   nor U9543 ( n9673,n8667,n9684 );
   nand U9544 ( n9684,n9685,n9686 );
   nand U9545 ( n9686,n7113,n9460 );
   not U9546 ( n7113,n9687 );
   nand U9547 ( n9685,n9461,n6095 );
   nor U9548 ( n8667,state_reg,n9688 );
   nor U9549 ( n9690,n9691,n9692 );
   nand U9550 ( n9692,n9693,n9694 );
   nand U9551 ( n9694,n9470,n9695 );
   xor U9552 ( n9695,n9696,n9697 );
   nand U9553 ( n9696,n9698,n9699 );
   nand U9554 ( n9693,n9461,n6035 );
   nor U9555 ( n9691,n6342,n9489 );
   nor U9556 ( n9689,n9700,n9701 );
   nand U9557 ( n9701,n9702,n9703 );
   nand U9558 ( n9703,n9494,n7844 );
   nand U9559 ( n9702,n7852,n9495 );
   not U9560 ( n7852,n9704 );
   nor U9561 ( n9700,state_reg,n9705 );
   nor U9562 ( n9707,n9708,n9709 );
   nand U9563 ( n9709,n9710,n9711 );
   nand U9564 ( n9711,n9712,n9470 );
   nor U9565 ( n9712,n9713,n9714 );
   nor U9566 ( n9714,n9715,n9716 );
   nor U9567 ( n9715,n9717,n9718 );
   nor U9568 ( n9713,n9719,n9720 );
   nand U9569 ( n9720,n9721,n9722 );
   nand U9570 ( n9721,n9723,n9724 );
   or U9571 ( n9719,n9718,n9717 );
   nand U9572 ( n9710,n9461,n6056 );
   nor U9573 ( n9708,n6440,n9489 );
   nor U9574 ( n9706,n9725,n9726 );
   nand U9575 ( n9726,n9727,n9728 );
   nand U9576 ( n9728,n9494,n7582 );
   nand U9577 ( n9727,n7581,n9460 );
   nor U9578 ( n9725,state_reg,n9729 );
   nor U9579 ( n9731,n9732,n9733 );
   nand U9580 ( n9733,n9734,n9735 );
   nand U9581 ( n9735,n9736,n9470 );
   xor U9582 ( n9736,n9737,n9738 );
   xor U9583 ( n9738,n9739,n9740 );
   nand U9584 ( n9734,n9454,n6098 );
   nor U9585 ( n9732,n6583,n5985 );
   nor U9586 ( n9730,n9741,n9742 );
   nand U9587 ( n9742,n9743,n9744 );
   nand U9588 ( n9744,n7140,n9460 );
   nand U9589 ( n9743,n9461,n6092 );
   nor U9590 ( n9741,state_reg,n9745 );
   nor U9591 ( n9747,n9748,n9749 );
   nand U9592 ( n9749,n9750,n9751 );
   nand U9593 ( n9751,n9470,n9752 );
   nand U9594 ( n9752,n9753,n9754 );
   nand U9595 ( n9754,n9755,n9756 );
   nor U9596 ( n9753,n9757,n9758 );
   nor U9597 ( n9758,n9759,n9760 );
   xor U9598 ( n9760,n9761,n9756 );
   not U9599 ( n9759,n9762 );
   nor U9600 ( n9757,n9762,n9763 );
   nand U9601 ( n9763,n9724,n9761 );
   nand U9602 ( n9750,n9454,n6065 );
   nor U9603 ( n9748,n6429,n9455 );
   nor U9604 ( n9746,n9764,n9765 );
   nand U9605 ( n9765,n9766,n9767 );
   nand U9606 ( n9767,n7549,n9460 );
   not U9607 ( n7549,n9768 );
   nand U9608 ( n9766,n9461,n6059 );
   nor U9609 ( n9764,state_reg,n9769 );
   nor U9610 ( n9771,n9772,n9773 );
   nand U9611 ( n9773,n9774,n9775 );
   nand U9612 ( n9775,n9470,n9776 );
   nand U9613 ( n9776,n9777,n9778 );
   nand U9614 ( n9778,n9779,n9478 );
   nor U9615 ( n9777,n9780,n9781 );
   nor U9616 ( n9781,n9782,n9783 );
   xor U9617 ( n9783,n9478,n9480 );
   nor U9618 ( n9780,n9479,n9784 );
   nand U9619 ( n9784,n9487,n9480 );
   not U9620 ( n9487,n9478 );
   nand U9621 ( n9774,n9494,n7879 );
   nor U9622 ( n9772,n9591,n7878 );
   not U9623 ( n9591,n9495 );
   nor U9624 ( n9770,n9785,n9786 );
   nand U9625 ( n9786,n9787,n9788 );
   nand U9626 ( n9788,n9454,n6038 );
   nand U9627 ( n9787,n9461,n6032 );
   nor U9628 ( n9785,state_reg,n9789 );
   nor U9629 ( n9791,n9792,n9793 );
   nand U9630 ( n9793,n9794,n9795 );
   nand U9631 ( n9795,n9796,n9470 );
   nor U9632 ( n9796,n9797,n9798 );
   nor U9633 ( n9798,n9610,n9799 );
   xor U9634 ( n9799,n9800,n9801 );
   not U9635 ( n9610,n9618 );
   nor U9636 ( n9797,n9618,n9802 );
   nand U9637 ( n9802,n9611,n9609 );
   nor U9638 ( n9618,n9573,n9803 );
   and U9639 ( n9803,n9571,n9804 );
   nand U9640 ( n9804,n9570,n9805 );
   not U9641 ( n9571,n9567 );
   nand U9642 ( n9567,n9806,n9807 );
   nand U9643 ( n9807,n9808,n9809 );
   nand U9644 ( n9794,n9454,n6077 );
   nor U9645 ( n9792,n6485,n9455 );
   nor U9646 ( n9790,n9810,n9811 );
   nand U9647 ( n9811,n9812,n9813 );
   nand U9648 ( n9813,n7417,n9460 );
   not U9649 ( n7417,n9814 );
   nand U9650 ( n9812,n9461,n6071 );
   nor U9651 ( n9810,state_reg,n9815 );
   nor U9652 ( n9817,n9818,n9819 );
   nand U9653 ( n9819,n9820,n9821 );
   nand U9654 ( n9821,n9822,n5984 );
   nor U9655 ( n9822,n9823,n9824 );
   nor U9656 ( n9824,n9825,n9826 );
   nand U9657 ( n9826,n9827,n9828 );
   nand U9658 ( n9827,n9829,n9634 );
   nor U9659 ( n9825,n9830,n9831 );
   nor U9660 ( n9823,n9832,n9833 );
   nand U9661 ( n9833,n9834,n9835 );
   nand U9662 ( n9834,n9642,n9828 );
   not U9663 ( n9828,n9633 );
   not U9664 ( n9642,n9634 );
   nand U9665 ( n9634,n9836,n9837 );
   nand U9666 ( n9820,n9461,n6044 );
   nor U9667 ( n9818,n6384,n9489 );
   nor U9668 ( n9816,n9838,n9839 );
   nand U9669 ( n9839,n9840,n9841 );
   nand U9670 ( n9841,n9494,n7706 );
   nand U9671 ( n9840,n7705,n9495 );
   nor U9672 ( n9838,state_reg,n9842 );
   nor U9673 ( n9844,n9845,n9846 );
   nand U9674 ( n9846,n9847,n9848 );
   nand U9675 ( n9848,n9470,n9849 );
   xor U9676 ( n9849,n9850,n9851 );
   nand U9677 ( n9850,n9852,n9853 );
   nand U9678 ( n9847,reg3_reg_1_,n9554 );
   nand U9679 ( n9554,n9529,state_reg );
   nor U9680 ( n9845,n9290,n9489 );
   nor U9681 ( n9843,n9854,n9855 );
   nor U9682 ( n9855,n6636,n9557 );
   nor U9683 ( n9854,n6639,n9455 );
   nor U9684 ( n9857,n9858,n9859 );
   nand U9685 ( n9859,n9860,n9861 );
   nand U9686 ( n9861,n9862,n9470 );
   xor U9687 ( n9862,n9863,n9864 );
   nand U9688 ( n9864,n9865,n9866 );
   nand U9689 ( n9860,n9461,n6083 );
   nor U9690 ( n9858,n6541,n9455 );
   nor U9691 ( n9856,n9867,n9868 );
   nand U9692 ( n9868,n9869,n9870 );
   nand U9693 ( n9870,n9454,n6089 );
   nand U9694 ( n9869,n7262,n9460 );
   not U9695 ( n7262,n9871 );
   nor U9696 ( n9867,state_reg,n9872 );
   nor U9697 ( n9874,n9875,n9876 );
   nand U9698 ( n9876,n9877,n9878 );
   nand U9699 ( n9878,n9879,n9470 );
   xor U9700 ( n9879,n9880,n9881 );
   xor U9701 ( n9881,n9882,n9883 );
   nand U9702 ( n9883,n9884,n9885 );
   not U9703 ( n9885,n9886 );
   nor U9704 ( n9882,n9887,n9888 );
   nor U9705 ( n9888,n6272,n9889 );
   nor U9706 ( n9887,n6261,n9890 );
   xor U9707 ( n9880,n6011,n9891 );
   nor U9708 ( n9891,n9892,n9893 );
   nor U9709 ( n9893,n6272,n5982 );
   nor U9710 ( n9892,n5991,n6261 );
   nand U9711 ( n9877,n9461,n6023 );
   nand U9712 ( n6023,n9895,n9896 );
   nor U9713 ( n9896,n9897,n9898 );
   nor U9714 ( n9898,n5956,n9899 );
   not U9715 ( n9899,reg1_reg_29_ );
   nor U9716 ( n9897,n6004,n6684 );
   nand U9717 ( n6684,n9900,reg3_reg_28_ );
   nor U9718 ( n9895,n9901,n9902 );
   and U9719 ( n9902,n9415,reg2_reg_29_ );
   nor U9720 ( n9901,n5961,n9903 );
   not U9721 ( n9903,reg0_reg_29_ );
   nor U9722 ( n9875,n6261,n9455 );
   nand U9723 ( n6261,datai_28_,n5962 );
   nor U9724 ( n9873,n9904,n9905 );
   nand U9725 ( n9905,n9906,n9907 );
   nand U9726 ( n9907,n9454,n6029 );
   nand U9727 ( n9906,n8034,n9495 );
   and U9728 ( n9904,n5932,reg3_reg_28_ );
   nor U9729 ( n9909,n9910,n9911 );
   nand U9730 ( n9911,n9912,n9913 );
   nand U9731 ( n9913,n9470,n9914 );
   nand U9732 ( n9914,n9915,n9916 );
   nand U9733 ( n9916,n9917,n9918 );
   nor U9734 ( n9915,n9919,n9920 );
   nor U9735 ( n9920,n9921,n9922 );
   xor U9736 ( n9922,n9923,n9917 );
   nor U9737 ( n9919,n9924,n9925 );
   nand U9738 ( n9925,n9923,n9926 );
   nand U9739 ( n9912,n9454,n6056 );
   nor U9740 ( n9910,n6387,n9455 );
   nor U9741 ( n9908,n8267,n9927 );
   nand U9742 ( n9927,n9928,n9929 );
   nand U9743 ( n9929,n7642,n9460 );
   nand U9744 ( n9928,n9461,n6050 );
   nor U9745 ( n8267,state_reg,n9930 );
   nor U9746 ( n9932,n9933,n9934 );
   nand U9747 ( n9934,n9935,n9936 );
   nand U9748 ( n9936,n9937,n9470 );
   nor U9749 ( n9937,n9938,n9939 );
   nor U9750 ( n9939,n9940,n9941 );
   nor U9751 ( n9940,n9942,n9943 );
   nor U9752 ( n9938,n9944,n9945 );
   nand U9753 ( n9945,n9946,n9947 );
   nand U9754 ( n9946,n9553,n9948 );
   not U9755 ( n9553,n9545 );
   or U9756 ( n9944,n9943,n9942 );
   nand U9757 ( n9935,n9454,n6104 );
   nor U9758 ( n9933,n6611,n9455 );
   nor U9759 ( n9931,n9949,n9950 );
   nand U9760 ( n9950,n9951,n8694 );
   nand U9761 ( n8694,reg3_reg_3_,n5973 );
   nand U9762 ( n9951,n9460,n7078 );
   nor U9763 ( n9949,n6608,n9557 );
   nor U9764 ( n9953,n9954,n9955 );
   nand U9765 ( n9955,n9956,n9957 );
   nand U9766 ( n9957,n9470,n9958 );
   xor U9767 ( n9958,n9959,n9808 );
   nand U9768 ( n9959,n9809,n9806 );
   not U9769 ( n9806,n9960 );
   nand U9770 ( n9956,n9454,n6083 );
   nor U9771 ( n9954,n6513,n9455 );
   nor U9772 ( n9952,n9961,n9962 );
   nand U9773 ( n9962,n9963,n9964 );
   nand U9774 ( n9964,n7334,n9460 );
   not U9775 ( n7334,n9965 );
   nand U9776 ( n9963,n9461,n6077 );
   nor U9777 ( n9961,state_reg,n9966 );
   nor U9778 ( n9968,n9969,n9970 );
   nand U9779 ( n9970,n9971,n9972 );
   or U9780 ( n9972,n9973,n9449 );
   xor U9781 ( n9973,n9974,n9975 );
   xor U9782 ( n9975,n9976,n9977 );
   nand U9783 ( n9971,n9454,n6044 );
   nor U9784 ( n9969,n6331,n9455 );
   nor U9785 ( n9967,n9978,n9979 );
   nand U9786 ( n9979,n9980,n9981 );
   nand U9787 ( n9981,n7788,n9495 );
   nand U9788 ( n9980,n9461,n6038 );
   nor U9789 ( n9978,state_reg,n9982 );
   nor U9790 ( n9984,n9985,n9986 );
   nand U9791 ( n9986,n9987,n9988 );
   or U9792 ( n9988,n9449,n9989 );
   xor U9793 ( n9989,n9990,n9991 );
   xor U9794 ( n9990,n9992,n9993 );
   nand U9795 ( n9987,n9494,n7473 );
   nor U9796 ( n9985,n9529,n7479 );
   not U9797 ( n9529,n9460 );
   nor U9798 ( n9983,n9994,n9995 );
   nand U9799 ( n9995,n9996,n9997 );
   nand U9800 ( n9997,n9454,n6071 );
   nand U9801 ( n9996,n5993,n6065 );
   not U9802 ( n9461,n9557 );
   nor U9803 ( n9994,state_reg,n9998 );
   nor U9804 ( n10000,n10001,n10002 );
   nand U9805 ( n10002,n10003,n10004 );
   nand U9806 ( n10004,n9470,n10005 );
   nand U9807 ( n10005,n10006,n10007 );
   nand U9808 ( n10007,n10008,n10009 );
   nand U9809 ( n10008,n9884,n10010 );
   nand U9810 ( n10006,n9886,n9884 );
   nand U9811 ( n9884,n10011,n10012 );
   not U9812 ( n10012,n10013 );
   xor U9813 ( n10011,n10014,n10015 );
   nor U9814 ( n9886,n10009,n10016 );
   not U9815 ( n10016,n10010 );
   nand U9816 ( n10010,n10017,n10013 );
   nand U9817 ( n10013,n10018,n10019 );
   nand U9818 ( n10019,n5996,n6029 );
   nand U9819 ( n10018,n5940,n7972 );
   xor U9820 ( n10017,n6008,n10014 );
   and U9821 ( n10014,n10022,n10023 );
   nand U9822 ( n10023,n5940,n6029 );
   nand U9823 ( n6029,n10024,n10025 );
   nor U9824 ( n10025,n10026,n10027 );
   nor U9825 ( n10027,n5956,n10028 );
   not U9826 ( n10028,reg1_reg_27_ );
   nor U9827 ( n10026,n10029,n6005 );
   not U9828 ( n10029,n7971 );
   nor U9829 ( n10024,n10030,n10031 );
   and U9830 ( n10031,n9415,reg2_reg_27_ );
   nor U9831 ( n10030,n5961,n10032 );
   not U9832 ( n10032,reg0_reg_27_ );
   nand U9833 ( n10022,n7972,n10033 );
   nand U9834 ( n10009,n10034,n10035 );
   nand U9835 ( n10035,n9488,n9478 );
   nand U9836 ( n9478,n9698,n10036 );
   nand U9837 ( n10036,n10037,n9699 );
   or U9838 ( n9699,n10038,n10039 );
   not U9839 ( n10037,n9697 );
   nand U9840 ( n9697,n10040,n10041 );
   nand U9841 ( n10041,n9974,n10042 );
   nand U9842 ( n10042,n9976,n9977 );
   xor U9843 ( n9974,n10043,n10015 );
   nor U9844 ( n10043,n10044,n10045 );
   nor U9845 ( n10045,n6342,n9890 );
   not U9846 ( n6342,n6041 );
   nor U9847 ( n10044,n5991,n6331 );
   or U9848 ( n10040,n9977,n9976 );
   and U9849 ( n9976,n10046,n10047 );
   nand U9850 ( n10047,n10048,n10049 );
   nand U9851 ( n10049,n9587,n9590 );
   not U9852 ( n10048,n9589 );
   nand U9853 ( n9589,n10050,n10051 );
   nand U9854 ( n10051,n10052,n10053 );
   nand U9855 ( n10052,n10054,n10055 );
   or U9856 ( n10055,n9837,n9832 );
   not U9857 ( n9837,n9918 );
   nor U9858 ( n9918,n9924,n9923 );
   nor U9859 ( n10054,n9633,n9831 );
   not U9860 ( n9831,n9835 );
   nand U9861 ( n9835,n10056,n10057 );
   nor U9862 ( n9633,n9640,n9639 );
   or U9863 ( n10050,n9836,n9832 );
   nand U9864 ( n9832,n10053,n9829 );
   nand U9865 ( n9829,n9639,n9640 );
   not U9866 ( n9640,n9637 );
   xor U9867 ( n9637,n10058,n6008 );
   nor U9868 ( n10058,n10059,n10060 );
   nor U9869 ( n10060,n6384,n9890 );
   not U9870 ( n6384,n6050 );
   nor U9871 ( n10059,n5990,n6373 );
   and U9872 ( n9639,n10061,n10062 );
   nand U9873 ( n10062,n5940,n7662 );
   not U9874 ( n7662,n6373 );
   nand U9875 ( n6373,datai_20_,n5962 );
   nand U9876 ( n10061,n10020,n6050 );
   nand U9877 ( n6050,n10063,n10064 );
   nor U9878 ( n10064,n10065,n10066 );
   nor U9879 ( n10066,n5953,n10067 );
   not U9880 ( n10067,reg1_reg_20_ );
   nor U9881 ( n10065,n6005,n9647 );
   nand U9882 ( n9647,n10068,n10069 );
   nand U9883 ( n10068,n9648,n10070 );
   or U9884 ( n10070,n9930,n10071 );
   not U9885 ( n9648,reg3_reg_20_ );
   nor U9886 ( n10063,n10072,n10073 );
   and U9887 ( n10073,n9415,reg2_reg_20_ );
   nor U9888 ( n10072,n5958,n10074 );
   not U9889 ( n10074,reg0_reg_20_ );
   not U9890 ( n10053,n9830 );
   nor U9891 ( n9830,n10056,n10057 );
   nand U9892 ( n10057,n10075,n10076 );
   nand U9893 ( n10076,n5940,n7706 );
   nand U9894 ( n10075,n5996,n6047 );
   xor U9895 ( n10056,n6010,n10077 );
   and U9896 ( n10077,n10078,n10079 );
   nand U9897 ( n10079,n7706,n10033 );
   not U9898 ( n7706,n6359 );
   nand U9899 ( n6359,datai_21_,n5962 );
   nand U9900 ( n10078,n5940,n6047 );
   nand U9901 ( n6047,n10080,n10081 );
   nor U9902 ( n10081,n10082,n10083 );
   nor U9903 ( n10083,n5953,n10084 );
   not U9904 ( n10084,reg1_reg_21_ );
   nor U9905 ( n10082,n10085,n6006 );
   not U9906 ( n10085,n7705 );
   xor U9907 ( n7705,n9842,n10069 );
   nor U9908 ( n10080,n10086,n10087 );
   and U9909 ( n10087,n9415,reg2_reg_21_ );
   nor U9910 ( n10086,n5958,n10088 );
   not U9911 ( n10088,reg0_reg_21_ );
   nand U9912 ( n9836,n9917,n10089 );
   nand U9913 ( n10089,n9923,n9924 );
   not U9914 ( n9924,n9921 );
   xor U9915 ( n9921,n10090,n6010 );
   nor U9916 ( n10090,n10091,n10092 );
   nor U9917 ( n10092,n6398,n5982 );
   not U9918 ( n6398,n6053 );
   nor U9919 ( n10091,n5990,n6387 );
   and U9920 ( n9923,n10093,n10094 );
   nand U9921 ( n10094,n5940,n7643 );
   not U9922 ( n7643,n6387 );
   nand U9923 ( n6387,n10095,n10096 );
   or U9924 ( n10096,n5964,datai_19_ );
   nand U9925 ( n10095,n8247,n5965 );
   nand U9926 ( n10093,n5996,n6053 );
   nand U9927 ( n6053,n10097,n10098 );
   nor U9928 ( n10098,n10099,n10100 );
   nor U9929 ( n10100,n5955,n8259 );
   not U9930 ( n8259,reg1_reg_19_ );
   nor U9931 ( n10099,n10101,n6004 );
   not U9932 ( n10101,n7642 );
   xor U9933 ( n7642,n9930,n10071 );
   nor U9934 ( n10097,n10102,n10103 );
   and U9935 ( n10103,n9415,reg2_reg_19_ );
   nor U9936 ( n10102,n5960,n10104 );
   not U9937 ( n10104,reg0_reg_19_ );
   not U9938 ( n9917,n9926 );
   nand U9939 ( n9926,n10105,n10106 );
   nand U9940 ( n10106,n10107,n9528 );
   nand U9941 ( n9528,n10108,n10109 );
   not U9942 ( n10109,n9717 );
   nor U9943 ( n9717,n10110,n10111 );
   or U9944 ( n10108,n9716,n9718 );
   and U9945 ( n9718,n10111,n10110 );
   nand U9946 ( n10110,n10112,n10113 );
   nand U9947 ( n10113,n5940,n7582 );
   not U9948 ( n7582,n6415 );
   nand U9949 ( n10112,n5996,n6059 );
   xor U9950 ( n10111,n10114,n6011 );
   nor U9951 ( n10114,n10115,n10116 );
   nor U9952 ( n10116,n6426,n5982 );
   not U9953 ( n6426,n6059 );
   nand U9954 ( n6059,n10117,n10118 );
   nor U9955 ( n10118,n10119,n10120 );
   nor U9956 ( n10120,n5955,n8297 );
   not U9957 ( n8297,reg1_reg_17_ );
   nor U9958 ( n10119,n10121,n6005 );
   not U9959 ( n10121,n7581 );
   xor U9960 ( n7581,n9729,n10122 );
   nor U9961 ( n10117,n10123,n10124 );
   nor U9962 ( n10124,n10125,n8290 );
   not U9963 ( n8290,reg2_reg_17_ );
   nor U9964 ( n10123,n5960,n10126 );
   not U9965 ( n10126,reg0_reg_17_ );
   nor U9966 ( n10115,n9894,n6415 );
   nand U9967 ( n6415,n10127,n10128 );
   or U9968 ( n10128,n5963,datai_17_ );
   nand U9969 ( n10127,n8292,n5966 );
   nand U9970 ( n8292,n10129,n10130 );
   nand U9971 ( n10130,n6860,n5987 );
   not U9972 ( n6860,ir_reg_17_ );
   nand U9973 ( n10129,ir_reg_31_,n6861 );
   nand U9974 ( n6861,n10132,n6867 );
   nand U9975 ( n10132,ir_reg_17_,n10133 );
   nand U9976 ( n9716,n9723,n10134 );
   nand U9977 ( n10134,n9756,n9722 );
   not U9978 ( n9722,n9755 );
   nor U9979 ( n9755,n9761,n9762 );
   not U9980 ( n9756,n9724 );
   nand U9981 ( n9724,n10135,n10136 );
   nand U9982 ( n10136,n9450,n10137 );
   nand U9983 ( n10137,n9453,n9452 );
   xor U9984 ( n9450,n10138,n10015 );
   nor U9985 ( n10138,n10139,n10140 );
   nor U9986 ( n10140,n6454,n5982 );
   not U9987 ( n6454,n6065 );
   nor U9988 ( n10139,n5991,n6443 );
   or U9989 ( n10135,n9452,n9453 );
   and U9990 ( n9453,n10141,n10142 );
   nand U9991 ( n10142,n9993,n10143 );
   nand U9992 ( n10143,n9991,n9992 );
   and U9993 ( n9993,n10144,n10145 );
   or U9994 ( n10145,n9609,n9612 );
   nand U9995 ( n9609,n9801,n9800 );
   nor U9996 ( n10144,n9613,n10146 );
   nor U9997 ( n10146,n10147,n9614 );
   nand U9998 ( n9614,n9611,n10148 );
   not U9999 ( n10148,n9612 );
   nor U10000 ( n9612,n10149,n10150 );
   or U10001 ( n9611,n9800,n9801 );
   xor U10002 ( n9801,n10151,n6010 );
   nor U10003 ( n10151,n10152,n10153 );
   nor U10004 ( n10153,n6496,n5982 );
   not U10005 ( n6496,n6074 );
   nor U10006 ( n10152,n5990,n6485 );
   nand U10007 ( n9800,n10154,n10155 );
   nand U10008 ( n10155,n5940,n7411 );
   not U10009 ( n7411,n6485 );
   nand U10010 ( n6485,n10156,n10157 );
   or U10011 ( n10157,n5963,datai_12_ );
   nand U10012 ( n10156,n5965,n8430 );
   nand U10013 ( n8430,n10158,n10159 );
   nor U10014 ( n10158,n10160,n10161 );
   nor U10015 ( n10161,n10131,n10162 );
   nand U10016 ( n10162,ir_reg_12_,n6822 );
   nor U10017 ( n10160,ir_reg_31_,ir_reg_12_ );
   nand U10018 ( n10154,n5996,n6074 );
   nand U10019 ( n6074,n10163,n10164 );
   nor U10020 ( n10164,n10165,n10166 );
   nor U10021 ( n10166,n5954,n8461 );
   not U10022 ( n8461,reg1_reg_12_ );
   nor U10023 ( n10165,n6006,n9814 );
   nand U10024 ( n9814,n10167,n10168 );
   nand U10025 ( n10167,n9815,n10169 );
   or U10026 ( n10169,n9579,n10170 );
   not U10027 ( n9815,reg3_reg_12_ );
   nor U10028 ( n10163,n10171,n10172 );
   nor U10029 ( n10172,n5995,n8436 );
   not U10030 ( n8436,reg2_reg_12_ );
   nor U10031 ( n10171,n5959,n10173 );
   not U10032 ( n10173,reg0_reg_12_ );
   nor U10033 ( n10147,n10174,n9573 );
   nor U10034 ( n9573,n9805,n9570 );
   not U10035 ( n9570,n10175 );
   not U10036 ( n9805,n9569 );
   nor U10037 ( n10174,n10176,n9574 );
   nor U10038 ( n9574,n9569,n10175 );
   nand U10039 ( n10175,n10177,n10178 );
   nand U10040 ( n10178,n5940,n7381 );
   not U10041 ( n7381,n6499 );
   nand U10042 ( n10177,n5996,n6077 );
   xor U10043 ( n9569,n10179,n6010 );
   nor U10044 ( n10179,n10180,n10181 );
   nor U10045 ( n10181,n6510,n9890 );
   not U10046 ( n6510,n6077 );
   nand U10047 ( n6077,n10182,n10183 );
   nor U10048 ( n10183,n10184,n10185 );
   nor U10049 ( n10185,n5954,n8465 );
   not U10050 ( n8465,reg1_reg_11_ );
   nor U10051 ( n10184,n10186,n6005 );
   not U10052 ( n10186,n7380 );
   xor U10053 ( n7380,n9579,n10170 );
   nor U10054 ( n10182,n10187,n10188 );
   nor U10055 ( n10188,n5995,n8457 );
   not U10056 ( n8457,reg2_reg_11_ );
   nor U10057 ( n10187,n5959,n10189 );
   not U10058 ( n10189,reg0_reg_11_ );
   nor U10059 ( n10180,n5990,n6499 );
   nand U10060 ( n6499,n10190,n10191 );
   or U10061 ( n10191,n5964,datai_11_ );
   nand U10062 ( n10190,n8459,n5964 );
   nand U10063 ( n8459,n10192,n10193 );
   nand U10064 ( n10193,n6815,n5987 );
   not U10065 ( n6815,ir_reg_11_ );
   nand U10066 ( n10192,ir_reg_31_,n6816 );
   nand U10067 ( n6816,n10194,n6822 );
   nand U10068 ( n10194,ir_reg_11_,n10195 );
   nor U10069 ( n10176,n10196,n10197 );
   not U10070 ( n10197,n9809 );
   nand U10071 ( n9809,n10198,n10199 );
   nor U10072 ( n10196,n9960,n9808 );
   nand U10073 ( n9808,n10200,n10201 );
   nand U10074 ( n10201,n10202,n9668 );
   nand U10075 ( n9668,n10203,n9865 );
   or U10076 ( n9865,n10204,n10205 );
   nand U10077 ( n10203,n9863,n9866 );
   nand U10078 ( n9866,n10205,n10204 );
   nand U10079 ( n10204,n10206,n10207 );
   nand U10080 ( n10207,n5940,n7256 );
   not U10081 ( n7256,n6541 );
   nand U10082 ( n10206,n5996,n6086 );
   xor U10083 ( n10205,n10208,n6010 );
   nor U10084 ( n10208,n10209,n10210 );
   nor U10085 ( n10210,n6552,n9890 );
   nor U10086 ( n10209,n9894,n6541 );
   nand U10087 ( n6541,n10211,n10212 );
   or U10088 ( n10212,n5965,datai_8_ );
   nand U10089 ( n10211,n5966,n8549 );
   nand U10090 ( n8549,n10213,n10214 );
   nor U10091 ( n10213,n10215,n10216 );
   nor U10092 ( n10216,n6794,n10217 );
   nand U10093 ( n10217,ir_reg_31_,n6792 );
   not U10094 ( n6794,ir_reg_8_ );
   nor U10095 ( n10215,ir_reg_8_,ir_reg_31_ );
   and U10096 ( n9863,n10218,n10219 );
   nand U10097 ( n10219,n10220,n10221 );
   nand U10098 ( n10220,n10222,n9509 );
   or U10099 ( n10218,n9506,n10223 );
   nand U10100 ( n10202,n9666,n9667 );
   or U10101 ( n10200,n9667,n9666 );
   xor U10102 ( n9666,n10224,n6008 );
   nor U10103 ( n10224,n10225,n10226 );
   nor U10104 ( n10226,n6538,n5982 );
   not U10105 ( n6538,n6083 );
   nor U10106 ( n10225,n5991,n6527 );
   nand U10107 ( n9667,n10227,n10228 );
   nand U10108 ( n10228,n5940,n7302 );
   not U10109 ( n7302,n6527 );
   nand U10110 ( n6527,n10229,n10230 );
   or U10111 ( n10230,n5966,datai_9_ );
   nand U10112 ( n10229,n8516,n5964 );
   nand U10113 ( n8516,n10231,n10232 );
   nand U10114 ( n10232,n5987,n6800 );
   not U10115 ( n6800,ir_reg_9_ );
   nand U10116 ( n10231,ir_reg_31_,n6801 );
   nand U10117 ( n6801,n10233,n6807 );
   nand U10118 ( n10233,ir_reg_9_,n10214 );
   nand U10119 ( n10227,n5996,n6083 );
   nand U10120 ( n6083,n10234,n10235 );
   nor U10121 ( n10235,n10236,n10237 );
   nor U10122 ( n10237,n5956,n8538 );
   not U10123 ( n8538,reg1_reg_9_ );
   nor U10124 ( n10236,n7301,n6004 );
   xor U10125 ( n7301,reg3_reg_9_,n10238 );
   nor U10126 ( n10234,n10239,n10240 );
   nor U10127 ( n10240,n10125,n8514 );
   not U10128 ( n8514,reg2_reg_9_ );
   nor U10129 ( n10239,n5961,n10241 );
   not U10130 ( n10241,reg0_reg_9_ );
   nor U10131 ( n9960,n10198,n10199 );
   nand U10132 ( n10199,n10242,n10243 );
   nand U10133 ( n10243,n5940,n7327 );
   nand U10134 ( n10242,n5996,n6080 );
   xor U10135 ( n10198,n6009,n10244 );
   and U10136 ( n10244,n10245,n10246 );
   nand U10137 ( n10246,n7327,n10033 );
   not U10138 ( n7327,n6513 );
   nand U10139 ( n6513,n10247,n10248 );
   or U10140 ( n10248,n5963,datai_10_ );
   nand U10141 ( n10247,n5964,n8493 );
   nand U10142 ( n8493,n10249,n10195 );
   nor U10143 ( n10249,n10250,n10251 );
   nor U10144 ( n10251,n10131,n10252 );
   nand U10145 ( n10252,ir_reg_10_,n6807 );
   nor U10146 ( n10250,ir_reg_31_,ir_reg_10_ );
   nand U10147 ( n10245,n5940,n6080 );
   nand U10148 ( n6080,n10253,n10254 );
   nor U10149 ( n10254,n10255,n10256 );
   nor U10150 ( n10256,n5956,n8505 );
   not U10151 ( n8505,reg1_reg_10_ );
   nor U10152 ( n10255,n6004,n9965 );
   nand U10153 ( n9965,n10257,n10170 );
   nand U10154 ( n10257,n9966,n10258 );
   nand U10155 ( n10258,reg3_reg_9_,n10259 );
   nor U10156 ( n10253,n10260,n10261 );
   nor U10157 ( n10261,n10125,n8492 );
   not U10158 ( n8492,reg2_reg_10_ );
   nor U10159 ( n10260,n5961,n10262 );
   not U10160 ( n10262,reg0_reg_10_ );
   not U10161 ( n9613,n9617 );
   nand U10162 ( n9617,n10150,n10149 );
   nand U10163 ( n10149,n10263,n10264 );
   nand U10164 ( n10264,n5940,n7442 );
   not U10165 ( n7442,n6471 );
   nand U10166 ( n10263,n5996,n6071 );
   xor U10167 ( n10150,n10265,n6008 );
   nor U10168 ( n10265,n10266,n10267 );
   nor U10169 ( n10267,n6482,n9890 );
   not U10170 ( n6482,n6071 );
   nand U10171 ( n6071,n10268,n10269 );
   nor U10172 ( n10269,n10270,n10271 );
   nor U10173 ( n10271,n5954,n8426 );
   not U10174 ( n8426,reg1_reg_13_ );
   nor U10175 ( n10270,n10272,n6005 );
   not U10176 ( n10272,n7441 );
   xor U10177 ( n7441,n9623,n10168 );
   nor U10178 ( n10268,n10273,n10274 );
   nor U10179 ( n10274,n10125,n8402 );
   not U10180 ( n8402,reg2_reg_13_ );
   nor U10181 ( n10273,n5959,n10275 );
   not U10182 ( n10275,reg0_reg_13_ );
   nor U10183 ( n10266,n5990,n6471 );
   nand U10184 ( n6471,n10276,n10277 );
   or U10185 ( n10277,n5966,datai_13_ );
   nand U10186 ( n10276,n8404,n5965 );
   nand U10187 ( n8404,n10278,n10279 );
   nand U10188 ( n10279,n6830,n5987 );
   not U10189 ( n6830,ir_reg_13_ );
   nand U10190 ( n10278,ir_reg_31_,n6831 );
   nand U10191 ( n6831,n10280,n6837 );
   nand U10192 ( n10280,ir_reg_13_,n10159 );
   or U10193 ( n10141,n9992,n9991 );
   xor U10194 ( n9991,n10281,n6009 );
   nor U10195 ( n10281,n10282,n10283 );
   nor U10196 ( n10283,n6468,n5982 );
   not U10197 ( n6468,n6068 );
   nor U10198 ( n10282,n9894,n6457 );
   nand U10199 ( n9992,n10284,n10285 );
   nand U10200 ( n10285,n5940,n7473 );
   not U10201 ( n7473,n6457 );
   nand U10202 ( n6457,n10286,n10287 );
   or U10203 ( n10287,n5965,datai_14_ );
   nand U10204 ( n10286,n5965,n8381 );
   nand U10205 ( n8381,n10288,n10289 );
   nor U10206 ( n10288,n10290,n10291 );
   nor U10207 ( n10291,n10131,n10292 );
   nand U10208 ( n10292,ir_reg_14_,n6837 );
   nor U10209 ( n10290,ir_reg_31_,ir_reg_14_ );
   nand U10210 ( n10284,n5996,n6068 );
   nand U10211 ( n6068,n10293,n10294 );
   nor U10212 ( n10294,n10295,n10296 );
   nor U10213 ( n10296,n5955,n8393 );
   not U10214 ( n8393,reg1_reg_14_ );
   nor U10215 ( n10295,n6004,n7479 );
   nand U10216 ( n7479,n10297,n10298 );
   nand U10217 ( n10297,n9998,n10299 );
   or U10218 ( n10299,n9623,n10168 );
   not U10219 ( n9998,reg3_reg_14_ );
   nor U10220 ( n10293,n10300,n10301 );
   nor U10221 ( n10301,n10125,n8380 );
   not U10222 ( n8380,reg2_reg_14_ );
   nor U10223 ( n10300,n5960,n10302 );
   not U10224 ( n10302,reg0_reg_14_ );
   nand U10225 ( n9452,n10303,n10304 );
   nand U10226 ( n10304,n10021,n7509 );
   not U10227 ( n7509,n6443 );
   nand U10228 ( n6443,n10305,n10306 );
   or U10229 ( n10306,n5966,datai_15_ );
   nand U10230 ( n10305,n8348,n5966 );
   nand U10231 ( n8348,n10307,n10308 );
   nand U10232 ( n10308,n6845,n5987 );
   not U10233 ( n6845,ir_reg_15_ );
   nand U10234 ( n10307,ir_reg_31_,n6846 );
   nand U10235 ( n6846,n10309,n6852 );
   nand U10236 ( n10309,ir_reg_15_,n10289 );
   nand U10237 ( n10303,n10020,n6065 );
   nand U10238 ( n6065,n10310,n10311 );
   nor U10239 ( n10311,n10312,n10313 );
   nor U10240 ( n10313,n5955,n8370 );
   not U10241 ( n8370,reg1_reg_15_ );
   nor U10242 ( n10312,n10314,n6006 );
   not U10243 ( n10314,n7508 );
   xor U10244 ( n7508,n9462,n10298 );
   nor U10245 ( n10310,n10315,n10316 );
   nor U10246 ( n10316,n10125,n8346 );
   not U10247 ( n8346,reg2_reg_15_ );
   nor U10248 ( n10315,n5960,n10317 );
   not U10249 ( n10317,reg0_reg_15_ );
   nand U10250 ( n9723,n9762,n9761 );
   nand U10251 ( n9761,n10318,n10319 );
   nand U10252 ( n10319,n10021,n7542 );
   not U10253 ( n7542,n6429 );
   nand U10254 ( n10318,n10020,n6062 );
   xor U10255 ( n9762,n10320,n6011 );
   nor U10256 ( n10320,n10321,n10322 );
   nor U10257 ( n10322,n6440,n5982 );
   not U10258 ( n6440,n6062 );
   nand U10259 ( n6062,n10323,n10324 );
   nor U10260 ( n10324,n10325,n10326 );
   nor U10261 ( n10326,n5953,n8318 );
   not U10262 ( n8318,reg1_reg_16_ );
   nor U10263 ( n10325,n6004,n9768 );
   nand U10264 ( n9768,n10327,n10122 );
   nand U10265 ( n10327,n9769,n10328 );
   or U10266 ( n10328,n9462,n10298 );
   not U10267 ( n9769,reg3_reg_16_ );
   nor U10268 ( n10323,n10329,n10330 );
   nor U10269 ( n10330,n10125,n8325 );
   not U10270 ( n8325,reg2_reg_16_ );
   nor U10271 ( n10329,n5958,n10331 );
   not U10272 ( n10331,reg0_reg_16_ );
   nor U10273 ( n10321,n5991,n6429 );
   nand U10274 ( n6429,n10332,n10333 );
   or U10275 ( n10333,n5966,datai_16_ );
   nand U10276 ( n10332,n5963,n8326 );
   nand U10277 ( n8326,n10334,n10133 );
   nor U10278 ( n10334,n10335,n10336 );
   nor U10279 ( n10336,n10131,n10337 );
   nand U10280 ( n10337,ir_reg_16_,n6852 );
   nor U10281 ( n10335,ir_reg_31_,ir_reg_16_ );
   nand U10282 ( n10107,n9526,n9527 );
   or U10283 ( n10105,n9527,n9526 );
   xor U10284 ( n9526,n10338,n6009 );
   nor U10285 ( n10338,n10339,n10340 );
   nor U10286 ( n10340,n6412,n5982 );
   not U10287 ( n6412,n6056 );
   nor U10288 ( n10339,n5990,n6401 );
   nand U10289 ( n9527,n10341,n10342 );
   nand U10290 ( n10342,n10021,n7614 );
   not U10291 ( n7614,n6401 );
   nand U10292 ( n6401,n10343,n10344 );
   or U10293 ( n10344,n5965,datai_18_ );
   nand U10294 ( n10343,n5964,n8253 );
   nand U10295 ( n8253,n10345,n10346 );
   nor U10296 ( n10345,n10347,n10348 );
   nor U10297 ( n10348,n10131,n10349 );
   nand U10298 ( n10349,ir_reg_18_,n6867 );
   nor U10299 ( n10347,ir_reg_31_,ir_reg_18_ );
   nand U10300 ( n10341,n10020,n6056 );
   nand U10301 ( n6056,n10350,n10351 );
   nor U10302 ( n10351,n10352,n10353 );
   nor U10303 ( n10353,n5953,n8263 );
   not U10304 ( n8263,reg1_reg_18_ );
   nor U10305 ( n10352,n6005,n7621 );
   nand U10306 ( n7621,n10354,n10071 );
   nand U10307 ( n10354,n9534,n10355 );
   or U10308 ( n10355,n9729,n10122 );
   not U10309 ( n9534,reg3_reg_18_ );
   nor U10310 ( n10350,n10356,n10357 );
   nor U10311 ( n10357,n10125,n8252 );
   not U10312 ( n8252,reg2_reg_18_ );
   nor U10313 ( n10356,n5958,n10358 );
   not U10314 ( n10358,reg0_reg_18_ );
   or U10315 ( n10046,n9590,n9587 );
   xor U10316 ( n9587,n10359,n6008 );
   nor U10317 ( n10359,n10360,n10361 );
   nor U10318 ( n10361,n6356,n5982 );
   not U10319 ( n6356,n6044 );
   nor U10320 ( n10360,n9894,n6345 );
   nand U10321 ( n9590,n10362,n10363 );
   nand U10322 ( n10363,n10021,n7740 );
   not U10323 ( n7740,n6345 );
   nand U10324 ( n6345,datai_22_,n5962 );
   nand U10325 ( n10362,n10020,n6044 );
   nand U10326 ( n6044,n10364,n10365 );
   nor U10327 ( n10365,n10366,n10367 );
   nor U10328 ( n10367,n5956,n10368 );
   not U10329 ( n10368,reg1_reg_22_ );
   nor U10330 ( n10366,n6005,n7746 );
   nand U10331 ( n7746,n10369,n10370 );
   nand U10332 ( n10369,n9596,n10371 );
   or U10333 ( n10371,n9842,n10069 );
   not U10334 ( n9596,reg3_reg_22_ );
   nor U10335 ( n10364,n10372,n10373 );
   and U10336 ( n10373,n9415,reg2_reg_22_ );
   nor U10337 ( n10372,n5961,n10374 );
   not U10338 ( n10374,reg0_reg_22_ );
   nand U10339 ( n9977,n10375,n10376 );
   nand U10340 ( n10376,n10021,n7789 );
   not U10341 ( n7789,n6331 );
   nand U10342 ( n6331,datai_23_,n5962 );
   nand U10343 ( n10375,n10020,n6041 );
   nand U10344 ( n6041,n10377,n10378 );
   nor U10345 ( n10378,n10379,n10380 );
   nor U10346 ( n10380,n5956,n10381 );
   not U10347 ( n10381,reg1_reg_23_ );
   nor U10348 ( n10379,n10382,n6004 );
   not U10349 ( n10382,n7788 );
   xor U10350 ( n7788,n9982,n10370 );
   nor U10351 ( n10377,n10383,n10384 );
   and U10352 ( n10384,n9415,reg2_reg_23_ );
   nor U10353 ( n10383,n5961,n10385 );
   not U10354 ( n10385,reg0_reg_23_ );
   nand U10355 ( n9698,n10039,n10038 );
   nand U10356 ( n10038,n10386,n10387 );
   nand U10357 ( n10387,n10021,n7844 );
   not U10358 ( n7844,n6317 );
   nand U10359 ( n10386,n10020,n6038 );
   xor U10360 ( n10039,n10388,n6010 );
   nor U10361 ( n10388,n10389,n10390 );
   nor U10362 ( n10390,n6328,n9890 );
   not U10363 ( n6328,n6038 );
   nand U10364 ( n6038,n10391,n10392 );
   nor U10365 ( n10392,n10393,n10394 );
   nor U10366 ( n10394,n5954,n10395 );
   not U10367 ( n10395,reg1_reg_24_ );
   nor U10368 ( n10393,n6006,n9704 );
   nand U10369 ( n9704,n10396,n10397 );
   nand U10370 ( n10396,n9705,n10398 );
   or U10371 ( n10398,n9982,n10370 );
   not U10372 ( n9705,reg3_reg_24_ );
   nor U10373 ( n10391,n10399,n10400 );
   and U10374 ( n10400,n9415,reg2_reg_24_ );
   nor U10375 ( n10399,n5959,n10401 );
   not U10376 ( n10401,reg0_reg_24_ );
   nor U10377 ( n10389,n9894,n6317 );
   nand U10378 ( n6317,datai_24_,n5962 );
   nor U10379 ( n9488,n9481,n10402 );
   and U10380 ( n10402,n9479,n9480 );
   nor U10381 ( n10034,n9482,n10403 );
   nor U10382 ( n10403,n9481,n9476 );
   not U10383 ( n9476,n9779 );
   nor U10384 ( n9779,n9480,n9479 );
   not U10385 ( n9479,n9782 );
   nand U10386 ( n9782,n10404,n10405 );
   nand U10387 ( n10405,n10021,n7879 );
   not U10388 ( n7879,n6303 );
   nand U10389 ( n10404,n10020,n6035 );
   xor U10390 ( n9480,n10406,n10015 );
   nor U10391 ( n10406,n10407,n10408 );
   nor U10392 ( n10408,n6314,n5982 );
   not U10393 ( n6314,n6035 );
   nand U10394 ( n6035,n10409,n10410 );
   nor U10395 ( n10410,n10411,n10412 );
   nor U10396 ( n10412,n5954,n10413 );
   not U10397 ( n10413,reg1_reg_25_ );
   nor U10398 ( n10411,n7878,n6006 );
   xor U10399 ( n7878,reg3_reg_25_,n10397 );
   nor U10400 ( n10409,n10414,n10415 );
   and U10401 ( n10415,n9415,reg2_reg_25_ );
   nor U10402 ( n10414,n5959,n10416 );
   not U10403 ( n10416,reg0_reg_25_ );
   nor U10404 ( n10407,n5990,n6303 );
   nand U10405 ( n6303,datai_25_,n5962 );
   nor U10406 ( n9481,n10417,n10418 );
   not U10407 ( n9482,n9486 );
   nand U10408 ( n9486,n10418,n10417 );
   nand U10409 ( n10417,n10419,n10420 );
   nand U10410 ( n10420,n10021,n7905 );
   not U10411 ( n7905,n6289 );
   nand U10412 ( n10419,n10020,n6032 );
   xor U10413 ( n10418,n10421,n6011 );
   nor U10414 ( n10421,n10422,n10423 );
   nor U10415 ( n10423,n6300,n5982 );
   not U10416 ( n6300,n6032 );
   nor U10417 ( n10422,n5991,n6289 );
   nand U10418 ( n6289,datai_26_,n5962 );
   nand U10419 ( n10003,n9454,n6032 );
   nand U10420 ( n6032,n10424,n10425 );
   nor U10421 ( n10425,n10426,n10427 );
   nor U10422 ( n10427,n5953,n10428 );
   not U10423 ( n10428,reg1_reg_26_ );
   nor U10424 ( n10426,n6004,n9496 );
   nand U10425 ( n9496,n10429,n10430 );
   or U10426 ( n10430,n10431,reg3_reg_26_ );
   nor U10427 ( n10424,n10432,n10433 );
   and U10428 ( n10433,n5979,reg2_reg_26_ );
   nor U10429 ( n10432,n5958,n10434 );
   not U10430 ( n10434,reg0_reg_26_ );
   nor U10431 ( n10001,n6272,n9557 );
   not U10432 ( n6272,n6026 );
   nand U10433 ( n6026,n10435,n10436 );
   nor U10434 ( n10436,n10437,n10438 );
   nor U10435 ( n10438,n5955,n10439 );
   not U10436 ( n10439,reg1_reg_28_ );
   nor U10437 ( n10437,n10440,n6006 );
   not U10438 ( n10440,n8034 );
   xor U10439 ( n8034,n9900,reg3_reg_28_ );
   nor U10440 ( n9900,n10429,n10441 );
   nor U10441 ( n10435,n10442,n10443 );
   and U10442 ( n10443,n9415,reg2_reg_28_ );
   nor U10443 ( n10442,n5960,n10444 );
   not U10444 ( n10444,reg0_reg_28_ );
   nor U10445 ( n9999,n10445,n10446 );
   nand U10446 ( n10446,n10447,n10448 );
   nand U10447 ( n10448,n7971,n9495 );
   nand U10448 ( n9495,n10449,n10450 );
   nand U10449 ( n10450,n10451,n6218 );
   nor U10450 ( n10451,n5975,n10452 );
   xor U10451 ( n7971,n10441,n10429 );
   nand U10452 ( n10429,reg3_reg_26_,n10431 );
   nor U10453 ( n10431,n9789,n10397 );
   nand U10454 ( n10397,n10453,reg3_reg_24_ );
   nor U10455 ( n10453,n10370,n9982 );
   not U10456 ( n9982,reg3_reg_23_ );
   nand U10457 ( n10370,n10454,reg3_reg_22_ );
   nor U10458 ( n10454,n10069,n9842 );
   not U10459 ( n9842,reg3_reg_21_ );
   nand U10460 ( n10069,n10455,reg3_reg_20_ );
   nor U10461 ( n10455,n10071,n9930 );
   not U10462 ( n9930,reg3_reg_19_ );
   nand U10463 ( n10071,n10456,reg3_reg_18_ );
   nor U10464 ( n10456,n10122,n9729 );
   not U10465 ( n9729,reg3_reg_17_ );
   nand U10466 ( n10122,n10457,reg3_reg_16_ );
   nor U10467 ( n10457,n10298,n9462 );
   not U10468 ( n9462,reg3_reg_15_ );
   nand U10469 ( n10298,n10458,reg3_reg_14_ );
   nor U10470 ( n10458,n10168,n9623 );
   not U10471 ( n9623,reg3_reg_13_ );
   nand U10472 ( n10168,n10459,reg3_reg_12_ );
   nor U10473 ( n10459,n10170,n9579 );
   not U10474 ( n9579,reg3_reg_11_ );
   nand U10475 ( n10170,n10460,reg3_reg_9_ );
   nor U10476 ( n10460,n10238,n9966 );
   not U10477 ( n9966,reg3_reg_10_ );
   not U10478 ( n9789,reg3_reg_25_ );
   nand U10479 ( n10447,n9494,n7972 );
   not U10480 ( n7972,n6275 );
   nand U10481 ( n6275,datai_27_,n5962 );
   nor U10482 ( n10445,state_reg,n10441 );
   not U10483 ( n10441,reg3_reg_27_ );
   nor U10484 ( n10462,n10463,n10464 );
   nand U10485 ( n10464,n10465,n10466 );
   nand U10486 ( n10466,n10467,n9470 );
   not U10487 ( n9470,n9449 );
   nand U10488 ( n9449,n10468,n10452 );
   nor U10489 ( n10468,n10469,n6979 );
   nor U10490 ( n10467,n10470,n10471 );
   nor U10491 ( n10471,n10472,n10473 );
   nand U10492 ( n10473,n10474,n9509 );
   nand U10493 ( n10474,n9510,n9508 );
   not U10494 ( n9510,n9506 );
   and U10495 ( n10472,n10221,n10222 );
   nor U10496 ( n10470,n10223,n10475 );
   nand U10497 ( n10475,n10476,n10222 );
   nand U10498 ( n10222,n10477,n10478 );
   nand U10499 ( n10476,n9506,n9509 );
   nand U10500 ( n9509,n9513,n9512 );
   nand U10501 ( n9506,n10479,n10480 );
   nand U10502 ( n10480,n9739,n10481 );
   nand U10503 ( n10481,n10482,n9737 );
   and U10504 ( n9739,n10483,n10484 );
   nand U10505 ( n10484,n10021,n7141 );
   not U10506 ( n7141,n6583 );
   nand U10507 ( n10483,n10020,n6095 );
   or U10508 ( n10479,n9737,n10482 );
   not U10509 ( n10482,n9740 );
   nand U10510 ( n9740,n10485,n10486 );
   nand U10511 ( n10486,n10487,n10488 );
   or U10512 ( n10488,n9683,n9681 );
   not U10513 ( n10487,n9682 );
   nand U10514 ( n9682,n10489,n10490 );
   nand U10515 ( n10490,n10021,n7106 );
   not U10516 ( n7106,n6597 );
   nand U10517 ( n10489,n10020,n6098 );
   nand U10518 ( n10485,n9681,n9683 );
   nand U10519 ( n9683,n10491,n10492 );
   not U10520 ( n10492,n9942 );
   nor U10521 ( n9942,n10493,n10494 );
   or U10522 ( n10491,n9941,n9943 );
   and U10523 ( n9943,n10494,n10493 );
   nand U10524 ( n10493,n10495,n10496 );
   nand U10525 ( n10496,n10021,n7079 );
   not U10526 ( n7079,n6611 );
   nand U10527 ( n10495,n10020,n6101 );
   xor U10528 ( n10494,n10497,n6011 );
   nor U10529 ( n10497,n10498,n10499 );
   nor U10530 ( n10499,n6622,n9890 );
   not U10531 ( n6622,n6101 );
   nand U10532 ( n6101,n10500,n10501 );
   nor U10533 ( n10501,n10502,n10503 );
   nor U10534 ( n10503,n5960,n10504 );
   not U10535 ( n10504,reg0_reg_3_ );
   nor U10536 ( n10502,n5955,n10505 );
   not U10537 ( n10505,reg1_reg_3_ );
   nor U10538 ( n10500,n10506,n10507 );
   nor U10539 ( n10507,n5995,n8684 );
   not U10540 ( n8684,reg2_reg_3_ );
   nor U10541 ( n10506,reg3_reg_3_,n6005 );
   nor U10542 ( n10498,n9894,n6611 );
   nand U10543 ( n6611,n10508,n10509 );
   or U10544 ( n10509,n5965,datai_3_ );
   nand U10545 ( n10508,n8686,n5966 );
   not U10546 ( n8686,n8690 );
   nand U10547 ( n8690,n10510,n10511 );
   nand U10548 ( n10511,ir_reg_3_,n5987 );
   nand U10549 ( n10510,n10512,ir_reg_31_ );
   and U10550 ( n10512,n6757,n6756 );
   nand U10551 ( n6756,ir_reg_3_,n10513 );
   nand U10552 ( n9941,n9948,n10514 );
   nand U10553 ( n10514,n9947,n9545 );
   nand U10554 ( n9545,n10515,n9853 );
   nand U10555 ( n9853,n10516,n10517 );
   nand U10556 ( n10515,n10518,n9852 );
   or U10557 ( n9852,n10517,n10516 );
   xor U10558 ( n10516,n10519,n6009 );
   nor U10559 ( n10519,n10520,n10521 );
   nor U10560 ( n10521,n6650,n9890 );
   not U10561 ( n6650,n6107 );
   nor U10562 ( n10520,n5990,n6639 );
   nand U10563 ( n10517,n10522,n10523 );
   nand U10564 ( n10523,n10021,n7011 );
   not U10565 ( n7011,n6639 );
   nand U10566 ( n6639,n10524,n10525 );
   or U10567 ( n10525,n5964,datai_1_ );
   nand U10568 ( n10524,n8760,n5963 );
   not U10569 ( n8760,n8759 );
   xor U10570 ( n8759,n6742,n10526 );
   nand U10571 ( n10526,ir_reg_0_,ir_reg_31_ );
   nand U10572 ( n10522,n10020,n6107 );
   nand U10573 ( n6107,n10527,n10528 );
   nor U10574 ( n10528,n10529,n10530 );
   nor U10575 ( n10530,n5959,n10531 );
   not U10576 ( n10531,reg0_reg_1_ );
   nor U10577 ( n10529,n5954,n8757 );
   not U10578 ( n8757,reg1_reg_1_ );
   nor U10579 ( n10527,n10532,n10533 );
   nor U10580 ( n10533,n5995,n8766 );
   not U10581 ( n8766,reg2_reg_1_ );
   nor U10582 ( n10532,n6005,n8795 );
   not U10583 ( n8795,reg3_reg_1_ );
   not U10584 ( n10518,n9851 );
   nand U10585 ( n9851,n10534,n10535 );
   nand U10586 ( n10535,n6010,n10536 );
   nand U10587 ( n10536,n9654,n9655 );
   or U10588 ( n10534,n9654,n9655 );
   nand U10589 ( n9655,n10537,n10538 );
   nand U10590 ( n10538,ir_reg_0_,n10539 );
   nor U10591 ( n10537,n10540,n10541 );
   nor U10592 ( n10541,n9290,n9889 );
   nor U10593 ( n10540,n6647,n9890 );
   xor U10594 ( n9654,n10015,n10542 );
   nand U10595 ( n10542,n10543,n10544 );
   nand U10596 ( n10544,reg1_reg_0_,n10539 );
   nor U10597 ( n10543,n10545,n10546 );
   nor U10598 ( n10546,n9290,n5982 );
   not U10599 ( n9290,n6110 );
   nand U10600 ( n6110,n10547,n10548 );
   nor U10601 ( n10548,n10549,n10550 );
   nor U10602 ( n10550,n5959,n10551 );
   not U10603 ( n10551,reg0_reg_0_ );
   nor U10604 ( n10549,n5954,n8805 );
   not U10605 ( n8805,reg1_reg_0_ );
   nor U10606 ( n10547,n10552,n10553 );
   and U10607 ( n10553,n9415,reg2_reg_0_ );
   nor U10608 ( n10552,n6006,n6996 );
   not U10609 ( n6996,reg3_reg_0_ );
   nor U10610 ( n10545,n5991,n6647 );
   nand U10611 ( n6647,n10554,n10555 );
   nand U10612 ( n10555,n5963,n8740 );
   or U10613 ( n10554,n5963,datai_0_ );
   not U10614 ( n9947,n9544 );
   nor U10615 ( n9544,n9550,n9551 );
   nand U10616 ( n9948,n9551,n9550 );
   nand U10617 ( n9550,n10556,n10557 );
   nand U10618 ( n10557,n10021,n7032 );
   not U10619 ( n7032,n6625 );
   nand U10620 ( n10556,n10020,n6104 );
   xor U10621 ( n9551,n10558,n6011 );
   nor U10622 ( n10558,n10559,n10560 );
   nor U10623 ( n10560,n6636,n9890 );
   not U10624 ( n6636,n6104 );
   nand U10625 ( n6104,n10561,n10562 );
   nor U10626 ( n10562,n10563,n10564 );
   nor U10627 ( n10564,n5961,n10565 );
   not U10628 ( n10565,reg0_reg_2_ );
   nor U10629 ( n10563,n5956,n8714 );
   not U10630 ( n8714,reg1_reg_2_ );
   nor U10631 ( n10561,n10566,n10567 );
   nor U10632 ( n10567,n5995,n8723 );
   not U10633 ( n8723,reg2_reg_2_ );
   nor U10634 ( n10566,n6006,n8767 );
   not U10635 ( n8767,reg3_reg_2_ );
   nor U10636 ( n10559,n9894,n6625 );
   nand U10637 ( n6625,n10568,n10569 );
   or U10638 ( n10569,n5964,datai_2_ );
   nand U10639 ( n10568,n8718,n5963 );
   nand U10640 ( n8718,n10570,n10571 );
   nand U10641 ( n10571,n6749,n5987 );
   not U10642 ( n6749,ir_reg_2_ );
   nand U10643 ( n10570,ir_reg_31_,n6750 );
   nand U10644 ( n6750,n10513,n10572 );
   nand U10645 ( n10572,ir_reg_2_,n10573 );
   nand U10646 ( n10573,n6742,n8740 );
   not U10647 ( n6742,ir_reg_1_ );
   xor U10648 ( n9681,n10574,n10015 );
   nor U10649 ( n10574,n10575,n10576 );
   nor U10650 ( n10576,n6608,n5982 );
   not U10651 ( n6608,n6098 );
   nand U10652 ( n6098,n10577,n10578 );
   nor U10653 ( n10578,n10579,n10580 );
   nor U10654 ( n10580,n5956,n8675 );
   not U10655 ( n8675,reg1_reg_4_ );
   nor U10656 ( n10579,n6006,n9687 );
   nand U10657 ( n9687,n10581,n10582 );
   nand U10658 ( n10582,n7078,n9688 );
   not U10659 ( n9688,reg3_reg_4_ );
   not U10660 ( n7078,reg3_reg_3_ );
   nor U10661 ( n10577,n10583,n10584 );
   nor U10662 ( n10584,n5995,n8660 );
   not U10663 ( n8660,reg2_reg_4_ );
   nor U10664 ( n10583,n5961,n10585 );
   not U10665 ( n10585,reg0_reg_4_ );
   nor U10666 ( n10575,n5990,n6597 );
   nand U10667 ( n6597,n10586,n10587 );
   or U10668 ( n10587,n5966,datai_4_ );
   nand U10669 ( n10586,n5963,n8661 );
   nand U10670 ( n8661,n10588,n10589 );
   nor U10671 ( n10588,n10590,n10591 );
   nor U10672 ( n10591,n6764,n10592 );
   nand U10673 ( n10592,ir_reg_31_,n6757 );
   not U10674 ( n6764,ir_reg_4_ );
   nor U10675 ( n10590,ir_reg_4_,ir_reg_31_ );
   xor U10676 ( n9737,n10593,n6009 );
   nor U10677 ( n10593,n10594,n10595 );
   nor U10678 ( n10595,n6594,n9890 );
   not U10679 ( n6594,n6095 );
   nand U10680 ( n6095,n10596,n10597 );
   nor U10681 ( n10597,n10598,n10599 );
   nor U10682 ( n10599,n5953,n8650 );
   not U10683 ( n8650,reg1_reg_5_ );
   nor U10684 ( n10598,n10600,n6004 );
   not U10685 ( n10600,n7140 );
   xor U10686 ( n7140,n9745,n10581 );
   nor U10687 ( n10596,n10601,n10602 );
   nor U10688 ( n10602,n5995,n8626 );
   not U10689 ( n8626,reg2_reg_5_ );
   nor U10690 ( n10601,n5958,n10603 );
   not U10691 ( n10603,reg0_reg_5_ );
   nor U10692 ( n10594,n5991,n6583 );
   nand U10693 ( n6583,n10604,n10605 );
   or U10694 ( n10605,n5963,datai_5_ );
   nand U10695 ( n10604,n8628,n5965 );
   nand U10696 ( n8628,n10606,n10607 );
   nand U10697 ( n10607,n5987,n6770 );
   not U10698 ( n6770,ir_reg_5_ );
   nand U10699 ( n10606,ir_reg_31_,n6771 );
   nand U10700 ( n6771,n10608,n6777 );
   nand U10701 ( n10608,ir_reg_5_,n10589 );
   nand U10702 ( n10223,n10221,n9508 );
   nand U10703 ( n9508,n10609,n10610 );
   not U10704 ( n10610,n9513 );
   xor U10705 ( n9513,n10611,n6009 );
   nor U10706 ( n10611,n10612,n10613 );
   nor U10707 ( n10613,n6580,n9890 );
   not U10708 ( n6580,n6092 );
   nor U10709 ( n10612,n9894,n6569 );
   not U10710 ( n9894,n10033 );
   not U10711 ( n10609,n9512 );
   nand U10712 ( n9512,n10614,n10615 );
   nand U10713 ( n10615,n10021,n7175 );
   not U10714 ( n7175,n6569 );
   nand U10715 ( n6569,n10616,n10617 );
   or U10716 ( n10617,n5965,datai_6_ );
   nand U10717 ( n10616,n5965,n8606 );
   nand U10718 ( n8606,n10618,n10619 );
   nor U10719 ( n10618,n10620,n10621 );
   nor U10720 ( n10621,n6779,n10622 );
   nand U10721 ( n10622,ir_reg_31_,n6777 );
   not U10722 ( n6779,ir_reg_6_ );
   nor U10723 ( n10620,ir_reg_6_,ir_reg_31_ );
   nand U10724 ( n10614,n10020,n6092 );
   or U10725 ( n10221,n10477,n10478 );
   nand U10726 ( n10478,n10623,n10624 );
   nand U10727 ( n10624,n5996,n6089 );
   not U10728 ( n10020,n9889 );
   nand U10729 ( n10623,n10021,n7216 );
   xor U10730 ( n10477,n6009,n10625 );
   and U10731 ( n10625,n10626,n10627 );
   nand U10732 ( n10627,n10021,n6089 );
   nand U10733 ( n6089,n10628,n10629 );
   nor U10734 ( n10629,n10630,n10631 );
   nor U10735 ( n10631,n5958,n10632 );
   not U10736 ( n10632,reg0_reg_7_ );
   nor U10737 ( n10630,n5953,n8589 );
   not U10738 ( n8589,reg1_reg_7_ );
   nor U10739 ( n10628,n10633,n10634 );
   nor U10740 ( n10634,n5995,n8570 );
   not U10741 ( n8570,reg2_reg_7_ );
   nor U10742 ( n10633,n10635,n6006 );
   not U10743 ( n10021,n9890 );
   nand U10744 ( n9890,n10636,n10637 );
   nand U10745 ( n10637,n8029,n10638 );
   nand U10746 ( n10626,n7216,n10033 );
   nand U10747 ( n10033,n9889,n10639 );
   nand U10748 ( n10639,n10640,n10636 );
   nand U10749 ( n9889,n10641,n10636 );
   nand U10750 ( n10641,n10642,n8820 );
   nor U10751 ( n8820,n7058,n7835 );
   nor U10752 ( n10642,n6664,n9092 );
   nand U10753 ( n10015,n10643,n10644 );
   nand U10754 ( n10644,n10640,n10645 );
   nand U10755 ( n10465,n9454,n6092 );
   nand U10756 ( n6092,n10646,n10647 );
   nor U10757 ( n10647,n10648,n10649 );
   nor U10758 ( n10649,n5955,n8598 );
   not U10759 ( n8598,reg1_reg_6_ );
   nor U10760 ( n10648,n10650,n6004 );
   not U10761 ( n10650,n7181 );
   xor U10762 ( n7181,n10651,reg3_reg_6_ );
   nor U10763 ( n10646,n10652,n10653 );
   nor U10764 ( n10653,n5995,n8605 );
   not U10765 ( n8605,reg2_reg_6_ );
   nor U10766 ( n10652,n5960,n10654 );
   not U10767 ( n10654,reg0_reg_6_ );
   not U10768 ( n9454,n9489 );
   nand U10769 ( n9489,n10655,n10656 );
   nor U10770 ( n10655,n10657,n8040 );
   nor U10771 ( n10463,n6552,n9557 );
   nand U10772 ( n9557,n10658,n10656 );
   nor U10773 ( n10658,n8732,n10657 );
   not U10774 ( n6552,n6086 );
   nand U10775 ( n6086,n10659,n10660 );
   nor U10776 ( n10660,n10661,n10662 );
   nor U10777 ( n10662,n5960,n10663 );
   not U10778 ( n10663,reg0_reg_8_ );
   nor U10779 ( n10661,n5955,n8561 );
   not U10780 ( n8561,reg1_reg_8_ );
   nor U10781 ( n10659,n10667,n10668 );
   nor U10782 ( n10668,n10125,n8548 );
   not U10783 ( n8548,reg2_reg_8_ );
   not U10784 ( n10125,n9415 );
   nor U10785 ( n9415,n10665,n10666 );
   nor U10786 ( n10667,n6005,n9871 );
   nand U10787 ( n9871,n10669,n10238 );
   not U10788 ( n10238,n10259 );
   nor U10789 ( n10259,n9872,n10670 );
   nand U10790 ( n10669,n9872,n10670 );
   nand U10791 ( n10670,n10671,reg3_reg_7_ );
   and U10792 ( n10671,n10651,reg3_reg_6_ );
   not U10793 ( n9872,reg3_reg_8_ );
   not U10794 ( n10664,n10666 );
   xor U10795 ( n10666,ir_reg_31_,ir_reg_29_ );
   nand U10796 ( n10665,n10672,n10673 );
   nand U10797 ( n10673,n6957,n5987 );
   not U10798 ( n6957,ir_reg_30_ );
   nand U10799 ( n10672,ir_reg_31_,n6958 );
   nand U10800 ( n6958,n6961,n10674 );
   nand U10801 ( n10674,ir_reg_30_,n10675 );
   nand U10802 ( n10675,n10676,n6951 );
   not U10803 ( n6951,ir_reg_29_ );
   nand U10804 ( n6961,n10677,n10676 );
   not U10805 ( n10676,n6949 );
   nor U10806 ( n10677,ir_reg_30_,ir_reg_29_ );
   nor U10807 ( n10461,n10678,n10679 );
   nand U10808 ( n10679,n10680,n10681 );
   nand U10809 ( n10681,n7215,n9460 );
   nand U10810 ( n9460,n10449,n10682 );
   nand U10811 ( n10682,n10683,n6218 );
   nor U10812 ( n10683,n10452,n6979 );
   and U10813 ( n10449,n10684,n10685 );
   nand U10814 ( n10685,n10656,n10657 );
   and U10815 ( n10656,n10686,n8823 );
   nor U10816 ( n10686,n9160,n6979 );
   nand U10817 ( n10684,n10687,state_reg );
   nand U10818 ( n10687,n10688,n10689 );
   nor U10819 ( n10689,n8826,n8236 );
   nor U10820 ( n8236,n8041,n6663 );
   not U10821 ( n8041,n6666 );
   nor U10822 ( n10688,n10690,n8812 );
   nor U10823 ( n10690,n10469,n10452 );
   and U10824 ( n10469,n10691,n10692 );
   nor U10825 ( n10692,n10693,n10694 );
   nand U10826 ( n10694,n8211,n8120 );
   nand U10827 ( n8120,n8823,n9160 );
   not U10828 ( n8823,n10638 );
   nand U10829 ( n10638,n6663,n6668 );
   nor U10830 ( n6663,n6653,n9157 );
   nand U10831 ( n8211,n6254,n8247 );
   not U10832 ( n10693,n7519 );
   nand U10833 ( n7519,n10695,n9092 );
   nor U10834 ( n10695,n6668,n6653 );
   nor U10835 ( n10691,n10696,n10697 );
   nand U10836 ( n10697,n10698,n10699 );
   nand U10837 ( n10699,n7058,n9160 );
   nor U10838 ( n7058,n10643,n6653 );
   nand U10839 ( n10698,n9160,n10700 );
   nand U10840 ( n10700,n8029,n7045 );
   not U10841 ( n7045,n7835 );
   nor U10842 ( n7835,n8247,n10643 );
   nand U10843 ( n10643,n6668,n9157 );
   nand U10844 ( n8029,n10701,n6653 );
   nor U10845 ( n10701,n9157,n10640 );
   nor U10846 ( n10696,n10702,n6668 );
   nor U10847 ( n10702,n8118,n7059 );
   nand U10848 ( n7059,n7770,n7769 );
   nand U10849 ( n7769,n10703,n6653 );
   nor U10850 ( n10703,n8956,n9160 );
   not U10851 ( n7770,n7807 );
   nor U10852 ( n7807,n8247,n5950 );
   not U10853 ( n8819,n9092 );
   nor U10854 ( n9092,n9160,n9157 );
   nor U10855 ( n8118,n10645,n8956 );
   nand U10856 ( n10645,n6667,n8247 );
   not U10857 ( n7215,n10635 );
   xor U10858 ( n10635,reg3_reg_7_,n10704 );
   nand U10859 ( n10704,reg3_reg_6_,n10651 );
   nor U10860 ( n10651,n9745,n10581 );
   nand U10861 ( n10581,reg3_reg_4_,reg3_reg_3_ );
   not U10862 ( n9745,reg3_reg_5_ );
   nand U10863 ( n10680,n9494,n7216 );
   not U10864 ( n7216,n6555 );
   nand U10865 ( n6555,n10705,n10706 );
   or U10866 ( n10706,n5964,datai_7_ );
   nand U10867 ( n10705,n8572,n5964 );
   nand U10868 ( n8572,n10707,n10708 );
   nand U10869 ( n10708,n10131,n6785 );
   not U10870 ( n6785,ir_reg_7_ );
   nand U10871 ( n10707,ir_reg_31_,n6786 );
   nand U10872 ( n6786,n10709,n6792 );
   nand U10873 ( n10709,ir_reg_7_,n10619 );
   not U10874 ( n9494,n9455 );
   nand U10875 ( n9455,n6210,n10710 );
   nand U10876 ( n10710,n8035,n10711 );
   nand U10877 ( n10711,n10452,n6218 );
   nor U10878 ( n6218,n9382,n6667 );
   not U10879 ( n9382,n6664 );
   nor U10880 ( n6664,n8956,n6668 );
   not U10881 ( n6668,n10640 );
   not U10882 ( n10452,n10657 );
   nand U10883 ( n10657,n10712,n6659 );
   not U10884 ( n6659,n8237 );
   nand U10885 ( n8237,n6673,n10713 );
   or U10886 ( n10713,n10714,d_reg_1_ );
   nand U10887 ( n6673,n10715,n10716 );
   nor U10888 ( n10712,n6658,n6212 );
   nand U10889 ( n6212,n6676,n10717 );
   or U10890 ( n10717,n10714,d_reg_0_ );
   nand U10891 ( n6676,n10715,n10718 );
   nand U10892 ( n6658,n10719,n10720 );
   nand U10893 ( n10720,n6980,n10721 );
   nand U10894 ( n10721,n10722,n10723 );
   nor U10895 ( n10723,n10724,n10725 );
   nand U10896 ( n10725,n10726,n10727 );
   nor U10897 ( n10727,d_reg_27_,n10728 );
   nand U10898 ( n10728,n6975,n6976 );
   not U10899 ( n6976,d_reg_29_ );
   not U10900 ( n6975,d_reg_28_ );
   nor U10901 ( n10726,d_reg_26_,d_reg_25_ );
   nand U10902 ( n10724,n10729,n10730 );
   nor U10903 ( n10730,d_reg_3_,n10731 );
   nand U10904 ( n10731,n6962,n6963 );
   not U10905 ( n6963,d_reg_5_ );
   not U10906 ( n6962,d_reg_4_ );
   nor U10907 ( n10729,d_reg_2_,n10732 );
   nand U10908 ( n10732,n6977,n6978 );
   not U10909 ( n6978,d_reg_31_ );
   not U10910 ( n6977,d_reg_30_ );
   nor U10911 ( n10722,n10733,n10734 );
   nand U10912 ( n10734,n10735,n10736 );
   nor U10913 ( n10736,d_reg_17_,n10737 );
   nand U10914 ( n10737,n6971,n6972 );
   not U10915 ( n6972,d_reg_19_ );
   not U10916 ( n6971,d_reg_18_ );
   nor U10917 ( n10735,d_reg_16_,d_reg_13_ );
   nand U10918 ( n10733,n10738,n10739 );
   nor U10919 ( n10739,d_reg_22_,n10740 );
   nand U10920 ( n10740,n6973,n6974 );
   not U10921 ( n6974,d_reg_24_ );
   not U10922 ( n6973,d_reg_23_ );
   nor U10923 ( n10738,d_reg_21_,d_reg_20_ );
   nand U10924 ( n10719,n6980,n10741 );
   nand U10925 ( n10741,n10742,n10743 );
   nor U10926 ( n10743,n10744,n10745 );
   nand U10927 ( n10745,n6970,n6964 );
   not U10928 ( n6964,d_reg_6_ );
   not U10929 ( n6970,d_reg_15_ );
   nand U10930 ( n10744,n10746,n6965 );
   not U10931 ( n6965,d_reg_7_ );
   nor U10932 ( n10746,d_reg_9_,d_reg_8_ );
   nor U10933 ( n10742,n10747,n10748 );
   nand U10934 ( n10748,n6966,n6967 );
   not U10935 ( n6967,d_reg_11_ );
   not U10936 ( n6966,d_reg_10_ );
   nand U10937 ( n10747,n6968,n6969 );
   not U10938 ( n6969,d_reg_14_ );
   not U10939 ( n6968,d_reg_12_ );
   not U10940 ( n6980,n10714 );
   nand U10941 ( n10714,n10749,n10750 );
   nor U10942 ( n10749,n10751,n10752 );
   nor U10943 ( n10752,n10753,n10754 );
   nand U10944 ( n10754,n10716,n10718 );
   not U10945 ( n10753,b_reg );
   nor U10946 ( n10751,b_reg,n10718 );
   nand U10947 ( n8035,n6653,n5997 );
   not U10948 ( n6254,n6223 );
   nand U10949 ( n6223,n6652,n10640 );
   nor U10950 ( n6652,n6667,n9157 );
   not U10951 ( n9157,n8956 );
   nand U10952 ( n8956,n10755,n10756 );
   nor U10953 ( n10755,n10757,n10758 );
   nor U10954 ( n10758,n10131,n10759 );
   nand U10955 ( n10759,ir_reg_20_,n6882 );
   nor U10956 ( n10757,ir_reg_31_,ir_reg_20_ );
   not U10957 ( n6667,n9160 );
   not U10958 ( n6653,n8247 );
   nand U10959 ( n8247,n10760,n10761 );
   nand U10960 ( n10761,n6875,n5987 );
   not U10961 ( n6875,ir_reg_19_ );
   nand U10962 ( n10760,ir_reg_31_,n6876 );
   nand U10963 ( n6876,n10762,n6882 );
   nand U10964 ( n10762,ir_reg_19_,n10346 );
   not U10965 ( n6210,n6979 );
   nand U10966 ( n6979,n10763,n9270 );
   nor U10967 ( n10763,n5932,n10539 );
   and U10968 ( n10678,n5932,reg3_reg_7_ );
   nand U10969 ( n6016,n8826,state_reg );
   nor U10970 ( n8826,n10636,n8812 );
   not U10971 ( n8812,n9270 );
   not U10972 ( n10636,n10539 );
   nor U10973 ( n10539,n10765,n10718 );
   nand U10974 ( n10718,n10766,n10767 );
   nor U10975 ( n10766,n10768,n10769 );
   nor U10976 ( n10769,n10131,n10770 );
   nand U10977 ( n10770,ir_reg_24_,n6912 );
   nor U10978 ( n10768,ir_reg_31_,ir_reg_24_ );
   or U10979 ( n10765,n10715,n10716 );
   nand U10980 ( n10716,n10771,n10772 );
   nand U10981 ( n10772,n6920,n5987 );
   not U10982 ( n6920,ir_reg_25_ );
   nand U10983 ( n10771,ir_reg_31_,n6921 );
   nand U10984 ( n6921,n10773,n10774 );
   nand U10985 ( n10774,ir_reg_25_,n10767 );
   not U10986 ( n10715,n10750 );
   nand U10987 ( n10750,n10775,n10776 );
   nand U10988 ( n10776,n10777,n6927 );
   nand U10989 ( n6927,ir_reg_26_,n10773 );
   nand U10990 ( n10775,ir_reg_26_,n5987 );
   nand U10991 ( n10764,n10778,state_reg );
   nand U10992 ( n10778,n10779,n5962 );
   not U10993 ( n8732,n8040 );
   nand U10994 ( n8040,n10780,n10781 );
   nand U10995 ( n10781,n6942,n5987 );
   not U10996 ( n6942,ir_reg_28_ );
   nand U10997 ( n10780,ir_reg_31_,n6943 );
   nand U10998 ( n6943,n10782,n6949 );
   nand U10999 ( n6949,n10783,n6937 );
   nor U11000 ( n10783,ir_reg_28_,ir_reg_27_ );
   nand U11001 ( n10782,ir_reg_28_,n10784 );
   nand U11002 ( n10784,n6937,n6935 );
   not U11003 ( n6935,ir_reg_27_ );
   xor U11004 ( n8734,n10777,ir_reg_27_ );
   nor U11005 ( n10777,n10131,n6937 );
   nor U11006 ( n6937,n10773,ir_reg_26_ );
   or U11007 ( n10773,n10767,ir_reg_25_ );
   or U11008 ( n10767,n6912,ir_reg_24_ );
   nand U11009 ( n10779,n6666,n9270 );
   nand U11010 ( n9270,n10785,n10786 );
   nand U11011 ( n10786,n6905,n5987 );
   not U11012 ( n6905,ir_reg_23_ );
   nand U11013 ( n10785,ir_reg_31_,n6906 );
   nand U11014 ( n6906,n6912,n10787 );
   nand U11015 ( n10787,ir_reg_23_,n10788 );
   or U11016 ( n6912,n10788,ir_reg_23_ );
   nor U11017 ( n6666,n9160,n10640 );
   nand U11018 ( n10640,n10789,n10790 );
   nand U11019 ( n10790,n6890,n5987 );
   not U11020 ( n6890,ir_reg_21_ );
   nand U11021 ( n10789,ir_reg_31_,n6891 );
   nand U11022 ( n6891,n10791,n6897 );
   nand U11023 ( n10791,ir_reg_21_,n10756 );
   nand U11024 ( n9160,n10792,n10788 );
   or U11025 ( n10788,n6897,ir_reg_22_ );
   nor U11026 ( n10792,n10793,n10794 );
   nor U11027 ( n10794,n10131,n10795 );
   nand U11028 ( n10795,ir_reg_22_,n6897 );
   or U11029 ( n6897,n10756,ir_reg_21_ );
   or U11030 ( n10756,n6882,ir_reg_20_ );
   or U11031 ( n6882,n10346,ir_reg_19_ );
   or U11032 ( n10346,n6867,ir_reg_18_ );
   or U11033 ( n6867,n10133,ir_reg_17_ );
   or U11034 ( n10133,n6852,ir_reg_16_ );
   or U11035 ( n6852,n10289,ir_reg_15_ );
   or U11036 ( n10289,n6837,ir_reg_14_ );
   or U11037 ( n6837,n10159,ir_reg_13_ );
   or U11038 ( n10159,n6822,ir_reg_12_ );
   or U11039 ( n6822,n10195,ir_reg_11_ );
   or U11040 ( n10195,n6807,ir_reg_10_ );
   or U11041 ( n6807,n10214,ir_reg_9_ );
   or U11042 ( n10214,n6792,ir_reg_8_ );
   or U11043 ( n6792,n10619,ir_reg_7_ );
   or U11044 ( n10619,n6777,ir_reg_6_ );
   or U11045 ( n6777,n10589,ir_reg_5_ );
   or U11046 ( n10589,n6757,ir_reg_4_ );
   or U11047 ( n6757,n10513,ir_reg_3_ );
   nand U11048 ( n10513,n10796,n8740 );
   not U11049 ( n8740,ir_reg_0_ );
   nor U11050 ( n10796,ir_reg_2_,ir_reg_1_ );
   not U11051 ( n10131,ir_reg_31_ );
   nor U11052 ( n10793,ir_reg_31_,ir_reg_22_ );
endmodule
