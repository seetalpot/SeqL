
module b15 ( datai_31_, datai_30_, datai_29_, datai_28_, datai_27_, datai_26_,
datai_25_, datai_24_, datai_23_, datai_22_, datai_21_, datai_20_,
datai_19_, datai_18_, datai_17_, datai_16_, datai_15_, datai_14_,
datai_13_, datai_12_, datai_11_, datai_10_, datai_9_, datai_8_,
datai_7_, datai_6_, datai_5_, datai_4_, datai_3_, datai_2_, datai_1_,
datai_0_, na_n, bs16_n, ready_n, hold, be_n_reg_3_, be_n_reg_2_,
be_n_reg_1_, be_n_reg_0_, address_reg_29_, address_reg_28_,
address_reg_27_, address_reg_26_, address_reg_25_, address_reg_24_,
address_reg_23_, address_reg_22_, address_reg_21_, address_reg_20_,
address_reg_19_, address_reg_18_, address_reg_17_, address_reg_16_,
address_reg_15_, address_reg_14_, address_reg_13_, address_reg_12_,
address_reg_11_, address_reg_10_, address_reg_9_, address_reg_8_,
address_reg_7_, address_reg_6_, address_reg_5_, address_reg_4_,
address_reg_3_, address_reg_2_, address_reg_1_, address_reg_0_,
state_reg_2_, state_reg_1_, state_reg_0_, datawidth_reg_0_,
datawidth_reg_1_, datawidth_reg_2_, datawidth_reg_3_, datawidth_reg_4_,
datawidth_reg_5_, datawidth_reg_6_, datawidth_reg_7_, datawidth_reg_8_,
datawidth_reg_9_, datawidth_reg_10_, datawidth_reg_11_,
datawidth_reg_12_, datawidth_reg_13_, datawidth_reg_14_,
datawidth_reg_15_, datawidth_reg_16_, datawidth_reg_17_,
datawidth_reg_18_, datawidth_reg_19_, datawidth_reg_20_,
datawidth_reg_21_, datawidth_reg_22_, datawidth_reg_23_,
datawidth_reg_24_, datawidth_reg_25_, datawidth_reg_26_,
datawidth_reg_27_, datawidth_reg_28_, datawidth_reg_29_,
datawidth_reg_30_, datawidth_reg_31_, state2_reg_3_, state2_reg_2_,
state2_reg_1_, state2_reg_0_, instqueue_reg_15__7_,
instqueue_reg_15__6_, instqueue_reg_15__5_, instqueue_reg_15__4_,
instqueue_reg_15__3_, instqueue_reg_15__2_, instqueue_reg_15__1_,
instqueue_reg_15__0_, instqueue_reg_14__7_, instqueue_reg_14__6_,
instqueue_reg_14__5_, instqueue_reg_14__4_, instqueue_reg_14__3_,
instqueue_reg_14__2_, instqueue_reg_14__1_, instqueue_reg_14__0_,
instqueue_reg_13__7_, instqueue_reg_13__6_, instqueue_reg_13__5_,
instqueue_reg_13__4_, instqueue_reg_13__3_, instqueue_reg_13__2_,
instqueue_reg_13__1_, instqueue_reg_13__0_, instqueue_reg_12__7_,
instqueue_reg_12__6_, instqueue_reg_12__5_, instqueue_reg_12__4_,
instqueue_reg_12__3_, instqueue_reg_12__2_, instqueue_reg_12__1_,
instqueue_reg_12__0_, instqueue_reg_11__7_, instqueue_reg_11__6_,
instqueue_reg_11__5_, instqueue_reg_11__4_, instqueue_reg_11__3_,
instqueue_reg_11__2_, instqueue_reg_11__1_, instqueue_reg_11__0_,
instqueue_reg_10__7_, instqueue_reg_10__6_, instqueue_reg_10__5_,
instqueue_reg_10__4_, instqueue_reg_10__3_, instqueue_reg_10__2_,
instqueue_reg_10__1_, instqueue_reg_10__0_, instqueue_reg_9__7_,
instqueue_reg_9__6_, instqueue_reg_9__5_, instqueue_reg_9__4_,
instqueue_reg_9__3_, instqueue_reg_9__2_, instqueue_reg_9__1_,
instqueue_reg_9__0_, instqueue_reg_8__7_, instqueue_reg_8__6_,
instqueue_reg_8__5_, instqueue_reg_8__4_, instqueue_reg_8__3_,
instqueue_reg_8__2_, instqueue_reg_8__1_, instqueue_reg_8__0_,
instqueue_reg_7__7_, instqueue_reg_7__6_, instqueue_reg_7__5_,
instqueue_reg_7__4_, instqueue_reg_7__3_, instqueue_reg_7__2_,
instqueue_reg_7__1_, instqueue_reg_7__0_, instqueue_reg_6__7_,
instqueue_reg_6__6_, instqueue_reg_6__5_, instqueue_reg_6__4_,
instqueue_reg_6__3_, instqueue_reg_6__2_, instqueue_reg_6__1_,
instqueue_reg_6__0_, instqueue_reg_5__7_, instqueue_reg_5__6_,
instqueue_reg_5__5_, instqueue_reg_5__4_, instqueue_reg_5__3_,
instqueue_reg_5__2_, instqueue_reg_5__1_, instqueue_reg_5__0_,
instqueue_reg_4__7_, instqueue_reg_4__6_, instqueue_reg_4__5_,
instqueue_reg_4__4_, instqueue_reg_4__3_, instqueue_reg_4__2_,
instqueue_reg_4__1_, instqueue_reg_4__0_, instqueue_reg_3__7_,
instqueue_reg_3__6_, instqueue_reg_3__5_, instqueue_reg_3__4_,
instqueue_reg_3__3_, instqueue_reg_3__2_, instqueue_reg_3__1_,
instqueue_reg_3__0_, instqueue_reg_2__7_, instqueue_reg_2__6_,
instqueue_reg_2__5_, instqueue_reg_2__4_, instqueue_reg_2__3_,
instqueue_reg_2__2_, instqueue_reg_2__1_, instqueue_reg_2__0_,
instqueue_reg_1__7_, instqueue_reg_1__6_, instqueue_reg_1__5_,
instqueue_reg_1__4_, instqueue_reg_1__3_, instqueue_reg_1__2_,
instqueue_reg_1__1_, instqueue_reg_1__0_, instqueue_reg_0__7_,
instqueue_reg_0__6_, instqueue_reg_0__5_, instqueue_reg_0__4_,
instqueue_reg_0__3_, instqueue_reg_0__2_, instqueue_reg_0__1_,
instqueue_reg_0__0_, instqueuerd_addr_reg_4_, instqueuerd_addr_reg_3_,
instqueuerd_addr_reg_2_, instqueuerd_addr_reg_1_,
instqueuerd_addr_reg_0_, instqueuewr_addr_reg_4_,
instqueuewr_addr_reg_3_, instqueuewr_addr_reg_2_,
instqueuewr_addr_reg_1_, instqueuewr_addr_reg_0_,
instaddrpointer_reg_0_, instaddrpointer_reg_1_, instaddrpointer_reg_2_,
instaddrpointer_reg_3_, instaddrpointer_reg_4_, instaddrpointer_reg_5_,
instaddrpointer_reg_6_, instaddrpointer_reg_7_, instaddrpointer_reg_8_,
instaddrpointer_reg_9_, instaddrpointer_reg_10_,
instaddrpointer_reg_11_, instaddrpointer_reg_12_,
instaddrpointer_reg_13_, instaddrpointer_reg_14_,
instaddrpointer_reg_15_, instaddrpointer_reg_16_,
instaddrpointer_reg_17_, instaddrpointer_reg_18_,
instaddrpointer_reg_19_, instaddrpointer_reg_20_,
instaddrpointer_reg_21_, instaddrpointer_reg_22_,
instaddrpointer_reg_23_, instaddrpointer_reg_24_,
instaddrpointer_reg_25_, instaddrpointer_reg_26_,
instaddrpointer_reg_27_, instaddrpointer_reg_28_,
instaddrpointer_reg_29_, instaddrpointer_reg_30_,
instaddrpointer_reg_31_, phyaddrpointer_reg_0_, phyaddrpointer_reg_1_,
phyaddrpointer_reg_2_, phyaddrpointer_reg_3_, phyaddrpointer_reg_4_,
phyaddrpointer_reg_5_, phyaddrpointer_reg_6_, phyaddrpointer_reg_7_,
phyaddrpointer_reg_8_, phyaddrpointer_reg_9_, phyaddrpointer_reg_10_,
phyaddrpointer_reg_11_, phyaddrpointer_reg_12_, phyaddrpointer_reg_13_,
phyaddrpointer_reg_14_, phyaddrpointer_reg_15_, phyaddrpointer_reg_16_,
phyaddrpointer_reg_17_, phyaddrpointer_reg_18_, phyaddrpointer_reg_19_,
phyaddrpointer_reg_20_, phyaddrpointer_reg_21_, phyaddrpointer_reg_22_,
phyaddrpointer_reg_23_, phyaddrpointer_reg_24_, phyaddrpointer_reg_25_,
phyaddrpointer_reg_26_, phyaddrpointer_reg_27_, phyaddrpointer_reg_28_,
phyaddrpointer_reg_29_, phyaddrpointer_reg_30_, phyaddrpointer_reg_31_,
lword_reg_15_, lword_reg_14_, lword_reg_13_, lword_reg_12_,
lword_reg_11_, lword_reg_10_, lword_reg_9_, lword_reg_8_, lword_reg_7_,
lword_reg_6_, lword_reg_5_, lword_reg_4_, lword_reg_3_, lword_reg_2_,
lword_reg_1_, lword_reg_0_, uword_reg_14_, uword_reg_13_,
uword_reg_12_, uword_reg_11_, uword_reg_10_, uword_reg_9_,
uword_reg_8_, uword_reg_7_, uword_reg_6_, uword_reg_5_, uword_reg_4_,
uword_reg_3_, uword_reg_2_, uword_reg_1_, uword_reg_0_, datao_reg_0_,
datao_reg_1_, datao_reg_2_, datao_reg_3_, datao_reg_4_, datao_reg_5_,
datao_reg_6_, datao_reg_7_, datao_reg_8_, datao_reg_9_, datao_reg_10_,
datao_reg_11_, datao_reg_12_, datao_reg_13_, datao_reg_14_,
datao_reg_15_, datao_reg_16_, datao_reg_17_, datao_reg_18_,
datao_reg_19_, datao_reg_20_, datao_reg_21_, datao_reg_22_,
datao_reg_23_, datao_reg_24_, datao_reg_25_, datao_reg_26_,
datao_reg_27_, datao_reg_28_, datao_reg_29_, datao_reg_30_,
datao_reg_31_, eax_reg_0_, eax_reg_1_, eax_reg_2_, eax_reg_3_,
eax_reg_4_, eax_reg_5_, eax_reg_6_, eax_reg_7_, eax_reg_8_, eax_reg_9_,
eax_reg_10_, eax_reg_11_, eax_reg_12_, eax_reg_13_, eax_reg_14_,
eax_reg_15_, eax_reg_16_, eax_reg_17_, eax_reg_18_, eax_reg_19_,
eax_reg_20_, eax_reg_21_, eax_reg_22_, eax_reg_23_, eax_reg_24_,
eax_reg_25_, eax_reg_26_, eax_reg_27_, eax_reg_28_, eax_reg_29_,
eax_reg_30_, eax_reg_31_, ebx_reg_0_, ebx_reg_1_, ebx_reg_2_,
ebx_reg_3_, ebx_reg_4_, ebx_reg_5_, ebx_reg_6_, ebx_reg_7_, ebx_reg_8_,
ebx_reg_9_, ebx_reg_10_, ebx_reg_11_, ebx_reg_12_, ebx_reg_13_,
ebx_reg_14_, ebx_reg_15_, ebx_reg_16_, ebx_reg_17_, ebx_reg_18_,
ebx_reg_19_, ebx_reg_20_, ebx_reg_21_, ebx_reg_22_, ebx_reg_23_,
ebx_reg_24_, ebx_reg_25_, ebx_reg_26_, ebx_reg_27_, ebx_reg_28_,
ebx_reg_29_, ebx_reg_30_, ebx_reg_31_, reip_reg_0_, reip_reg_1_,
reip_reg_2_, reip_reg_3_, reip_reg_4_, reip_reg_5_, reip_reg_6_,
reip_reg_7_, reip_reg_8_, reip_reg_9_, reip_reg_10_, reip_reg_11_,
reip_reg_12_, reip_reg_13_, reip_reg_14_, reip_reg_15_, reip_reg_16_,
reip_reg_17_, reip_reg_18_, reip_reg_19_, reip_reg_20_, reip_reg_21_,
reip_reg_22_, reip_reg_23_, reip_reg_24_, reip_reg_25_, reip_reg_26_,
reip_reg_27_, reip_reg_28_, reip_reg_29_, reip_reg_30_, reip_reg_31_,
byteenable_reg_3_, byteenable_reg_2_, byteenable_reg_1_,
byteenable_reg_0_, w_r_n_reg, flush_reg, more_reg, statebs16_reg,
requestpending_reg, d_c_n_reg, m_io_n_reg, codefetch_reg, ads_n_reg,
readrequest_reg, memoryfetch_reg, u3445, u3446, u3447, u3448, u3213,
u3212, u3211, u3210, u3209, u3208, u3207, u3206, u3205, u3204, u3203,
u3202, u3201, u3200, u3199, u3198, u3197, u3196, u3195, u3194, u3193,
u3192, u3191, u3190, u3189, u3188, u3187, u3186, u3185, u3184, u3183,
u3182, u3181, u3451, u3452, u3180, u3179, u3178, u3177, u3176, u3175,
u3174, u3173, u3172, u3171, u3170, u3169, u3168, u3167, u3166, u3165,
u3164, u3163, u3162, u3161, u3160, u3159, u3158, u3157, u3156, u3155,
u3154, u3153, u3152, u3151, u3453, u3150, u3149, u3148, u3147, u3146,
u3145, u3144, u3143, u3142, u3141, u3140, u3139, u3138, u3137, u3136,
u3135, u3134, u3133, u3132, u3131, u3130, u3129, u3128, u3127, u3126,
u3125, u3124, u3123, u3122, u3121, u3120, u3119, u3118, u3117, u3116,
u3115, u3114, u3113, u3112, u3111, u3110, u3109, u3108, u3107, u3106,
u3105, u3104, u3103, u3102, u3101, u3100, u3099, u3098, u3097, u3096,
u3095, u3094, u3093, u3092, u3091, u3090, u3089, u3088, u3087, u3086,
u3085, u3084, u3083, u3082, u3081, u3080, u3079, u3078, u3077, u3076,
u3075, u3074, u3073, u3072, u3071, u3070, u3069, u3068, u3067, u3066,
u3065, u3064, u3063, u3062, u3061, u3060, u3059, u3058, u3057, u3056,
u3055, u3054, u3053, u3052, u3051, u3050, u3049, u3048, u3047, u3046,
u3045, u3044, u3043, u3042, u3041, u3040, u3039, u3038, u3037, u3036,
u3035, u3034, u3033, u3032, u3031, u3030, u3029, u3028, u3027, u3026,
u3025, u3024, u3023, u3022, u3021, u3020, u3455, u3456, u3459, u3460,
u3461, u3019, u3462, u3463, u3464, u3465, u3018, u3017, u3016, u3015,
u3014, u3013, u3012, u3011, u3010, u3009, u3008, u3007, u3006, u3005,
u3004, u3003, u3002, u3001, u3000, u2999, u2998, u2997, u2996, u2995,
u2994, u2993, u2992, u2991, u2990, u2989, u2988, u2987, u2986, u2985,
u2984, u2983, u2982, u2981, u2980, u2979, u2978, u2977, u2976, u2975,
u2974, u2973, u2972, u2971, u2970, u2969, u2968, u2967, u2966, u2965,
u2964, u2963, u2962, u2961, u2960, u2959, u2958, u2957, u2956, u2955,
u2954, u2953, u2952, u2951, u2950, u2949, u2948, u2947, u2946, u2945,
u2944, u2943, u2942, u2941, u2940, u2939, u2938, u2937, u2936, u2935,
u2934, u2933, u2932, u2931, u2930, u2929, u2928, u2927, u2926, u2925,
u2924, u2923, u2922, u2921, u2920, u2919, u2918, u2917, u2916, u2915,
u2914, u2913, u2912, u2911, u2910, u2909, u2908, u2907, u2906, u2905,
u2904, u2903, u2902, u2901, u2900, u2899, u2898, u2897, u2896, u2895,
u2894, u2893, u2892, u2891, u2890, u2889, u2888, u2887, u2886, u2885,
u2884, u2883, u2882, u2881, u2880, u2879, u2878, u2877, u2876, u2875,
u2874, u2873, u2872, u2871, u2870, u2869, u2868, u2867, u2866, u2865,
u2864, u2863, u2862, u2861, u2860, u2859, u2858, u2857, u2856, u2855,
u2854, u2853, u2852, u2851, u2850, u2849, u2848, u2847, u2846, u2845,
u2844, u2843, u2842, u2841, u2840, u2839, u2838, u2837, u2836, u2835,
u2834, u2833, u2832, u2831, u2830, u2829, u2828, u2827, u2826, u2825,
u2824, u2823, u2822, u2821, u2820, u2819, u2818, u2817, u2816, u2815,
u2814, u2813, u2812, u2811, u2810, u2809, u2808, u2807, u2806, u2805,
u2804, u2803, u2802, u2801, u2800, u2799, u2798, u2797, u2796, u2795,
u3468, u2794, u3469, u3470, u2793, u3471, u2792, u3472, u2791, u3473,
u2790, u2789, u3474, u2788 );
input datai_31_, datai_30_, datai_29_, datai_28_, datai_27_, datai_26_,
datai_25_, datai_24_, datai_23_, datai_22_, datai_21_, datai_20_,
datai_19_, datai_18_, datai_17_, datai_16_, datai_15_, datai_14_,
datai_13_, datai_12_, datai_11_, datai_10_, datai_9_, datai_8_,
datai_7_, datai_6_, datai_5_, datai_4_, datai_3_, datai_2_, datai_1_,
datai_0_, na_n, bs16_n, ready_n, hold, be_n_reg_3_, be_n_reg_2_,
be_n_reg_1_, be_n_reg_0_, address_reg_29_, address_reg_28_,
address_reg_27_, address_reg_26_, address_reg_25_, address_reg_24_,
address_reg_23_, address_reg_22_, address_reg_21_, address_reg_20_,
address_reg_19_, address_reg_18_, address_reg_17_, address_reg_16_,
address_reg_15_, address_reg_14_, address_reg_13_, address_reg_12_,
address_reg_11_, address_reg_10_, address_reg_9_, address_reg_8_,
address_reg_7_, address_reg_6_, address_reg_5_, address_reg_4_,
address_reg_3_, address_reg_2_, address_reg_1_, address_reg_0_,
state_reg_2_, state_reg_1_, state_reg_0_, datawidth_reg_0_,
datawidth_reg_1_, datawidth_reg_2_, datawidth_reg_3_,
datawidth_reg_4_, datawidth_reg_5_, datawidth_reg_6_,
datawidth_reg_7_, datawidth_reg_8_, datawidth_reg_9_,
datawidth_reg_10_, datawidth_reg_11_, datawidth_reg_12_,
datawidth_reg_13_, datawidth_reg_14_, datawidth_reg_15_,
datawidth_reg_16_, datawidth_reg_17_, datawidth_reg_18_,
datawidth_reg_19_, datawidth_reg_20_, datawidth_reg_21_,
datawidth_reg_22_, datawidth_reg_23_, datawidth_reg_24_,
datawidth_reg_25_, datawidth_reg_26_, datawidth_reg_27_,
datawidth_reg_28_, datawidth_reg_29_, datawidth_reg_30_,
datawidth_reg_31_, state2_reg_3_, state2_reg_2_, state2_reg_1_,
state2_reg_0_, instqueue_reg_15__7_, instqueue_reg_15__6_,
instqueue_reg_15__5_, instqueue_reg_15__4_, instqueue_reg_15__3_,
instqueue_reg_15__2_, instqueue_reg_15__1_, instqueue_reg_15__0_,
instqueue_reg_14__7_, instqueue_reg_14__6_, instqueue_reg_14__5_,
instqueue_reg_14__4_, instqueue_reg_14__3_, instqueue_reg_14__2_,
instqueue_reg_14__1_, instqueue_reg_14__0_, instqueue_reg_13__7_,
instqueue_reg_13__6_, instqueue_reg_13__5_, instqueue_reg_13__4_,
instqueue_reg_13__3_, instqueue_reg_13__2_, instqueue_reg_13__1_,
instqueue_reg_13__0_, instqueue_reg_12__7_, instqueue_reg_12__6_,
instqueue_reg_12__5_, instqueue_reg_12__4_, instqueue_reg_12__3_,
instqueue_reg_12__2_, instqueue_reg_12__1_, instqueue_reg_12__0_,
instqueue_reg_11__7_, instqueue_reg_11__6_, instqueue_reg_11__5_,
instqueue_reg_11__4_, instqueue_reg_11__3_, instqueue_reg_11__2_,
instqueue_reg_11__1_, instqueue_reg_11__0_, instqueue_reg_10__7_,
instqueue_reg_10__6_, instqueue_reg_10__5_, instqueue_reg_10__4_,
instqueue_reg_10__3_, instqueue_reg_10__2_, instqueue_reg_10__1_,
instqueue_reg_10__0_, instqueue_reg_9__7_, instqueue_reg_9__6_,
instqueue_reg_9__5_, instqueue_reg_9__4_, instqueue_reg_9__3_,
instqueue_reg_9__2_, instqueue_reg_9__1_, instqueue_reg_9__0_,
instqueue_reg_8__7_, instqueue_reg_8__6_, instqueue_reg_8__5_,
instqueue_reg_8__4_, instqueue_reg_8__3_, instqueue_reg_8__2_,
instqueue_reg_8__1_, instqueue_reg_8__0_, instqueue_reg_7__7_,
instqueue_reg_7__6_, instqueue_reg_7__5_, instqueue_reg_7__4_,
instqueue_reg_7__3_, instqueue_reg_7__2_, instqueue_reg_7__1_,
instqueue_reg_7__0_, instqueue_reg_6__7_, instqueue_reg_6__6_,
instqueue_reg_6__5_, instqueue_reg_6__4_, instqueue_reg_6__3_,
instqueue_reg_6__2_, instqueue_reg_6__1_, instqueue_reg_6__0_,
instqueue_reg_5__7_, instqueue_reg_5__6_, instqueue_reg_5__5_,
instqueue_reg_5__4_, instqueue_reg_5__3_, instqueue_reg_5__2_,
instqueue_reg_5__1_, instqueue_reg_5__0_, instqueue_reg_4__7_,
instqueue_reg_4__6_, instqueue_reg_4__5_, instqueue_reg_4__4_,
instqueue_reg_4__3_, instqueue_reg_4__2_, instqueue_reg_4__1_,
instqueue_reg_4__0_, instqueue_reg_3__7_, instqueue_reg_3__6_,
instqueue_reg_3__5_, instqueue_reg_3__4_, instqueue_reg_3__3_,
instqueue_reg_3__2_, instqueue_reg_3__1_, instqueue_reg_3__0_,
instqueue_reg_2__7_, instqueue_reg_2__6_, instqueue_reg_2__5_,
instqueue_reg_2__4_, instqueue_reg_2__3_, instqueue_reg_2__2_,
instqueue_reg_2__1_, instqueue_reg_2__0_, instqueue_reg_1__7_,
instqueue_reg_1__6_, instqueue_reg_1__5_, instqueue_reg_1__4_,
instqueue_reg_1__3_, instqueue_reg_1__2_, instqueue_reg_1__1_,
instqueue_reg_1__0_, instqueue_reg_0__7_, instqueue_reg_0__6_,
instqueue_reg_0__5_, instqueue_reg_0__4_, instqueue_reg_0__3_,
instqueue_reg_0__2_, instqueue_reg_0__1_, instqueue_reg_0__0_,
instqueuerd_addr_reg_4_, instqueuerd_addr_reg_3_,
instqueuerd_addr_reg_2_, instqueuerd_addr_reg_1_,
instqueuerd_addr_reg_0_, instqueuewr_addr_reg_4_,
instqueuewr_addr_reg_3_, instqueuewr_addr_reg_2_,
instqueuewr_addr_reg_1_, instqueuewr_addr_reg_0_,
instaddrpointer_reg_0_, instaddrpointer_reg_1_,
instaddrpointer_reg_2_, instaddrpointer_reg_3_,
instaddrpointer_reg_4_, instaddrpointer_reg_5_,
instaddrpointer_reg_6_, instaddrpointer_reg_7_,
instaddrpointer_reg_8_, instaddrpointer_reg_9_,
instaddrpointer_reg_10_, instaddrpointer_reg_11_,
instaddrpointer_reg_12_, instaddrpointer_reg_13_,
instaddrpointer_reg_14_, instaddrpointer_reg_15_,
instaddrpointer_reg_16_, instaddrpointer_reg_17_,
instaddrpointer_reg_18_, instaddrpointer_reg_19_,
instaddrpointer_reg_20_, instaddrpointer_reg_21_,
instaddrpointer_reg_22_, instaddrpointer_reg_23_,
instaddrpointer_reg_24_, instaddrpointer_reg_25_,
instaddrpointer_reg_26_, instaddrpointer_reg_27_,
instaddrpointer_reg_28_, instaddrpointer_reg_29_,
instaddrpointer_reg_30_, instaddrpointer_reg_31_,
phyaddrpointer_reg_0_, phyaddrpointer_reg_1_, phyaddrpointer_reg_2_,
phyaddrpointer_reg_3_, phyaddrpointer_reg_4_, phyaddrpointer_reg_5_,
phyaddrpointer_reg_6_, phyaddrpointer_reg_7_, phyaddrpointer_reg_8_,
phyaddrpointer_reg_9_, phyaddrpointer_reg_10_, phyaddrpointer_reg_11_,
phyaddrpointer_reg_12_, phyaddrpointer_reg_13_,
phyaddrpointer_reg_14_, phyaddrpointer_reg_15_,
phyaddrpointer_reg_16_, phyaddrpointer_reg_17_,
phyaddrpointer_reg_18_, phyaddrpointer_reg_19_,
phyaddrpointer_reg_20_, phyaddrpointer_reg_21_,
phyaddrpointer_reg_22_, phyaddrpointer_reg_23_,
phyaddrpointer_reg_24_, phyaddrpointer_reg_25_,
phyaddrpointer_reg_26_, phyaddrpointer_reg_27_,
phyaddrpointer_reg_28_, phyaddrpointer_reg_29_,
phyaddrpointer_reg_30_, phyaddrpointer_reg_31_, lword_reg_15_,
lword_reg_14_, lword_reg_13_, lword_reg_12_, lword_reg_11_,
lword_reg_10_, lword_reg_9_, lword_reg_8_, lword_reg_7_, lword_reg_6_,
lword_reg_5_, lword_reg_4_, lword_reg_3_, lword_reg_2_, lword_reg_1_,
lword_reg_0_, uword_reg_14_, uword_reg_13_, uword_reg_12_,
uword_reg_11_, uword_reg_10_, uword_reg_9_, uword_reg_8_,
uword_reg_7_, uword_reg_6_, uword_reg_5_, uword_reg_4_, uword_reg_3_,
uword_reg_2_, uword_reg_1_, uword_reg_0_, datao_reg_0_, datao_reg_1_,
datao_reg_2_, datao_reg_3_, datao_reg_4_, datao_reg_5_, datao_reg_6_,
datao_reg_7_, datao_reg_8_, datao_reg_9_, datao_reg_10_,
datao_reg_11_, datao_reg_12_, datao_reg_13_, datao_reg_14_,
datao_reg_15_, datao_reg_16_, datao_reg_17_, datao_reg_18_,
datao_reg_19_, datao_reg_20_, datao_reg_21_, datao_reg_22_,
datao_reg_23_, datao_reg_24_, datao_reg_25_, datao_reg_26_,
datao_reg_27_, datao_reg_28_, datao_reg_29_, datao_reg_30_,
datao_reg_31_, eax_reg_0_, eax_reg_1_, eax_reg_2_, eax_reg_3_,
eax_reg_4_, eax_reg_5_, eax_reg_6_, eax_reg_7_, eax_reg_8_,
eax_reg_9_, eax_reg_10_, eax_reg_11_, eax_reg_12_, eax_reg_13_,
eax_reg_14_, eax_reg_15_, eax_reg_16_, eax_reg_17_, eax_reg_18_,
eax_reg_19_, eax_reg_20_, eax_reg_21_, eax_reg_22_, eax_reg_23_,
eax_reg_24_, eax_reg_25_, eax_reg_26_, eax_reg_27_, eax_reg_28_,
eax_reg_29_, eax_reg_30_, eax_reg_31_, ebx_reg_0_, ebx_reg_1_,
ebx_reg_2_, ebx_reg_3_, ebx_reg_4_, ebx_reg_5_, ebx_reg_6_,
ebx_reg_7_, ebx_reg_8_, ebx_reg_9_, ebx_reg_10_, ebx_reg_11_,
ebx_reg_12_, ebx_reg_13_, ebx_reg_14_, ebx_reg_15_, ebx_reg_16_,
ebx_reg_17_, ebx_reg_18_, ebx_reg_19_, ebx_reg_20_, ebx_reg_21_,
ebx_reg_22_, ebx_reg_23_, ebx_reg_24_, ebx_reg_25_, ebx_reg_26_,
ebx_reg_27_, ebx_reg_28_, ebx_reg_29_, ebx_reg_30_, ebx_reg_31_,
reip_reg_0_, reip_reg_1_, reip_reg_2_, reip_reg_3_, reip_reg_4_,
reip_reg_5_, reip_reg_6_, reip_reg_7_, reip_reg_8_, reip_reg_9_,
reip_reg_10_, reip_reg_11_, reip_reg_12_, reip_reg_13_, reip_reg_14_,
reip_reg_15_, reip_reg_16_, reip_reg_17_, reip_reg_18_, reip_reg_19_,
reip_reg_20_, reip_reg_21_, reip_reg_22_, reip_reg_23_, reip_reg_24_,
reip_reg_25_, reip_reg_26_, reip_reg_27_, reip_reg_28_, reip_reg_29_,
reip_reg_30_, reip_reg_31_, byteenable_reg_3_, byteenable_reg_2_,
byteenable_reg_1_, byteenable_reg_0_, w_r_n_reg, flush_reg, more_reg,
statebs16_reg, requestpending_reg, d_c_n_reg, m_io_n_reg,
codefetch_reg, ads_n_reg, readrequest_reg, memoryfetch_reg;
output u3445, u3446, u3447, u3448, u3213, u3212, u3211, u3210, u3209, u3208,
u3207, u3206, u3205, u3204, u3203, u3202, u3201, u3200, u3199, u3198,
u3197, u3196, u3195, u3194, u3193, u3192, u3191, u3190, u3189, u3188,
u3187, u3186, u3185, u3184, u3183, u3182, u3181, u3451, u3452, u3180,
u3179, u3178, u3177, u3176, u3175, u3174, u3173, u3172, u3171, u3170,
u3169, u3168, u3167, u3166, u3165, u3164, u3163, u3162, u3161, u3160,
u3159, u3158, u3157, u3156, u3155, u3154, u3153, u3152, u3151, u3453,
u3150, u3149, u3148, u3147, u3146, u3145, u3144, u3143, u3142, u3141,
u3140, u3139, u3138, u3137, u3136, u3135, u3134, u3133, u3132, u3131,
u3130, u3129, u3128, u3127, u3126, u3125, u3124, u3123, u3122, u3121,
u3120, u3119, u3118, u3117, u3116, u3115, u3114, u3113, u3112, u3111,
u3110, u3109, u3108, u3107, u3106, u3105, u3104, u3103, u3102, u3101,
u3100, u3099, u3098, u3097, u3096, u3095, u3094, u3093, u3092, u3091,
u3090, u3089, u3088, u3087, u3086, u3085, u3084, u3083, u3082, u3081,
u3080, u3079, u3078, u3077, u3076, u3075, u3074, u3073, u3072, u3071,
u3070, u3069, u3068, u3067, u3066, u3065, u3064, u3063, u3062, u3061,
u3060, u3059, u3058, u3057, u3056, u3055, u3054, u3053, u3052, u3051,
u3050, u3049, u3048, u3047, u3046, u3045, u3044, u3043, u3042, u3041,
u3040, u3039, u3038, u3037, u3036, u3035, u3034, u3033, u3032, u3031,
u3030, u3029, u3028, u3027, u3026, u3025, u3024, u3023, u3022, u3021,
u3020, u3455, u3456, u3459, u3460, u3461, u3019, u3462, u3463, u3464,
u3465, u3018, u3017, u3016, u3015, u3014, u3013, u3012, u3011, u3010,
u3009, u3008, u3007, u3006, u3005, u3004, u3003, u3002, u3001, u3000,
u2999, u2998, u2997, u2996, u2995, u2994, u2993, u2992, u2991, u2990,
u2989, u2988, u2987, u2986, u2985, u2984, u2983, u2982, u2981, u2980,
u2979, u2978, u2977, u2976, u2975, u2974, u2973, u2972, u2971, u2970,
u2969, u2968, u2967, u2966, u2965, u2964, u2963, u2962, u2961, u2960,
u2959, u2958, u2957, u2956, u2955, u2954, u2953, u2952, u2951, u2950,
u2949, u2948, u2947, u2946, u2945, u2944, u2943, u2942, u2941, u2940,
u2939, u2938, u2937, u2936, u2935, u2934, u2933, u2932, u2931, u2930,
u2929, u2928, u2927, u2926, u2925, u2924, u2923, u2922, u2921, u2920,
u2919, u2918, u2917, u2916, u2915, u2914, u2913, u2912, u2911, u2910,
u2909, u2908, u2907, u2906, u2905, u2904, u2903, u2902, u2901, u2900,
u2899, u2898, u2897, u2896, u2895, u2894, u2893, u2892, u2891, u2890,
u2889, u2888, u2887, u2886, u2885, u2884, u2883, u2882, u2881, u2880,
u2879, u2878, u2877, u2876, u2875, u2874, u2873, u2872, u2871, u2870,
u2869, u2868, u2867, u2866, u2865, u2864, u2863, u2862, u2861, u2860,
u2859, u2858, u2857, u2856, u2855, u2854, u2853, u2852, u2851, u2850,
u2849, u2848, u2847, u2846, u2845, u2844, u2843, u2842, u2841, u2840,
u2839, u2838, u2837, u2836, u2835, u2834, u2833, u2832, u2831, u2830,
u2829, u2828, u2827, u2826, u2825, u2824, u2823, u2822, u2821, u2820,
u2819, u2818, u2817, u2816, u2815, u2814, u2813, u2812, u2811, u2810,
u2809, u2808, u2807, u2806, u2805, u2804, u2803, u2802, u2801, u2800,
u2799, u2798, u2797, u2796, u2795, u3468, u2794, u3469, u3470, u2793,
u3471, u2792, u3472, u2791, u3473, u2790, u2789, u3474, u2788;
wire   n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
n16522, n16523, n16524, n16525, n7819, n7820, n7821, n7822, n7823,
n7824, n7825, n7826, n7827, n7828, n7829, n7831, n7833, n7835, n7837,
n7839, n7841, n7843, n7845, n7847, n7849, n7851, n7853, n7855, n7857,
n7859, n7861, n7863, n7865, n7867, n7869, n7871, n7873, n7875, n7877,
n7879, n7881, n7883, n7885, n7887, n7889, n7891, n7893, n7895, n7897,
n7899, n7901, n7903, n7905, n7907, n7909, n7911, n7913, n7915, n7917,
n7919, n7921, n7923, n7925, n7927, n7929, n7931, n7933, n7935, n7937,
n7939, n7941, n7943, n7945, n7947, n7949, n7951, n7953, n7955, n7957,
n7959, n7961, n7963, n7965, n7967, n7969, n7971, n7973, n7975, n7977,
n7979, n7981, n7983, n7985, n7987, n7989, n7991, n7993, n7995, n7997,
n7999, n8001, n8003, n8005, n8007, n8009, n8011, n8013, n8015, n8017,
n8019, n8021, n8023, n8025, n8027, n8029, n8031, n8033, n8035, n8037,
n8039, n8041, n8043, n8045, n8047, n8049, n8051, n8053, n8055, n8057,
n8059, n8061, n8063, n8065, n8067, n8069, n8071, n8073, n8075, n8077,
n8079, n8081, n8083, n8085, n8087, n8089, n8091, n8093, n8095, n8097,
n8099, n8101, n8103, n8105, n8107, n8109, n8111, n8113, n8115, n8117,
n8119, n8121, n8123, n8125, n8127, n8129, n8131, n8133, n8135, n8137,
n8139, n8141, n8143, n8145, n8147, n8149, n8151, n8153, n8155, n8157,
n8159, n8161, n8163, n8165, n8167, n8169, n8171, n8173, n8175, n8177,
n8179, n8181, n8183, n8185, n8187, n8189, n8191, n8193, n8195, n8197,
n8199, n8201, n8203, n8205, n8207, n8209, n8211, n8213, n8215, n8217,
n8219, n8221, n8223, n8225, n8227, n8229, n8231, n8233, n8235, n8237,
n8239, n8241, n8243, n8245, n8247, n8249, n8251, n8253, n8255, n8257,
n8259, n8261, n8263, n8265, n8267, n8269, n8271, n8273, n8275, n8277,
n8279, n8281, n8283, n8285, n8287, n8289, n8291, n8293, n8295, n8297,
n8299, n8301, n8303, n8305, n8307, n8309, n8311, n8313, n8315, n8317,
n8319, n8321, n8323, n8325, n8327, n8329, n8331, n8333, n8335, n8337,
n8339, n8341, n8343, n8345, n8347, n8349, n8351, n8353, n8355, n8357,
n8359, n8361, n8363, n8365, n8367, n8369, n8371, n8373, n8375, n8377,
n8379, n8381, n8383, n8385, n8387, n8389, n8391, n8393, n8395, n8397,
n8399, n8401, n8403, n8405, n8407, n8409, n8411, n8413, n8415, n8417,
n8419, n8421, n8423, n8425, n8427, n8429, n8431, n8433, n8435, n8437,
n8439, n8441, n8443, n8445, n8447, n8449, n8451, n8453, n8455, n8457,
n8459, n8461, n8463, n8465, n8467, n8469, n8471, n8473, n8475, n8477,
n8479, n8481, n8483, n8485, n8487, n8489, n8491, n8493, n8495, n8497,
n8499, n8501, n8503, n8505, n8507, n8509, n8511, n8513, n8515, n8517,
n8519, n8521, n8523, n8525, n8527, n8529, n8531, n8533, n8535, n8537,
n8539, n8541, n8543, n8545, n8547, n8549, n8551, n8553, n8555, n8557,
n8559, n8561, n8563, n8565, n8567, n8569, n8571, n8573, n8575, n8577,
n8579, n8581, n8583, n8585, n8587, n8589, n8591, n8593, n8595, n8597,
n8599, n8601, n8603, n8605, n8607, n8609, n8611, n8613, n8615, n8617,
n8619, n8621, n8623, n8625, n8627, n8629, n8631, n8633, n8635, n8637,
n8639, n8641, n8643, n8645, n8647, n8649, n8651, n8653, n8655, n8657,
n8659, n8661, n8663, n8665, n8667, n8669, n8671, n8673, n8675, n8677,
n8679, n8681, n8683, n8685, n8687, n8689, n8691, n8693, n8695, n8697,
n8699, n8701, n8703, n8705, n8707, n8709, n8711, n8713, n8715, n8717,
n8719, n8721, n8723, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
n16497;

   and U8268 ( n7819,statebs16_reg,n8790 );
   and U8269 ( n7820,n7821,n12980 );
   not U8270 ( n7821,n8813 );
   buf U8271 ( n7822,n9445 );
   buf U8272 ( n7823,n9457 );
   buf U8273 ( n7824,n9433 );
   buf U8274 ( n7825,n9469 );
   buf U8275 ( n7826,n9421 );
   buf U8276 ( n7827,n9481 );
   buf U8277 ( n7828,n9408 );
   and U8278 ( n7829,n8939,n8940 );
   not U8279 ( u3462,n7829 );
   and U8280 ( n7831,n8925,n8926 );
   not U8281 ( u3463,n7831 );
   and U8282 ( n7833,n8911,n8912 );
   not U8283 ( u3464,n7833 );
   and U8284 ( n7835,n8898,n8899 );
   not U8285 ( u3465,n7835 );
   and U8286 ( n7837,n10922,n10923 );
   not U8287 ( u3018,n7837 );
   and U8288 ( n7839,n10937,n10938 );
   not U8289 ( u3017,n7839 );
   and U8290 ( n7841,n10953,n10954 );
   not U8291 ( u3016,n7841 );
   and U8292 ( n7843,n10983,n10984 );
   not U8293 ( u3015,n7843 );
   and U8294 ( n7845,n11005,n11006 );
   not U8295 ( u3014,n7845 );
   and U8296 ( n7847,n11033,n11034 );
   not U8297 ( u3013,n7847 );
   and U8298 ( n7849,n11052,n11053 );
   not U8299 ( u3012,n7849 );
   and U8300 ( n7851,n11080,n11081 );
   not U8301 ( u3011,n7851 );
   and U8302 ( n7853,n11099,n11100 );
   not U8303 ( u3010,n7853 );
   and U8304 ( n7855,n11126,n11127 );
   not U8305 ( u3009,n7855 );
   and U8306 ( n7857,n11145,n11146 );
   not U8307 ( u3008,n7857 );
   and U8308 ( n7859,n11172,n11173 );
   not U8309 ( u3007,n7859 );
   and U8310 ( n7861,n11191,n11192 );
   not U8311 ( u3006,n7861 );
   and U8312 ( n7863,n11218,n11219 );
   not U8313 ( u3005,n7863 );
   and U8314 ( n7865,n11237,n11238 );
   not U8315 ( u3004,n7865 );
   and U8316 ( n7867,n11264,n11265 );
   not U8317 ( u3003,n7867 );
   and U8318 ( n7869,n11283,n11284 );
   not U8319 ( u3002,n7869 );
   and U8320 ( n7871,n11310,n11311 );
   not U8321 ( u3001,n7871 );
   and U8322 ( n7873,n11329,n11330 );
   not U8323 ( u3000,n7873 );
   and U8324 ( n7875,n11356,n11357 );
   not U8325 ( u2999,n7875 );
   and U8326 ( n7877,n11375,n11376 );
   not U8327 ( u2998,n7877 );
   and U8328 ( n7879,n11404,n11405 );
   not U8329 ( u2997,n7879 );
   and U8330 ( n7881,n11423,n11424 );
   not U8331 ( u2996,n7881 );
   and U8332 ( n7883,n11449,n11450 );
   not U8333 ( u2995,n7883 );
   and U8334 ( n7885,n11468,n11469 );
   not U8335 ( u2994,n7885 );
   and U8336 ( n7887,n11496,n11497 );
   not U8337 ( u2993,n7887 );
   and U8338 ( n7889,n11515,n11516 );
   not U8339 ( u2992,n7889 );
   and U8340 ( n7891,n11542,n11543 );
   not U8341 ( u2991,n7891 );
   and U8342 ( n7893,n11560,n11561 );
   not U8343 ( u2990,n7893 );
   and U8344 ( n7895,n11585,n11586 );
   not U8345 ( u2989,n7895 );
   and U8346 ( n7897,n11598,n11599 );
   not U8347 ( u2988,n7897 );
   and U8348 ( n7899,n11611,n11612 );
   not U8349 ( u2987,n7899 );
   and U8350 ( n7901,n11751,n11752 );
   not U8351 ( u2986,n7901 );
   and U8352 ( n7903,n11765,n11766 );
   not U8353 ( u2985,n7903 );
   and U8354 ( n7905,n11780,n11781 );
   not U8355 ( u2984,n7905 );
   and U8356 ( n7907,n11797,n11798 );
   not U8357 ( u2983,n7907 );
   and U8358 ( n7909,n11818,n11819 );
   not U8359 ( u2982,n7909 );
   and U8360 ( n7911,n11839,n11840 );
   not U8361 ( u2981,n7911 );
   and U8362 ( n7913,n11854,n11855 );
   not U8363 ( u2980,n7913 );
   and U8364 ( n7915,n11869,n11870 );
   not U8365 ( u2979,n7915 );
   and U8366 ( n7917,n11885,n11886 );
   not U8367 ( u2978,n7917 );
   and U8368 ( n7919,n11909,n11910 );
   not U8369 ( u2977,n7919 );
   and U8370 ( n7921,n11924,n11925 );
   not U8371 ( u2976,n7921 );
   and U8372 ( n7923,n11942,n11943 );
   not U8373 ( u2975,n7923 );
   and U8374 ( n7925,n11960,n11961 );
   not U8375 ( u2974,n7925 );
   and U8376 ( n7927,n11980,n11981 );
   not U8377 ( u2973,n7927 );
   and U8378 ( n7929,n11995,n11996 );
   not U8379 ( u2972,n7929 );
   and U8380 ( n7931,n12010,n12011 );
   not U8381 ( u2971,n7931 );
   and U8382 ( n7933,n12025,n12026 );
   not U8383 ( u2970,n7933 );
   and U8384 ( n7935,n12040,n12041 );
   not U8385 ( u2969,n7935 );
   and U8386 ( n7937,n12056,n12057 );
   not U8387 ( u2968,n7937 );
   and U8388 ( n7939,n12070,n12071 );
   not U8389 ( u2967,n7939 );
   and U8390 ( n7941,n12089,n12090 );
   not U8391 ( u2966,n7941 );
   and U8392 ( n7943,n12107,n12108 );
   not U8393 ( u2965,n7943 );
   and U8394 ( n7945,n12124,n12125 );
   not U8395 ( u2964,n7945 );
   and U8396 ( n7947,n12145,n12146 );
   not U8397 ( u2963,n7947 );
   and U8398 ( n7949,n12163,n12164 );
   not U8399 ( u2962,n7949 );
   and U8400 ( n7951,n12180,n12181 );
   not U8401 ( u2961,n7951 );
   and U8402 ( n7953,n12208,n12209 );
   not U8403 ( u2960,n7953 );
   and U8404 ( n7955,n12227,n12228 );
   not U8405 ( u2959,n7955 );
   and U8406 ( n7957,n12243,n12244 );
   not U8407 ( u2958,n7957 );
   and U8408 ( n7959,n12266,n12267 );
   not U8409 ( u2957,n7959 );
   and U8410 ( n7961,n12283,n12284 );
   not U8411 ( u2956,n7961 );
   and U8412 ( n7963,n12302,n12303 );
   not U8413 ( u2955,n7963 );
   and U8414 ( n7965,n12471,n12472 );
   not U8415 ( u2954,n7965 );
   and U8416 ( n7967,n12479,n12480 );
   not U8417 ( u2953,n7967 );
   and U8418 ( n7969,n12484,n12485 );
   not U8419 ( u2952,n7969 );
   and U8420 ( n7971,n12489,n12490 );
   not U8421 ( u2951,n7971 );
   and U8422 ( n7973,n12494,n12495 );
   not U8423 ( u2950,n7973 );
   and U8424 ( n7975,n12499,n12500 );
   not U8425 ( u2949,n7975 );
   and U8426 ( n7977,n12504,n12505 );
   not U8427 ( u2948,n7977 );
   and U8428 ( n7979,n12509,n12510 );
   not U8429 ( u2947,n7979 );
   and U8430 ( n7981,n12514,n12515 );
   not U8431 ( u2946,n7981 );
   and U8432 ( n7983,n12519,n12520 );
   not U8433 ( u2945,n7983 );
   and U8434 ( n7985,n12524,n12525 );
   not U8435 ( u2944,n7985 );
   and U8436 ( n7987,n12529,n12530 );
   not U8437 ( u2943,n7987 );
   and U8438 ( n7989,n12534,n12535 );
   not U8439 ( u2942,n7989 );
   and U8440 ( n7991,n12539,n12540 );
   not U8441 ( u2941,n7991 );
   and U8442 ( n7993,n12544,n12545 );
   not U8443 ( u2940,n7993 );
   and U8444 ( n7995,n12549,n12550 );
   not U8445 ( u2939,n7995 );
   and U8446 ( n7997,n12554,n12555 );
   not U8447 ( u2938,n7997 );
   and U8448 ( n7999,n12559,n12560 );
   not U8449 ( u2937,n7999 );
   and U8450 ( n8001,n12564,n12565 );
   not U8451 ( u2936,n8001 );
   and U8452 ( n8003,n12569,n12570 );
   not U8453 ( u2935,n8003 );
   and U8454 ( n8005,n12574,n12575 );
   not U8455 ( u2934,n8005 );
   and U8456 ( n8007,n12579,n12580 );
   not U8457 ( u2933,n8007 );
   and U8458 ( n8009,n12584,n12585 );
   not U8459 ( u2932,n8009 );
   and U8460 ( n8011,n12589,n12590 );
   not U8461 ( u2931,n8011 );
   and U8462 ( n8013,n12594,n12595 );
   not U8463 ( u2930,n8013 );
   and U8464 ( n8015,n12599,n12600 );
   not U8465 ( u2929,n8015 );
   and U8466 ( n8017,n12604,n12605 );
   not U8467 ( u2928,n8017 );
   and U8468 ( n8019,n12609,n12610 );
   not U8469 ( u2927,n8019 );
   and U8470 ( n8021,n12614,n12615 );
   not U8471 ( u2926,n8021 );
   and U8472 ( n8023,n12619,n12620 );
   not U8473 ( u2925,n8023 );
   and U8474 ( n8025,n12624,n12625 );
   not U8475 ( u2924,n8025 );
   and U8476 ( n8027,n12632,n12633 );
   not U8477 ( u2923,n8027 );
   and U8478 ( n8029,n12640,n12641 );
   not U8479 ( u2922,n8029 );
   and U8480 ( n8031,n12645,n12646 );
   not U8481 ( u2921,n8031 );
   and U8482 ( n8033,n12650,n12651 );
   not U8483 ( u2920,n8033 );
   and U8484 ( n8035,n12655,n12656 );
   not U8485 ( u2919,n8035 );
   and U8486 ( n8037,n12660,n12661 );
   not U8487 ( u2918,n8037 );
   and U8488 ( n8039,n12665,n12666 );
   not U8489 ( u2917,n8039 );
   and U8490 ( n8041,n12670,n12671 );
   not U8491 ( u2916,n8041 );
   and U8492 ( n8043,n12675,n12676 );
   not U8493 ( u2915,n8043 );
   and U8494 ( n8045,n12679,n12680 );
   not U8495 ( u2914,n8045 );
   and U8496 ( n8047,n12684,n12685 );
   not U8497 ( u2913,n8047 );
   and U8498 ( n8049,n12688,n12689 );
   not U8499 ( u2912,n8049 );
   and U8500 ( n8051,n12693,n12694 );
   not U8501 ( u2911,n8051 );
   and U8502 ( n8053,n12698,n12699 );
   not U8503 ( u2910,n8053 );
   and U8504 ( n8055,n12703,n12704 );
   not U8505 ( u2909,n8055 );
   and U8506 ( n8057,n12707,n12708 );
   not U8507 ( u2908,n8057 );
   and U8508 ( n8059,n12711,n12712 );
   not U8509 ( u2907,n8059 );
   and U8510 ( n8061,n12717,n12718 );
   not U8511 ( u2906,n8061 );
   and U8512 ( n8063,n12722,n12723 );
   not U8513 ( u2905,n8063 );
   and U8514 ( n8065,n12727,n12728 );
   not U8515 ( u2904,n8065 );
   and U8516 ( n8067,n12732,n12733 );
   not U8517 ( u2903,n8067 );
   and U8518 ( n8069,n12737,n12738 );
   not U8519 ( u2902,n8069 );
   and U8520 ( n8071,n12742,n12743 );
   not U8521 ( u2901,n8071 );
   and U8522 ( n8073,n12747,n12748 );
   not U8523 ( u2900,n8073 );
   and U8524 ( n8075,n12752,n12753 );
   not U8525 ( u2899,n8075 );
   and U8526 ( n8077,n12757,n12758 );
   not U8527 ( u2898,n8077 );
   and U8528 ( n8079,n12762,n12763 );
   not U8529 ( u2897,n8079 );
   and U8530 ( n8081,n12767,n12768 );
   not U8531 ( u2896,n8081 );
   and U8532 ( n8083,n12772,n12773 );
   not U8533 ( u2895,n8083 );
   and U8534 ( n8085,n12777,n12778 );
   not U8535 ( u2894,n8085 );
   and U8536 ( n8087,n12782,n12783 );
   not U8537 ( u2893,n8087 );
   nand U8538 ( n8089,datao_reg_31_,n12634 );
   not U8539 ( u2892,n8089 );
   and U8540 ( n8091,n12792,n12793 );
   not U8541 ( u2891,n8091 );
   and U8542 ( n8093,n12798,n12799 );
   not U8543 ( u2890,n8093 );
   and U8544 ( n8095,n12802,n12803 );
   not U8545 ( u2889,n8095 );
   and U8546 ( n8097,n12807,n12808 );
   not U8547 ( u2888,n8097 );
   and U8548 ( n8099,n12812,n12813 );
   not U8549 ( u2887,n8099 );
   and U8550 ( n8101,n12817,n12818 );
   not U8551 ( u2886,n8101 );
   and U8552 ( n8103,n12822,n12823 );
   not U8553 ( u2885,n8103 );
   and U8554 ( n8105,n12827,n12828 );
   not U8555 ( u2884,n8105 );
   and U8556 ( n8107,n12832,n12833 );
   not U8557 ( u2883,n8107 );
   and U8558 ( n8109,n12837,n12838 );
   not U8559 ( u2882,n8109 );
   and U8560 ( n8111,n12842,n12843 );
   not U8561 ( u2881,n8111 );
   and U8562 ( n8113,n12847,n12848 );
   not U8563 ( u2880,n8113 );
   and U8564 ( n8115,n12852,n12853 );
   not U8565 ( u2879,n8115 );
   and U8566 ( n8117,n12857,n12858 );
   not U8567 ( u2878,n8117 );
   and U8568 ( n8119,n12862,n12863 );
   not U8569 ( u2877,n8119 );
   and U8570 ( n8121,n12867,n12868 );
   not U8571 ( u2876,n8121 );
   and U8572 ( n8123,n12875,n12876 );
   not U8573 ( u2875,n8123 );
   and U8574 ( n8125,n12884,n12885 );
   not U8575 ( u2874,n8125 );
   and U8576 ( n8127,n12891,n12892 );
   not U8577 ( u2873,n8127 );
   and U8578 ( n8129,n12898,n12899 );
   not U8579 ( u2872,n8129 );
   and U8580 ( n8131,n12905,n12906 );
   not U8581 ( u2871,n8131 );
   and U8582 ( n8133,n12912,n12913 );
   not U8583 ( u2870,n8133 );
   and U8584 ( n8135,n12919,n12920 );
   not U8585 ( u2869,n8135 );
   and U8586 ( n8137,n12926,n12927 );
   not U8587 ( u2868,n8137 );
   and U8588 ( n8139,n12933,n12934 );
   not U8589 ( u2867,n8139 );
   and U8590 ( n8141,n12940,n12941 );
   not U8591 ( u2866,n8141 );
   and U8592 ( n8143,n12947,n12948 );
   not U8593 ( u2865,n8143 );
   and U8594 ( n8145,n12954,n12955 );
   not U8595 ( u2864,n8145 );
   and U8596 ( n8147,n12961,n12962 );
   not U8597 ( u2863,n8147 );
   and U8598 ( n8149,n12968,n12969 );
   not U8599 ( u2862,n8149 );
   and U8600 ( n8151,n12975,n12976 );
   not U8601 ( u2861,n8151 );
   and U8602 ( n8153,n12984,n12985 );
   not U8603 ( u2860,n8153 );
   and U8604 ( n8155,n13004,n13005 );
   not U8605 ( u2859,n8155 );
   and U8606 ( n8157,n13010,n13011 );
   not U8607 ( u2858,n8157 );
   and U8608 ( n8159,n13015,n13016 );
   not U8609 ( u2857,n8159 );
   and U8610 ( n8161,n13020,n13021 );
   not U8611 ( u2856,n8161 );
   and U8612 ( n8163,n13025,n13026 );
   not U8613 ( u2855,n8163 );
   and U8614 ( n8165,n13029,n13030 );
   not U8615 ( u2854,n8165 );
   and U8616 ( n8167,n13034,n13035 );
   not U8617 ( u2853,n8167 );
   and U8618 ( n8169,n13038,n13039 );
   not U8619 ( u2852,n8169 );
   and U8620 ( n8171,n13043,n13044 );
   not U8621 ( u2851,n8171 );
   and U8622 ( n8173,n13047,n13048 );
   not U8623 ( u2850,n8173 );
   and U8624 ( n8175,n13052,n13053 );
   not U8625 ( u2849,n8175 );
   and U8626 ( n8177,n13056,n13057 );
   not U8627 ( u2848,n8177 );
   and U8628 ( n8179,n13061,n13062 );
   not U8629 ( u2847,n8179 );
   and U8630 ( n8181,n13065,n13066 );
   not U8631 ( u2846,n8181 );
   and U8632 ( n8183,n13070,n13071 );
   not U8633 ( u2845,n8183 );
   and U8634 ( n8185,n13074,n13075 );
   not U8635 ( u2844,n8185 );
   and U8636 ( n8187,n13079,n13080 );
   not U8637 ( u2843,n8187 );
   and U8638 ( n8189,n13083,n13084 );
   not U8639 ( u2842,n8189 );
   and U8640 ( n8191,n13088,n13089 );
   not U8641 ( u2841,n8191 );
   and U8642 ( n8193,n13092,n13093 );
   not U8643 ( u2840,n8193 );
   and U8644 ( n8195,n13097,n13098 );
   not U8645 ( u2839,n8195 );
   and U8646 ( n8197,n13101,n13102 );
   not U8647 ( u2838,n8197 );
   and U8648 ( n8199,n13106,n13107 );
   not U8649 ( u2837,n8199 );
   and U8650 ( n8201,n13110,n13111 );
   not U8651 ( u2836,n8201 );
   and U8652 ( n8203,n13115,n13116 );
   not U8653 ( u2835,n8203 );
   and U8654 ( n8205,n13119,n13120 );
   not U8655 ( u2834,n8205 );
   and U8656 ( n8207,n13124,n13125 );
   not U8657 ( u2833,n8207 );
   and U8658 ( n8209,n13128,n13129 );
   not U8659 ( u2832,n8209 );
   and U8660 ( n8211,n13133,n13134 );
   not U8661 ( u2831,n8211 );
   and U8662 ( n8213,n13137,n13138 );
   not U8663 ( u2830,n8213 );
   and U8664 ( n8215,n13142,n13143 );
   not U8665 ( u2829,n8215 );
   and U8666 ( n8217,n13148,n13149 );
   not U8667 ( u2828,n8217 );
   and U8668 ( n8219,n13157,n13158 );
   not U8669 ( u2827,n8219 );
   and U8670 ( n8221,n13184,n13185 );
   not U8671 ( u2826,n8221 );
   and U8672 ( n8223,n13211,n13212 );
   not U8673 ( u2825,n8223 );
   and U8674 ( n8225,n13238,n13239 );
   not U8675 ( u2824,n8225 );
   and U8676 ( n8227,n13267,n13268 );
   not U8677 ( u2823,n8227 );
   and U8678 ( n8229,n13298,n13299 );
   not U8679 ( u2822,n8229 );
   and U8680 ( n8231,n13328,n13329 );
   not U8681 ( u2821,n8231 );
   and U8682 ( n8233,n13354,n13355 );
   not U8683 ( u2820,n8233 );
   and U8684 ( n8235,n13380,n13381 );
   not U8685 ( u2819,n8235 );
   and U8686 ( n8237,n13403,n13404 );
   not U8687 ( u2818,n8237 );
   and U8688 ( n8239,n13426,n13427 );
   not U8689 ( u2817,n8239 );
   and U8690 ( n8241,n13449,n13450 );
   not U8691 ( u2816,n8241 );
   and U8692 ( n8243,n13474,n13475 );
   not U8693 ( u2815,n8243 );
   and U8694 ( n8245,n13498,n13499 );
   not U8695 ( u2814,n8245 );
   and U8696 ( n8247,n13521,n13522 );
   not U8697 ( u2813,n8247 );
   and U8698 ( n8249,n13544,n13545 );
   not U8699 ( u2812,n8249 );
   and U8700 ( n8251,n13571,n13572 );
   not U8701 ( u2811,n8251 );
   and U8702 ( n8253,n13600,n13601 );
   not U8703 ( u2810,n8253 );
   and U8704 ( n8255,n13623,n13624 );
   not U8705 ( u2809,n8255 );
   and U8706 ( n8257,n13648,n13649 );
   not U8707 ( u2808,n8257 );
   and U8708 ( n8259,n13672,n13673 );
   not U8709 ( u2807,n8259 );
   and U8710 ( n8261,n13694,n13695 );
   not U8711 ( u2806,n8261 );
   and U8712 ( n8263,n13716,n13717 );
   not U8713 ( u2805,n8263 );
   and U8714 ( n8265,n13742,n13743 );
   not U8715 ( u2804,n8265 );
   and U8716 ( n8267,n13763,n13764 );
   not U8717 ( u2803,n8267 );
   and U8718 ( n8269,n13792,n13793 );
   not U8719 ( u2802,n8269 );
   and U8720 ( n8271,n13814,n13815 );
   not U8721 ( u2801,n8271 );
   and U8722 ( n8273,n13836,n13837 );
   not U8723 ( u2800,n8273 );
   and U8724 ( n8275,n13863,n13864 );
   not U8725 ( u2799,n8275 );
   and U8726 ( n8277,n13890,n13891 );
   not U8727 ( u2798,n8277 );
   and U8728 ( n8279,n13911,n13912 );
   not U8729 ( u2797,n8279 );
   and U8730 ( n8281,n13968,n13969 );
   not U8731 ( u2796,n8281 );
   and U8732 ( n8283,n16077,n16078 );
   not U8733 ( u2795,n8283 );
   and U8734 ( n8285,n8890,n8891 );
   not U8735 ( u3468,n8285 );
   and U8736 ( n8287,n16082,n16083 );
   not U8737 ( u2794,n8287 );
   and U8738 ( n8289,n8884,n8885 );
   not U8739 ( u3469,n8289 );
   and U8740 ( n8291,n8882,n8883 );
   not U8741 ( u3470,n8291 );
   and U8742 ( n8293,n12470,n16116 );
   not U8743 ( u2793,n8293 );
   and U8744 ( n8295,n8877,n8878 );
   not U8745 ( u3471,n8295 );
   and U8746 ( n8297,n16126,n16127 );
   not U8747 ( u2792,n8297 );
   and U8748 ( n8299,n8850,n8851 );
   not U8749 ( u3472,n8299 );
   and U8750 ( n8301,n16130,n16127 );
   not U8751 ( u2791,n8301 );
   and U8752 ( n8303,n8846,n8847 );
   not U8753 ( u3473,n8303 );
   and U8754 ( n8305,n16133,n16134 );
   not U8755 ( u2790,n8305 );
   and U8756 ( n8307,n9023,n16141 );
   not U8757 ( u2789,n8307 );
   and U8758 ( n8309,n8837,n8838 );
   not U8759 ( u3474,n8309 );
   and U8760 ( n8311,n16144,n16145 );
   not U8761 ( u2788,n8311 );
   and U8762 ( n8313,n8955,n8956 );
   not U8763 ( u3461,n8313 );
   and U8764 ( n8315,n8971,n8972 );
   not U8765 ( u3460,n8315 );
   and U8766 ( n8317,n8984,n8985 );
   not U8767 ( u3459,n8317 );
   and U8768 ( n8319,n8999,n9000 );
   not U8769 ( u3456,n8319 );
   and U8770 ( n8321,n9006,n9007 );
   not U8771 ( u3455,n8321 );
   and U8772 ( n8323,n10812,n10813 );
   not U8773 ( u3020,n8323 );
   and U8774 ( n8325,n10802,n10803 );
   not U8775 ( u3021,n8325 );
   and U8776 ( n8327,n10792,n10793 );
   not U8777 ( u3022,n8327 );
   and U8778 ( n8329,n10782,n10783 );
   not U8779 ( u3023,n8329 );
   and U8780 ( n8331,n10772,n10773 );
   not U8781 ( u3024,n8331 );
   and U8782 ( n8333,n10762,n10763 );
   not U8783 ( u3025,n8333 );
   and U8784 ( n8335,n10752,n10753 );
   not U8785 ( u3026,n8335 );
   and U8786 ( n8337,n10735,n10736 );
   not U8787 ( u3027,n8337 );
   and U8788 ( n8339,n10711,n10712 );
   not U8789 ( u3028,n8339 );
   and U8790 ( n8341,n10702,n10703 );
   not U8791 ( u3029,n8341 );
   and U8792 ( n8343,n10693,n10694 );
   not U8793 ( u3030,n8343 );
   and U8794 ( n8345,n10684,n10685 );
   not U8795 ( u3031,n8345 );
   and U8796 ( n8347,n10675,n10676 );
   not U8797 ( u3032,n8347 );
   and U8798 ( n8349,n10666,n10667 );
   not U8799 ( u3033,n8349 );
   and U8800 ( n8351,n10657,n10658 );
   not U8801 ( u3034,n8351 );
   and U8802 ( n8353,n10643,n10644 );
   not U8803 ( u3035,n8353 );
   and U8804 ( n8355,n10620,n10621 );
   not U8805 ( u3036,n8355 );
   and U8806 ( n8357,n10612,n10613 );
   not U8807 ( u3037,n8357 );
   and U8808 ( n8359,n10604,n10605 );
   not U8809 ( u3038,n8359 );
   and U8810 ( n8361,n10596,n10597 );
   not U8811 ( u3039,n8361 );
   and U8812 ( n8363,n10588,n10589 );
   not U8813 ( u3040,n8363 );
   and U8814 ( n8365,n10580,n10581 );
   not U8815 ( u3041,n8365 );
   and U8816 ( n8367,n10572,n10573 );
   not U8817 ( u3042,n8367 );
   and U8818 ( n8369,n10559,n10560 );
   not U8819 ( u3043,n8369 );
   and U8820 ( n8371,n10532,n10533 );
   not U8821 ( u3044,n8371 );
   and U8822 ( n8373,n10524,n10525 );
   not U8823 ( u3045,n8373 );
   and U8824 ( n8375,n10516,n10517 );
   not U8825 ( u3046,n8375 );
   and U8826 ( n8377,n10508,n10509 );
   not U8827 ( u3047,n8377 );
   and U8828 ( n8379,n10500,n10501 );
   not U8829 ( u3048,n8379 );
   and U8830 ( n8381,n10492,n10493 );
   not U8831 ( u3049,n8381 );
   and U8832 ( n8383,n10484,n10485 );
   not U8833 ( u3050,n8383 );
   and U8834 ( n8385,n10471,n10472 );
   not U8835 ( u3051,n8385 );
   and U8836 ( n8387,n10448,n10449 );
   not U8837 ( u3052,n8387 );
   and U8838 ( n8389,n10440,n10441 );
   not U8839 ( u3053,n8389 );
   and U8840 ( n8391,n10432,n10433 );
   not U8841 ( u3054,n8391 );
   and U8842 ( n8393,n10424,n10425 );
   not U8843 ( u3055,n8393 );
   and U8844 ( n8395,n10416,n10417 );
   not U8845 ( u3056,n8395 );
   and U8846 ( n8397,n10408,n10409 );
   not U8847 ( u3057,n8397 );
   and U8848 ( n8399,n10400,n10401 );
   not U8849 ( u3058,n8399 );
   and U8850 ( n8401,n10387,n10388 );
   not U8851 ( u3059,n8401 );
   and U8852 ( n8403,n10364,n10365 );
   not U8853 ( u3060,n8403 );
   and U8854 ( n8405,n10356,n10357 );
   not U8855 ( u3061,n8405 );
   and U8856 ( n8407,n10348,n10349 );
   not U8857 ( u3062,n8407 );
   and U8858 ( n8409,n10340,n10341 );
   not U8859 ( u3063,n8409 );
   and U8860 ( n8411,n10332,n10333 );
   not U8861 ( u3064,n8411 );
   and U8862 ( n8413,n10324,n10325 );
   not U8863 ( u3065,n8413 );
   and U8864 ( n8415,n10316,n10317 );
   not U8865 ( u3066,n8415 );
   and U8866 ( n8417,n10303,n10304 );
   not U8867 ( u3067,n8417 );
   and U8868 ( n8419,n10278,n10279 );
   not U8869 ( u3068,n8419 );
   and U8870 ( n8421,n10270,n10271 );
   not U8871 ( u3069,n8421 );
   and U8872 ( n8423,n10262,n10263 );
   not U8873 ( u3070,n8423 );
   and U8874 ( n8425,n10254,n10255 );
   not U8875 ( u3071,n8425 );
   and U8876 ( n8427,n10246,n10247 );
   not U8877 ( u3072,n8427 );
   and U8878 ( n8429,n10238,n10239 );
   not U8879 ( u3073,n8429 );
   and U8880 ( n8431,n10230,n10231 );
   not U8881 ( u3074,n8431 );
   and U8882 ( n8433,n10217,n10218 );
   not U8883 ( u3075,n8433 );
   and U8884 ( n8435,n10189,n10190 );
   not U8885 ( u3076,n8435 );
   and U8886 ( n8437,n10181,n10182 );
   not U8887 ( u3077,n8437 );
   and U8888 ( n8439,n10173,n10174 );
   not U8889 ( u3078,n8439 );
   and U8890 ( n8441,n10165,n10166 );
   not U8891 ( u3079,n8441 );
   and U8892 ( n8443,n10157,n10158 );
   not U8893 ( u3080,n8443 );
   and U8894 ( n8445,n10149,n10150 );
   not U8895 ( u3081,n8445 );
   and U8896 ( n8447,n10141,n10142 );
   not U8897 ( u3082,n8447 );
   and U8898 ( n8449,n10129,n10130 );
   not U8899 ( u3083,n8449 );
   and U8900 ( n8451,n10107,n10108 );
   not U8901 ( u3084,n8451 );
   and U8902 ( n8453,n10099,n10100 );
   not U8903 ( u3085,n8453 );
   and U8904 ( n8455,n10091,n10092 );
   not U8905 ( u3086,n8455 );
   and U8906 ( n8457,n10083,n10084 );
   not U8907 ( u3087,n8457 );
   and U8908 ( n8459,n10075,n10076 );
   not U8909 ( u3088,n8459 );
   and U8910 ( n8461,n10067,n10068 );
   not U8911 ( u3089,n8461 );
   and U8912 ( n8463,n10059,n10060 );
   not U8913 ( u3090,n8463 );
   and U8914 ( n8465,n10046,n10047 );
   not U8915 ( u3091,n8465 );
   and U8916 ( n8467,n10024,n10025 );
   not U8917 ( u3092,n8467 );
   and U8918 ( n8469,n10016,n10017 );
   not U8919 ( u3093,n8469 );
   and U8920 ( n8471,n10008,n10009 );
   not U8921 ( u3094,n8471 );
   and U8922 ( n8473,n10000,n10001 );
   not U8923 ( u3095,n8473 );
   and U8924 ( n8475,n9992,n9993 );
   not U8925 ( u3096,n8475 );
   and U8926 ( n8477,n9984,n9985 );
   not U8927 ( u3097,n8477 );
   and U8928 ( n8479,n9976,n9977 );
   not U8929 ( u3098,n8479 );
   and U8930 ( n8481,n9963,n9964 );
   not U8931 ( u3099,n8481 );
   and U8932 ( n8483,n9938,n9939 );
   not U8933 ( u3100,n8483 );
   and U8934 ( n8485,n9930,n9931 );
   not U8935 ( u3101,n8485 );
   and U8936 ( n8487,n9922,n9923 );
   not U8937 ( u3102,n8487 );
   and U8938 ( n8489,n9914,n9915 );
   not U8939 ( u3103,n8489 );
   and U8940 ( n8491,n9906,n9907 );
   not U8941 ( u3104,n8491 );
   and U8942 ( n8493,n9898,n9899 );
   not U8943 ( u3105,n8493 );
   and U8944 ( n8495,n9890,n9891 );
   not U8945 ( u3106,n8495 );
   and U8946 ( n8497,n9877,n9878 );
   not U8947 ( u3107,n8497 );
   and U8948 ( n8499,n9850,n9851 );
   not U8949 ( u3108,n8499 );
   and U8950 ( n8501,n9842,n9843 );
   not U8951 ( u3109,n8501 );
   and U8952 ( n8503,n9834,n9835 );
   not U8953 ( u3110,n8503 );
   and U8954 ( n8505,n9826,n9827 );
   not U8955 ( u3111,n8505 );
   and U8956 ( n8507,n9818,n9819 );
   not U8957 ( u3112,n8507 );
   and U8958 ( n8509,n9810,n9811 );
   not U8959 ( u3113,n8509 );
   and U8960 ( n8511,n9802,n9803 );
   not U8961 ( u3114,n8511 );
   and U8962 ( n8513,n9789,n9790 );
   not U8963 ( u3115,n8513 );
   and U8964 ( n8515,n9760,n9761 );
   not U8965 ( u3116,n8515 );
   and U8966 ( n8517,n9752,n9753 );
   not U8967 ( u3117,n8517 );
   and U8968 ( n8519,n9744,n9745 );
   not U8969 ( u3118,n8519 );
   and U8970 ( n8521,n9736,n9737 );
   not U8971 ( u3119,n8521 );
   and U8972 ( n8523,n9728,n9729 );
   not U8973 ( u3120,n8523 );
   and U8974 ( n8525,n9720,n9721 );
   not U8975 ( u3121,n8525 );
   and U8976 ( n8527,n9712,n9713 );
   not U8977 ( u3122,n8527 );
   and U8978 ( n8529,n9699,n9700 );
   not U8979 ( u3123,n8529 );
   and U8980 ( n8531,n9673,n9674 );
   not U8981 ( u3124,n8531 );
   and U8982 ( n8533,n9665,n9666 );
   not U8983 ( u3125,n8533 );
   and U8984 ( n8535,n9657,n9658 );
   not U8985 ( u3126,n8535 );
   and U8986 ( n8537,n9649,n9650 );
   not U8987 ( u3127,n8537 );
   and U8988 ( n8539,n9641,n9642 );
   not U8989 ( u3128,n8539 );
   and U8990 ( n8541,n9633,n9634 );
   not U8991 ( u3129,n8541 );
   and U8992 ( n8543,n9625,n9626 );
   not U8993 ( u3130,n8543 );
   and U8994 ( n8545,n9612,n9613 );
   not U8995 ( u3131,n8545 );
   and U8996 ( n8547,n9583,n9584 );
   not U8997 ( u3132,n8547 );
   and U8998 ( n8549,n9575,n9576 );
   not U8999 ( u3133,n8549 );
   and U9000 ( n8551,n9567,n9568 );
   not U9001 ( u3134,n8551 );
   and U9002 ( n8553,n9559,n9560 );
   not U9003 ( u3135,n8553 );
   and U9004 ( n8555,n9551,n9552 );
   not U9005 ( u3136,n8555 );
   and U9006 ( n8557,n9543,n9544 );
   not U9007 ( u3137,n8557 );
   and U9008 ( n8559,n9535,n9536 );
   not U9009 ( u3138,n8559 );
   and U9010 ( n8561,n9522,n9523 );
   not U9011 ( u3139,n8561 );
   and U9012 ( n8563,n9483,n9484 );
   not U9013 ( u3140,n8563 );
   and U9014 ( n8565,n9471,n9472 );
   not U9015 ( u3141,n8565 );
   and U9016 ( n8567,n9459,n9460 );
   not U9017 ( u3142,n8567 );
   and U9018 ( n8569,n9447,n9448 );
   not U9019 ( u3143,n8569 );
   and U9020 ( n8571,n9435,n9436 );
   not U9021 ( u3144,n8571 );
   and U9022 ( n8573,n9423,n9424 );
   not U9023 ( u3145,n8573 );
   and U9024 ( n8575,n9411,n9412 );
   not U9025 ( u3146,n8575 );
   and U9026 ( n8577,n9394,n9395 );
   not U9027 ( u3147,n8577 );
   and U9028 ( n8579,n9289,n9290 );
   not U9029 ( u3148,n8579 );
   and U9030 ( n8581,n9278,n9279 );
   not U9031 ( u3149,n8581 );
   and U9032 ( n8583,n9268,n9269 );
   not U9033 ( u3150,n8583 );
   and U9034 ( n8585,n9016,n9017 );
   not U9035 ( u3453,n8585 );
   not U9036 ( n8587,n16525 );
   not U9037 ( u3151,n8587 );
   not U9038 ( n8589,n16524 );
   not U9039 ( u3152,n8589 );
   not U9040 ( n8591,n16523 );
   not U9041 ( u3153,n8591 );
   not U9042 ( n8593,n16522 );
   not U9043 ( u3154,n8593 );
   not U9044 ( n8595,n16521 );
   not U9045 ( u3155,n8595 );
   not U9046 ( n8597,n16520 );
   not U9047 ( u3156,n8597 );
   not U9048 ( n8599,n16519 );
   not U9049 ( u3157,n8599 );
   not U9050 ( n8601,n16518 );
   not U9051 ( u3158,n8601 );
   not U9052 ( n8603,n16517 );
   not U9053 ( u3159,n8603 );
   not U9054 ( n8605,n16516 );
   not U9055 ( u3160,n8605 );
   not U9056 ( n8607,n16515 );
   not U9057 ( u3161,n8607 );
   not U9058 ( n8609,n16514 );
   not U9059 ( u3162,n8609 );
   not U9060 ( n8611,n16513 );
   not U9061 ( u3163,n8611 );
   not U9062 ( n8613,n16512 );
   not U9063 ( u3164,n8613 );
   not U9064 ( n8615,n16511 );
   not U9065 ( u3165,n8615 );
   not U9066 ( n8617,n16510 );
   not U9067 ( u3166,n8617 );
   not U9068 ( n8619,n16509 );
   not U9069 ( u3167,n8619 );
   not U9070 ( n8621,n16508 );
   not U9071 ( u3168,n8621 );
   not U9072 ( n8623,n16507 );
   not U9073 ( u3169,n8623 );
   not U9074 ( n8625,n16506 );
   not U9075 ( u3170,n8625 );
   not U9076 ( n8627,n16505 );
   not U9077 ( u3171,n8627 );
   not U9078 ( n8629,n16504 );
   not U9079 ( u3172,n8629 );
   not U9080 ( n8631,n16503 );
   not U9081 ( u3173,n8631 );
   not U9082 ( n8633,n16502 );
   not U9083 ( u3174,n8633 );
   not U9084 ( n8635,n16501 );
   not U9085 ( u3175,n8635 );
   not U9086 ( n8637,n16500 );
   not U9087 ( u3176,n8637 );
   not U9088 ( n8639,n16499 );
   not U9089 ( u3177,n8639 );
   or U9090 ( n8641,n8756,n9240 );
   not U9091 ( u3178,n8641 );
   or U9092 ( n8643,n9025,n9239 );
   not U9093 ( u3179,n8643 );
   not U9094 ( n8645,n16498 );
   not U9095 ( u3180,n8645 );
   and U9096 ( n8647,n9021,n9022 );
   not U9097 ( u3452,n8647 );
   and U9098 ( n8649,n9028,n9029 );
   not U9099 ( u3451,n8649 );
   and U9100 ( n8651,n9230,n9231 );
   not U9101 ( u3181,n8651 );
   and U9102 ( n8653,n9212,n9213 );
   not U9103 ( u3182,n8653 );
   and U9104 ( n8655,n9193,n9194 );
   not U9105 ( u3183,n8655 );
   and U9106 ( n8657,n9188,n9189 );
   not U9107 ( u3184,n8657 );
   and U9108 ( n8659,n9183,n9184 );
   not U9109 ( u3185,n8659 );
   and U9110 ( n8661,n9178,n9179 );
   not U9111 ( u3186,n8661 );
   and U9112 ( n8663,n9173,n9174 );
   not U9113 ( u3187,n8663 );
   and U9114 ( n8665,n9168,n9169 );
   not U9115 ( u3188,n8665 );
   and U9116 ( n8667,n9163,n9164 );
   not U9117 ( u3189,n8667 );
   and U9118 ( n8669,n9158,n9159 );
   not U9119 ( u3190,n8669 );
   and U9120 ( n8671,n9153,n9154 );
   not U9121 ( u3191,n8671 );
   and U9122 ( n8673,n9148,n9149 );
   not U9123 ( u3192,n8673 );
   and U9124 ( n8675,n9143,n9144 );
   not U9125 ( u3193,n8675 );
   and U9126 ( n8677,n9138,n9139 );
   not U9127 ( u3194,n8677 );
   and U9128 ( n8679,n9133,n9134 );
   not U9129 ( u3195,n8679 );
   and U9130 ( n8681,n9128,n9129 );
   not U9131 ( u3196,n8681 );
   and U9132 ( n8683,n9123,n9124 );
   not U9133 ( u3197,n8683 );
   and U9134 ( n8685,n9118,n9119 );
   not U9135 ( u3198,n8685 );
   and U9136 ( n8687,n9113,n9114 );
   not U9137 ( u3199,n8687 );
   and U9138 ( n8689,n9108,n9109 );
   not U9139 ( u3200,n8689 );
   and U9140 ( n8691,n9103,n9104 );
   not U9141 ( u3201,n8691 );
   and U9142 ( n8693,n9098,n9099 );
   not U9143 ( u3202,n8693 );
   and U9144 ( n8695,n9093,n9094 );
   not U9145 ( u3203,n8695 );
   and U9146 ( n8697,n9088,n9089 );
   not U9147 ( u3204,n8697 );
   and U9148 ( n8699,n9083,n9084 );
   not U9149 ( u3205,n8699 );
   and U9150 ( n8701,n9078,n9079 );
   not U9151 ( u3206,n8701 );
   and U9152 ( n8703,n9073,n9074 );
   not U9153 ( u3207,n8703 );
   and U9154 ( n8705,n9068,n9069 );
   not U9155 ( u3208,n8705 );
   and U9156 ( n8707,n9063,n9064 );
   not U9157 ( u3209,n8707 );
   and U9158 ( n8709,n9058,n9059 );
   not U9159 ( u3210,n8709 );
   and U9160 ( n8711,n9053,n9054 );
   not U9161 ( u3211,n8711 );
   and U9162 ( n8713,n9048,n9049 );
   not U9163 ( u3212,n8713 );
   and U9164 ( n8715,n9040,n9041 );
   not U9165 ( u3213,n8715 );
   and U9166 ( n8717,n9032,n9033 );
   not U9167 ( u3448,n8717 );
   and U9168 ( n8719,n9034,n9035 );
   not U9169 ( u3447,n8719 );
   and U9170 ( n8721,n9036,n9037 );
   not U9171 ( u3446,n8721 );
   and U9172 ( n8723,n9038,n9039 );
   not U9173 ( u3445,n8723 );
   not U9174 ( n8725,n13179 );
   not U9175 ( n8727,n13146 );
   not U9176 ( n8726,n13146 );
   not U9177 ( n8728,n7820 );
   not U9178 ( n8730,n7820 );
   not U9179 ( n8729,n7820 );
   nor U9180 ( n8731,n13006,n11661 );
   not U9181 ( n8732,n8731 );
   not U9182 ( n8734,n8731 );
   not U9183 ( n8733,n8731 );
   nand U9184 ( n8736,n8821,n12787 );
   nand U9185 ( n8735,n8821,n12787 );
   nand U9186 ( n8738,n8868,n8808 );
   nand U9187 ( n8737,n8868,n8808 );
   nand U9188 ( n8740,n8789,n10934 );
   nand U9189 ( n8739,n8789,n10934 );
   nand U9190 ( n8742,state_reg_1_,n9202 );
   nand U9191 ( n8741,state_reg_1_,n9202 );
   nand U9192 ( n8744,n8849,n9208 );
   nand U9193 ( n8743,n8849,n9208 );
   not U9194 ( n8745,n8782 );
   not U9195 ( n8747,n8782 );
   not U9196 ( n8746,n13168 );
   nand U9197 ( n8749,state_reg_2_,n8849 );
   nand U9198 ( n8748,state_reg_2_,n8849 );
   nand U9199 ( n8750,n11706,n11707 );
   not U9200 ( n8751,n8750 );
   not U9201 ( n8754,n8750 );
   not U9202 ( n8752,n8750 );
   not U9203 ( n8753,n8750 );
   not U9204 ( n8756,n9023 );
   not U9205 ( n8755,n9023 );
   and U9206 ( n8757,n10788,n10808 );
   not U9207 ( n8758,n8757 );
   not U9208 ( n8761,n8757 );
   not U9209 ( n8759,n8757 );
   not U9210 ( n8760,n8757 );
   and U9211 ( n8762,n8871,n10838 );
   not U9212 ( n8763,n8762 );
   not U9213 ( n8766,n8762 );
   not U9214 ( n8764,n8762 );
   not U9215 ( n8765,n8762 );
   buf U9216 ( n8767,n9517 );
   buf U9217 ( n8768,n9410 );
   buf U9218 ( n8769,n9404 );
   buf U9219 ( n8770,n9422 );
   buf U9220 ( n8771,n9418 );
   buf U9221 ( n8772,n9434 );
   buf U9222 ( n8773,n9430 );
   not U9223 ( n8774,n13959 );
   not U9224 ( n8775,n10972 );
   buf U9225 ( n8776,n9446 );
   buf U9226 ( n8777,n9442 );
   buf U9227 ( n8778,n12880 );
   not U9228 ( n8779,n10927 );
   buf U9229 ( n8780,n9458 );
   buf U9230 ( n8781,n9454 );
   buf U9231 ( n8782,n13168 );
   buf U9232 ( n8783,n12797 );
   not U9233 ( n8784,n8811 );
   buf U9234 ( n8785,n12476 );
   buf U9235 ( n8786,n9470 );
   buf U9236 ( n8787,n9466 );
   buf U9237 ( n8788,n11755 );
   not U9238 ( n8790,state2_reg_2_ );
   not U9239 ( n8789,state2_reg_2_ );
   buf U9240 ( n8791,n12716 );
   not U9241 ( n8792,n10949 );
   buf U9242 ( n8793,n9482 );
   buf U9243 ( n8794,n9478 );
   not U9244 ( n8795,n12787 );
   not U9245 ( n8796,n12454 );
   buf U9246 ( n8797,n13006 );
   not U9247 ( n8798,n13164 );
   buf U9248 ( n8799,n12473 );
   nand U9249 ( n8800,n11619,n8961 );
   nand U9250 ( n8802,n11661,state2_reg_2_ );
   nand U9251 ( n8801,n11661,state2_reg_2_ );
   not U9252 ( n8803,n7819 );
   not U9253 ( n8805,n7819 );
   not U9254 ( n8804,n7819 );
   and U9255 ( n8806,n12467,n12468 );
   not U9256 ( n8807,n8806 );
   not U9257 ( n8810,n8806 );
   not U9258 ( n8808,n8806 );
   not U9259 ( n8809,n8806 );
   buf U9260 ( n8811,n14090 );
   buf U9261 ( n8812,n10927 );
   buf U9262 ( n8813,n12794 );
   buf U9263 ( n8814,n9519 );
   buf U9264 ( n8815,n9512 );
   not U9265 ( n8816,n10934 );
   buf U9266 ( n8817,n10980 );
   not U9267 ( n8818,n16012 );
   not U9268 ( n8819,n13314 );
   not U9269 ( n8820,n11764 );
   not U9270 ( n8821,state2_reg_0_ );
   not U9271 ( n8822,n13183 );
   buf U9272 ( n8823,n12064 );
   buf U9273 ( n8824,n13177 );
   nand U9274 ( n8826,n13958,n12461 );
   nand U9275 ( n8825,n13958,n12461 );
   nand U9276 ( n8828,n12462,n12463 );
   nand U9277 ( n8827,n12462,n12463 );
   not U9278 ( n8829,n8763 );
   not U9279 ( n8831,n8766 );
   not U9280 ( n8830,n8766 );
   nand U9281 ( n8832,n12629,n12630 );
   not U9282 ( n8833,n8832 );
   not U9283 ( n8836,n8832 );
   not U9284 ( n8834,n8832 );
   not U9285 ( n8835,n8832 );
   nand U9286 ( n8838,n8839,readrequest_reg );
   nand U9287 ( n8837,n8840,n8841 );
   not U9288 ( n8841,n8839 );
   nor U9289 ( n8839,n8842,n8843 );
   nand U9290 ( n8840,n8844,state2_reg_2_ );
   nor U9291 ( n8844,n8845,n8757 );
   nand U9292 ( n8847,m_io_n_reg,n8742 );
   nand U9293 ( n8846,memoryfetch_reg,n8849 );
   or U9294 ( n8851,n8852,n8853 );
   nand U9295 ( n8850,n8854,n8852 );
   nand U9296 ( n8852,n8855,n8856 );
   nor U9297 ( n8856,n8857,n8858 );
   nor U9298 ( n8855,n8842,n8859 );
   nor U9299 ( n8859,n8860,n8861 );
   nand U9300 ( n8861,n8862,n8821 );
   nand U9301 ( n8854,n8864,n8865 );
   nand U9302 ( n8865,n8866,n8867 );
   nor U9303 ( n8864,n8868,n8869 );
   nor U9304 ( n8869,n8870,n8863 );
   nor U9305 ( n8870,n8790,n8872 );
   nand U9306 ( n8872,n8873,n8862 );
   nand U9307 ( n8873,n8874,n8875 );
   nand U9308 ( n8875,statebs16_reg,n8876 );
   nand U9309 ( n8878,n8879,n8880 );
   nand U9310 ( n8877,more_reg,n8881 );
   or U9311 ( n8883,n8741,readrequest_reg );
   nand U9312 ( n8882,w_r_n_reg,n8742 );
   nor U9313 ( n8884,n8886,n8887 );
   nor U9314 ( n8887,n8888,n8889 );
   and U9315 ( n8886,n8888,byteenable_reg_0_ );
   nand U9316 ( n8891,n8892,reip_reg_0_ );
   nor U9317 ( n8890,n8893,n8894 );
   nor U9318 ( n8894,n8888,n8895 );
   nand U9319 ( n8895,n8896,n8897 );
   nand U9320 ( n8897,reip_reg_0_,datawidth_reg_0_ );
   nor U9321 ( n8896,reip_reg_1_,datawidth_reg_1_ );
   and U9322 ( n8893,n8888,byteenable_reg_2_ );
   nand U9323 ( n8899,n8900,instqueuewr_addr_reg_0_ );
   nand U9324 ( n8898,n8901,n8902 );
   nand U9325 ( n8901,n8903,n8904 );
   nand U9326 ( n8904,n8857,n8905 );
   nor U9327 ( n8903,n8906,n8907 );
   nor U9328 ( n8907,n8860,n8908 );
   nor U9329 ( n8906,n8909,n8910 );
   nand U9330 ( n8912,n8900,instqueuewr_addr_reg_1_ );
   nand U9331 ( n8911,n8913,n8902 );
   nand U9332 ( n8913,n8914,n8915 );
   nand U9333 ( n8915,n8916,n8917 );
   nor U9334 ( n8914,n8918,n8919 );
   nor U9335 ( n8919,n8909,n8920 );
   nor U9336 ( n8918,n8921,n8922 );
   nor U9337 ( n8921,n8923,n8924 );
   nand U9338 ( n8926,n8900,instqueuewr_addr_reg_2_ );
   nand U9339 ( n8925,n8927,n8902 );
   nand U9340 ( n8927,n8928,n8929 );
   nand U9341 ( n8929,n8916,n8930 );
   nor U9342 ( n8928,n8931,n8932 );
   nor U9343 ( n8932,n8909,n8933 );
   nor U9344 ( n8931,n8922,n8934 );
   nand U9345 ( n8934,n8935,n8936 );
   or U9346 ( n8935,n8937,n8938 );
   nand U9347 ( n8940,n8900,instqueuewr_addr_reg_3_ );
   nand U9348 ( n8939,n8941,n8902 );
   nand U9349 ( n8941,n8942,n8943 );
   nand U9350 ( n8943,n8944,n8916 );
   nor U9351 ( n8942,n8945,n8946 );
   nor U9352 ( n8946,n8909,n8947 );
   nor U9353 ( n8909,n8948,state2_reg_3_ );
   nor U9354 ( n8945,n8949,n8922 );
   nor U9355 ( n8949,n8950,n8951 );
   not U9356 ( n8951,n8952 );
   nor U9357 ( n8950,n8953,n8954 );
   nand U9358 ( n8956,instqueuerd_addr_reg_0_,n8957 );
   nand U9359 ( n8957,n8958,n8959 );
   nand U9360 ( n8959,n8960,n8961 );
   nand U9361 ( n8955,n8962,n8958 );
   nand U9362 ( n8962,n8963,n8964 );
   nand U9363 ( n8964,state2_reg_1_,n8965 );
   nor U9364 ( n8963,n8966,n8967 );
   and U9365 ( n8967,n8968,n8969 );
   and U9366 ( n8966,n8970,n8960 );
   nand U9367 ( n8972,n8973,instqueuerd_addr_reg_1_ );
   nand U9368 ( n8971,n8974,n8958 );
   nand U9369 ( n8974,n8975,n8976 );
   nand U9370 ( n8976,n8969,n8977 );
   nor U9371 ( n8975,n8978,n8979 );
   nor U9372 ( n8979,n8980,n8981 );
   nor U9373 ( n8978,n8965,n8982 );
   nand U9374 ( n8982,state2_reg_1_,n8983 );
   nand U9375 ( n8985,n8973,instqueuerd_addr_reg_2_ );
   nand U9376 ( n8984,n8986,n8958 );
   nand U9377 ( n8986,n8987,n8988 );
   nand U9378 ( n8988,n8969,n8989 );
   nor U9379 ( n8987,n8990,n8991 );
   nor U9380 ( n8991,n8992,n8981 );
   nor U9381 ( n8990,n8983,n8993 );
   nand U9382 ( n8993,instaddrpointer_reg_0_,state2_reg_1_ );
   nand U9383 ( n8983,n8994,n8995 );
   nand U9384 ( n8995,n8996,n8997 );
   nand U9385 ( n8994,instaddrpointer_reg_31_,n8998 );
   nand U9386 ( n9000,n8973,instqueuerd_addr_reg_3_ );
   nand U9387 ( n8999,n9001,n8958 );
   nand U9388 ( n9001,n9002,n9003 );
   nand U9389 ( n9003,n8960,n9004 );
   nand U9390 ( n9002,n8969,n9005 );
   nand U9391 ( n9007,n9008,n8958 );
   nor U9392 ( n9008,n8981,n9009 );
   nand U9393 ( n9006,n8973,instqueuerd_addr_reg_4_ );
   not U9394 ( n8973,n8958 );
   nand U9395 ( n8958,n9010,n9011 );
   nand U9396 ( n9011,state2_reg_3_,n8821 );
   nor U9397 ( n9010,n9012,n9013 );
   nor U9398 ( n9013,n9014,n9015 );
   or U9399 ( n9017,n9018,n9019 );
   nand U9400 ( n9016,n9019,n9020 );
   nand U9401 ( n9022,n9023,datawidth_reg_1_ );
   nand U9402 ( n9021,n9024,n8756 );
   nand U9403 ( n9024,n9026,n9027 );
   nand U9404 ( n9029,n9030,n9025 );
   nor U9405 ( n9030,bs16_n,n9031 );
   nand U9406 ( n9028,n9023,datawidth_reg_0_ );
   nand U9407 ( n9033,be_n_reg_0_,n8848 );
   nand U9408 ( n9032,byteenable_reg_0_,n8849 );
   nand U9409 ( n9035,be_n_reg_1_,n8742 );
   nand U9410 ( n9034,byteenable_reg_1_,n8849 );
   nand U9411 ( n9037,be_n_reg_2_,n8848 );
   nand U9412 ( n9036,byteenable_reg_2_,n8849 );
   nand U9413 ( n9039,be_n_reg_3_,n8742 );
   nand U9414 ( n9038,byteenable_reg_3_,n8849 );
   nand U9415 ( n9041,address_reg_29_,n8741 );
   nor U9416 ( n9040,n9042,n9043 );
   nor U9417 ( n9043,n8743,n9045 );
   nor U9418 ( n9042,n8749,n9047 );
   nand U9419 ( n9049,address_reg_28_,n8848 );
   nor U9420 ( n9048,n9050,n9051 );
   nor U9421 ( n9051,n9047,n8744 );
   nor U9422 ( n9050,n8748,n9052 );
   nand U9423 ( n9054,address_reg_27_,n8848 );
   nor U9424 ( n9053,n9055,n9056 );
   nor U9425 ( n9056,n8744,n9052 );
   nor U9426 ( n9055,n8748,n9057 );
   nand U9427 ( n9059,address_reg_26_,n8741 );
   nor U9428 ( n9058,n9060,n9061 );
   nor U9429 ( n9061,n9044,n9057 );
   nor U9430 ( n9060,n9046,n9062 );
   nand U9431 ( n9064,address_reg_25_,n8741 );
   nor U9432 ( n9063,n9065,n9066 );
   nor U9433 ( n9066,n8743,n9062 );
   nor U9434 ( n9065,n8748,n9067 );
   nand U9435 ( n9069,address_reg_24_,n8742 );
   nor U9436 ( n9068,n9070,n9071 );
   nor U9437 ( n9071,n8744,n9067 );
   nor U9438 ( n9070,n8749,n9072 );
   nand U9439 ( n9074,address_reg_23_,n8741 );
   nor U9440 ( n9073,n9075,n9076 );
   nor U9441 ( n9076,n9044,n9072 );
   nor U9442 ( n9075,n9046,n9077 );
   nand U9443 ( n9079,address_reg_22_,n8741 );
   nor U9444 ( n9078,n9080,n9081 );
   nor U9445 ( n9081,n9044,n9077 );
   nor U9446 ( n9080,n8748,n9082 );
   nand U9447 ( n9084,address_reg_21_,n8848 );
   nor U9448 ( n9083,n9085,n9086 );
   nor U9449 ( n9086,n8743,n9082 );
   nor U9450 ( n9085,n8749,n9087 );
   nand U9451 ( n9089,address_reg_20_,n8848 );
   nor U9452 ( n9088,n9090,n9091 );
   nor U9453 ( n9091,n8744,n9087 );
   nor U9454 ( n9090,n9046,n9092 );
   nand U9455 ( n9094,address_reg_19_,n8741 );
   nor U9456 ( n9093,n9095,n9096 );
   nor U9457 ( n9096,n9044,n9092 );
   nor U9458 ( n9095,n8748,n9097 );
   nand U9459 ( n9099,address_reg_18_,n8742 );
   nor U9460 ( n9098,n9100,n9101 );
   nor U9461 ( n9101,n8743,n9097 );
   nor U9462 ( n9100,n8749,n9102 );
   nand U9463 ( n9104,address_reg_17_,n8848 );
   nor U9464 ( n9103,n9105,n9106 );
   nor U9465 ( n9106,n8744,n9102 );
   nor U9466 ( n9105,n8748,n9107 );
   nand U9467 ( n9109,address_reg_16_,n8741 );
   nor U9468 ( n9108,n9110,n9111 );
   nor U9469 ( n9111,n9044,n9107 );
   nor U9470 ( n9110,n9046,n9112 );
   nand U9471 ( n9114,address_reg_15_,n8742 );
   nor U9472 ( n9113,n9115,n9116 );
   nor U9473 ( n9116,n8743,n9112 );
   nor U9474 ( n9115,n8748,n9117 );
   nand U9475 ( n9119,address_reg_14_,n8848 );
   nor U9476 ( n9118,n9120,n9121 );
   nor U9477 ( n9121,n8744,n9117 );
   nor U9478 ( n9120,n8749,n9122 );
   nand U9479 ( n9124,address_reg_13_,n8741 );
   nor U9480 ( n9123,n9125,n9126 );
   nor U9481 ( n9126,n8743,n9122 );
   nor U9482 ( n9125,n9046,n9127 );
   nand U9483 ( n9129,address_reg_12_,n8742 );
   nor U9484 ( n9128,n9130,n9131 );
   nor U9485 ( n9131,n9044,n9127 );
   nor U9486 ( n9130,n9046,n9132 );
   nand U9487 ( n9134,address_reg_11_,n8848 );
   nor U9488 ( n9133,n9135,n9136 );
   nor U9489 ( n9136,n9044,n9132 );
   nor U9490 ( n9135,n8749,n9137 );
   nand U9491 ( n9139,address_reg_10_,n8741 );
   nor U9492 ( n9138,n9140,n9141 );
   nor U9493 ( n9141,n8743,n9137 );
   nor U9494 ( n9140,n8748,n9142 );
   nand U9495 ( n9144,address_reg_9_,n8848 );
   nor U9496 ( n9143,n9145,n9146 );
   nor U9497 ( n9146,n8744,n9142 );
   nor U9498 ( n9145,n9046,n9147 );
   nand U9499 ( n9149,address_reg_8_,n8848 );
   nor U9500 ( n9148,n9150,n9151 );
   nor U9501 ( n9151,n9044,n9147 );
   nor U9502 ( n9150,n8749,n9152 );
   nand U9503 ( n9154,address_reg_7_,n8848 );
   nor U9504 ( n9153,n9155,n9156 );
   nor U9505 ( n9156,n8743,n9152 );
   nor U9506 ( n9155,n9046,n9157 );
   nand U9507 ( n9159,address_reg_6_,n8741 );
   nor U9508 ( n9158,n9160,n9161 );
   nor U9509 ( n9161,n8744,n9157 );
   nor U9510 ( n9160,n8748,n9162 );
   nand U9511 ( n9164,address_reg_5_,n8742 );
   nor U9512 ( n9163,n9165,n9166 );
   nor U9513 ( n9166,n9044,n9162 );
   nor U9514 ( n9165,n9046,n9167 );
   nand U9515 ( n9169,address_reg_4_,n8742 );
   nor U9516 ( n9168,n9170,n9171 );
   nor U9517 ( n9171,n8743,n9167 );
   nor U9518 ( n9170,n8749,n9172 );
   nand U9519 ( n9174,address_reg_3_,n8741 );
   nor U9520 ( n9173,n9175,n9176 );
   nor U9521 ( n9176,n8744,n9172 );
   nor U9522 ( n9175,n8748,n9177 );
   nand U9523 ( n9179,address_reg_2_,n8741 );
   nor U9524 ( n9178,n9180,n9181 );
   nor U9525 ( n9181,n9044,n9177 );
   nor U9526 ( n9180,n9046,n9182 );
   nand U9527 ( n9184,address_reg_1_,n8742 );
   nor U9528 ( n9183,n9185,n9186 );
   nor U9529 ( n9186,n8743,n9182 );
   nor U9530 ( n9185,n8749,n9187 );
   nand U9531 ( n9189,address_reg_0_,n8742 );
   nor U9532 ( n9188,n9190,n9191 );
   nor U9533 ( n9191,n8744,n9187 );
   nor U9534 ( n9190,n9192,n8748 );
   nand U9535 ( n9194,n9195,n9196 );
   nor U9536 ( n9196,n9197,n9198 );
   nor U9537 ( n9198,requestpending_reg,hold );
   nor U9538 ( n9197,n9199,n9200 );
   nor U9539 ( n9199,requestpending_reg,n9027 );
   nor U9540 ( n9195,n9201,n9202 );
   nor U9541 ( n9201,n9203,n9204 );
   nor U9542 ( n9193,n9205,n9206 );
   nor U9543 ( n9206,n9207,n9208 );
   nor U9544 ( n9207,n9200,n9209 );
   nand U9545 ( n9209,n9210,n9211 );
   nand U9546 ( n9211,n9204,n9202 );
   not U9547 ( n9204,na_n );
   nand U9548 ( n9210,hold,state_reg_0_ );
   nor U9549 ( n9200,n9203,n8862 );
   not U9550 ( n9205,n8749 );
   nand U9551 ( n9046,state_reg_2_,n8849 );
   nor U9552 ( n9213,n9214,n9215 );
   nand U9553 ( n9215,n9216,n8743 );
   nand U9554 ( n9044,n8849,n9208 );
   not U9555 ( n8849,n8742 );
   nand U9556 ( n9216,n9217,state_reg_1_ );
   nor U9557 ( n9217,n9218,n9219 );
   nor U9558 ( n9219,hold,n9220 );
   nand U9559 ( n9220,n8862,n8853 );
   nor U9560 ( n9218,n9221,n9208 );
   nor U9561 ( n9221,n9222,n9202 );
   and U9562 ( n9222,n8862,hold );
   nor U9563 ( n9214,n9027,n9223 );
   nand U9564 ( n9223,state_reg_0_,requestpending_reg );
   nor U9565 ( n9212,n9224,n9225 );
   nor U9566 ( n9225,n8848,n8862 );
   nor U9567 ( n9224,n9226,n9208 );
   nor U9568 ( n9226,n9227,n9228 );
   and U9569 ( n9227,n9203,n9229 );
   nand U9570 ( n9231,n9228,na_n );
   nor U9571 ( n9230,n9232,n9233 );
   nor U9572 ( n9233,state_reg_2_,n9234 );
   nor U9573 ( n9234,n9202,n9235 );
   nand U9574 ( n9235,requestpending_reg,n9236 );
   nand U9575 ( n9236,ready_n,state_reg_1_ );
   nor U9576 ( n9232,n9229,n9237 );
   nand U9577 ( n9237,n8848,n9027 );
   nor U9578 ( n9229,n8853,hold );
   not U9579 ( n8853,requestpending_reg );
   nor U9580 ( n16498,n8755,n9238 );
   nor U9581 ( n16499,n8755,n9241 );
   nor U9582 ( n16500,n9025,n9242 );
   nor U9583 ( n16501,n8756,n9243 );
   nor U9584 ( n16502,n8756,n9244 );
   nor U9585 ( n16503,n8755,n9245 );
   nor U9586 ( n16504,n9025,n9246 );
   nor U9587 ( n16505,n8756,n9247 );
   nor U9588 ( n16506,n8755,n9248 );
   nor U9589 ( n16507,n9025,n9249 );
   nor U9590 ( n16508,n8755,n9250 );
   nor U9591 ( n16509,n9025,n9251 );
   nor U9592 ( n16510,n9025,n9252 );
   nor U9593 ( n16511,n8755,n9253 );
   nor U9594 ( n16512,n8756,n9254 );
   nor U9595 ( n16513,n9025,n9255 );
   nor U9596 ( n16514,n8755,n9256 );
   nor U9597 ( n16515,n8756,n9257 );
   nor U9598 ( n16516,n8755,n9258 );
   nor U9599 ( n16517,n9025,n9259 );
   nor U9600 ( n16518,n8756,n9260 );
   nor U9601 ( n16519,n8755,n9261 );
   nor U9602 ( n16520,n9025,n9262 );
   nor U9603 ( n16521,n8756,n9263 );
   nor U9604 ( n16522,n8755,n9264 );
   nor U9605 ( n16523,n9025,n9265 );
   nor U9606 ( n16524,n8756,n9266 );
   nor U9607 ( n16525,n8756,n9267 );
   nor U9608 ( n9269,n9270,n9271 );
   nor U9609 ( n9271,n8863,n9272 );
   or U9610 ( n9272,n9273,ready_n );
   nor U9611 ( n9270,state2_reg_0_,n9274 );
   nand U9612 ( n9274,statebs16_reg,state2_reg_1_ );
   nor U9613 ( n9268,n9275,n9276 );
   nor U9614 ( n9276,n9019,n8789 );
   nor U9615 ( n9019,n8863,n9277 );
   nand U9616 ( n9279,state2_reg_1_,n9280 );
   nand U9617 ( n9280,n9281,n9282 );
   nor U9618 ( n9278,n9283,n9284 );
   nor U9619 ( n9284,n9277,n9285 );
   nor U9620 ( n9285,n9286,n9287 );
   nor U9621 ( n9286,ready_n,n9288 );
   nor U9622 ( n9290,n9291,n9292 );
   nand U9623 ( n9292,n9282,n9293 );
   nand U9624 ( n9282,n9294,ready_n );
   nor U9625 ( n9294,state2_reg_2_,n8863 );
   nor U9626 ( n9291,n9295,n8908 );
   nor U9627 ( n9289,n9296,n9297 );
   nand U9628 ( n9297,n9298,n9299 );
   nand U9629 ( n9299,n9300,n8821 );
   nor U9630 ( n9300,n9277,n9301 );
   and U9631 ( n9301,n8969,n8868 );
   nand U9632 ( n9298,n9277,state2_reg_0_ );
   not U9633 ( n9277,n9281 );
   nand U9634 ( n9281,n9302,n9303 );
   nor U9635 ( n9303,n9304,n9305 );
   nor U9636 ( n9305,state2_reg_0_,n9306 );
   nor U9637 ( n9306,n8948,n8862 );
   nor U9638 ( n9304,n9307,n8863 );
   nor U9639 ( n9307,state2_reg_1_,n9308 );
   nor U9640 ( n9302,n9309,n8790 );
   nor U9641 ( n9309,n9310,n9311 );
   and U9642 ( n9296,n9308,n9287 );
   nand U9643 ( n9308,n9312,n9313 );
   nor U9644 ( n9313,n9314,n9315 );
   nand U9645 ( n9315,n9316,n9317 );
   nand U9646 ( n9317,n9318,n9319 );
   nand U9647 ( n9319,n9320,instqueuewr_addr_reg_3_ );
   nor U9648 ( n9318,instqueuewr_addr_reg_4_,n9321 );
   nor U9649 ( n9321,n9322,n9323 );
   nand U9650 ( n9323,n9324,n9325 );
   nand U9651 ( n9325,n9326,n9327 );
   nor U9652 ( n9326,instqueuewr_addr_reg_2_,n9328 );
   nand U9653 ( n9324,n9329,n9330 );
   nand U9654 ( n9330,n9331,n9332 );
   nand U9655 ( n9332,n9333,n9334 );
   nand U9656 ( n9333,n9335,instqueuewr_addr_reg_0_ );
   nor U9657 ( n9335,n9336,n9337 );
   nor U9658 ( n9337,n9014,n8980 );
   not U9659 ( n8980,n9338 );
   nor U9660 ( n9336,n9339,n9340 );
   nor U9661 ( n9331,n9341,n9342 );
   nor U9662 ( n9342,n9014,n9343 );
   nor U9663 ( n9343,n9344,n8970 );
   nand U9664 ( n8970,n9345,n9346 );
   nand U9665 ( n9346,n9347,n8968 );
   nand U9666 ( n9345,n9348,n9349 );
   nor U9667 ( n9344,n8968,n9350 );
   nor U9668 ( n9341,n8968,n9340 );
   nor U9669 ( n9329,n9351,n9352 );
   nor U9670 ( n9352,n9353,n9354 );
   nor U9671 ( n9353,n9355,n9328 );
   not U9672 ( n9355,n9327 );
   nor U9673 ( n9351,n9356,n9357 );
   nand U9674 ( n9357,n9358,n9359 );
   nand U9675 ( n9359,n9014,instqueuerd_addr_reg_1_ );
   nand U9676 ( n9358,n9338,n9340 );
   nand U9677 ( n9338,n9360,n9361 );
   nand U9678 ( n9361,n8961,n9339 );
   nor U9679 ( n9360,n9362,n9363 );
   nor U9680 ( n9363,n9364,n8920 );
   and U9681 ( n9362,n9347,n8977 );
   nand U9682 ( n9347,n9365,n9366 );
   nand U9683 ( n9366,n9367,n8845 );
   nor U9684 ( n9322,instqueuewr_addr_reg_3_,n9320 );
   not U9685 ( n9320,n9368 );
   nand U9686 ( n9316,n9369,n9370 );
   or U9687 ( n9370,more_reg,flush_reg );
   not U9688 ( n9314,n9371 );
   nor U9689 ( n9312,n8880,n9372 );
   nand U9690 ( n9372,n9373,n9374 );
   nand U9691 ( n9374,n9375,n9376 );
   nand U9692 ( n8880,n9377,n9378 );
   nand U9693 ( n9378,n9379,n9380 );
   nor U9694 ( n9377,n9381,n9382 );
   nor U9695 ( n9382,n9383,n9384 );
   nor U9696 ( n9383,n9385,n9386 );
   nand U9697 ( n9386,n9387,n9350 );
   nand U9698 ( n9385,n9388,n9371 );
   nand U9699 ( n9371,n9389,n9390 );
   nor U9700 ( n9389,n9391,n9392 );
   nor U9701 ( n9381,n9393,n9365 );
   nor U9702 ( n9395,n9396,n9397 );
   nand U9703 ( n9397,n9398,n9399 );
   nand U9704 ( n9399,n9400,n9401 );
   nand U9705 ( n9398,instqueue_reg_15__7_,n9402 );
   nor U9706 ( n9396,n9403,n8769 );
   nor U9707 ( n9394,n9405,n9406 );
   nor U9708 ( n9406,n9407,n7828 );
   nor U9709 ( n9405,n9409,n8768 );
   nor U9710 ( n9412,n9413,n9414 );
   nand U9711 ( n9414,n9415,n9416 );
   nand U9712 ( n9416,n9417,n9401 );
   nand U9713 ( n9415,instqueue_reg_15__6_,n9402 );
   nor U9714 ( n9413,n9403,n8771 );
   nor U9715 ( n9411,n9419,n9420 );
   nor U9716 ( n9420,n9407,n7826 );
   nor U9717 ( n9419,n9409,n8770 );
   nor U9718 ( n9424,n9425,n9426 );
   nand U9719 ( n9426,n9427,n9428 );
   nand U9720 ( n9428,n9429,n9401 );
   nand U9721 ( n9427,instqueue_reg_15__5_,n9402 );
   nor U9722 ( n9425,n9403,n8773 );
   nor U9723 ( n9423,n9431,n9432 );
   nor U9724 ( n9432,n9407,n7824 );
   nor U9725 ( n9431,n9409,n8772 );
   nor U9726 ( n9436,n9437,n9438 );
   nand U9727 ( n9438,n9439,n9440 );
   nand U9728 ( n9440,n9441,n9401 );
   nand U9729 ( n9439,instqueue_reg_15__4_,n9402 );
   nor U9730 ( n9437,n9403,n8777 );
   nor U9731 ( n9435,n9443,n9444 );
   nor U9732 ( n9444,n9407,n7822 );
   nor U9733 ( n9443,n9409,n8776 );
   nor U9734 ( n9448,n9449,n9450 );
   nand U9735 ( n9450,n9451,n9452 );
   nand U9736 ( n9452,n9453,n9401 );
   nand U9737 ( n9451,instqueue_reg_15__3_,n9402 );
   nor U9738 ( n9449,n9403,n8781 );
   nor U9739 ( n9447,n9455,n9456 );
   nor U9740 ( n9456,n9407,n7823 );
   nor U9741 ( n9455,n9409,n8780 );
   nor U9742 ( n9460,n9461,n9462 );
   nand U9743 ( n9462,n9463,n9464 );
   nand U9744 ( n9464,n9465,n9401 );
   nand U9745 ( n9463,instqueue_reg_15__2_,n9402 );
   nor U9746 ( n9461,n9403,n8787 );
   nor U9747 ( n9459,n9467,n9468 );
   nor U9748 ( n9468,n9407,n7825 );
   nor U9749 ( n9467,n9409,n8786 );
   nor U9750 ( n9472,n9473,n9474 );
   nand U9751 ( n9474,n9475,n9476 );
   nand U9752 ( n9476,n9477,n9401 );
   nand U9753 ( n9475,instqueue_reg_15__1_,n9402 );
   nor U9754 ( n9473,n9403,n8794 );
   nor U9755 ( n9471,n9479,n9480 );
   nor U9756 ( n9480,n9407,n7827 );
   nor U9757 ( n9479,n9409,n8793 );
   nor U9758 ( n9484,n9485,n9486 );
   nand U9759 ( n9486,n9487,n9488 );
   nand U9760 ( n9488,n9489,n9401 );
   nand U9761 ( n9401,n9490,n9491 );
   nand U9762 ( n9491,state2_reg_2_,n9492 );
   nand U9763 ( n9490,n9493,n9494 );
   nand U9764 ( n9487,instqueue_reg_15__0_,n9402 );
   nand U9765 ( n9402,n9495,n9496 );
   nand U9766 ( n9496,state2_reg_3_,n9409 );
   nor U9767 ( n9495,n9497,n9498 );
   nor U9768 ( n9498,n9499,n9500 );
   nand U9769 ( n9500,n9501,n9502 );
   nand U9770 ( n9501,n9503,n9504 );
   nand U9771 ( n9504,n9407,n9403 );
   and U9772 ( n9499,n9494,n9505 );
   nand U9773 ( n9494,n9409,n9506 );
   nand U9774 ( n9506,n9507,n9508 );
   nor U9775 ( n9497,n8790,n9492 );
   nand U9776 ( n9492,n9409,n9509 );
   nand U9777 ( n9509,n9510,n9511 );
   nor U9778 ( n9485,n9403,n8815 );
   nand U9779 ( n9403,n9513,n9514 );
   nor U9780 ( n9483,n9515,n9516 );
   nor U9781 ( n9516,n9407,n8767 );
   nand U9782 ( n9407,n8953,n9518 );
   nor U9783 ( n9515,n9409,n8814 );
   nand U9784 ( n9409,n9520,n9521 );
   nor U9785 ( n9523,n9524,n9525 );
   nand U9786 ( n9525,n9526,n9527 );
   nand U9787 ( n9527,n9400,n9528 );
   nand U9788 ( n9526,instqueue_reg_14__7_,n9529 );
   nor U9789 ( n9524,n9404,n9530 );
   nor U9790 ( n9522,n9531,n9532 );
   nor U9791 ( n9532,n7828,n9533 );
   nor U9792 ( n9531,n8768,n9534 );
   nor U9793 ( n9536,n9537,n9538 );
   nand U9794 ( n9538,n9539,n9540 );
   nand U9795 ( n9540,n9417,n9528 );
   nand U9796 ( n9539,instqueue_reg_14__6_,n9529 );
   nor U9797 ( n9537,n9418,n9530 );
   nor U9798 ( n9535,n9541,n9542 );
   nor U9799 ( n9542,n7826,n9533 );
   nor U9800 ( n9541,n8770,n9534 );
   nor U9801 ( n9544,n9545,n9546 );
   nand U9802 ( n9546,n9547,n9548 );
   nand U9803 ( n9548,n9429,n9528 );
   nand U9804 ( n9547,instqueue_reg_14__5_,n9529 );
   nor U9805 ( n9545,n9430,n9530 );
   nor U9806 ( n9543,n9549,n9550 );
   nor U9807 ( n9550,n7824,n9533 );
   nor U9808 ( n9549,n8772,n9534 );
   nor U9809 ( n9552,n9553,n9554 );
   nand U9810 ( n9554,n9555,n9556 );
   nand U9811 ( n9556,n9441,n9528 );
   nand U9812 ( n9555,instqueue_reg_14__4_,n9529 );
   nor U9813 ( n9553,n9442,n9530 );
   nor U9814 ( n9551,n9557,n9558 );
   nor U9815 ( n9558,n7822,n9533 );
   nor U9816 ( n9557,n8776,n9534 );
   nor U9817 ( n9560,n9561,n9562 );
   nand U9818 ( n9562,n9563,n9564 );
   nand U9819 ( n9564,n9453,n9528 );
   nand U9820 ( n9563,instqueue_reg_14__3_,n9529 );
   nor U9821 ( n9561,n9454,n9530 );
   nor U9822 ( n9559,n9565,n9566 );
   nor U9823 ( n9566,n7823,n9533 );
   nor U9824 ( n9565,n8780,n9534 );
   nor U9825 ( n9568,n9569,n9570 );
   nand U9826 ( n9570,n9571,n9572 );
   nand U9827 ( n9572,n9465,n9528 );
   nand U9828 ( n9571,instqueue_reg_14__2_,n9529 );
   nor U9829 ( n9569,n9466,n9530 );
   nor U9830 ( n9567,n9573,n9574 );
   nor U9831 ( n9574,n7825,n9533 );
   nor U9832 ( n9573,n8786,n9534 );
   nor U9833 ( n9576,n9577,n9578 );
   nand U9834 ( n9578,n9579,n9580 );
   nand U9835 ( n9580,n9477,n9528 );
   nand U9836 ( n9579,instqueue_reg_14__1_,n9529 );
   nor U9837 ( n9577,n9478,n9530 );
   nor U9838 ( n9575,n9581,n9582 );
   nor U9839 ( n9582,n7827,n9533 );
   nor U9840 ( n9581,n8793,n9534 );
   nor U9841 ( n9584,n9585,n9586 );
   nand U9842 ( n9586,n9587,n9588 );
   nand U9843 ( n9588,n9489,n9528 );
   nand U9844 ( n9528,n9589,n9590 );
   nand U9845 ( n9590,n9591,n9511 );
   nand U9846 ( n9589,n9592,n9493 );
   not U9847 ( n9592,n9593 );
   nand U9848 ( n9587,instqueue_reg_14__0_,n9529 );
   nand U9849 ( n9529,n9594,n9595 );
   nand U9850 ( n9595,state2_reg_3_,n9534 );
   nor U9851 ( n9594,n9596,n9597 );
   nor U9852 ( n9597,n9598,n9599 );
   nand U9853 ( n9599,n9600,n9502 );
   nand U9854 ( n9600,n9503,n9601 );
   nand U9855 ( n9601,n9533,n9530 );
   nor U9856 ( n9598,n9593,n9602 );
   nand U9857 ( n9593,n9507,n9603 );
   nor U9858 ( n9596,n9604,n8871 );
   nor U9859 ( n9604,n9605,n9606 );
   nor U9860 ( n9585,n9512,n9530 );
   nand U9861 ( n9530,n9607,n9513 );
   nor U9862 ( n9583,n9608,n9609 );
   nor U9863 ( n9609,n8767,n9533 );
   nand U9864 ( n9533,n8923,n9610 );
   nor U9865 ( n9608,n8814,n9534 );
   nand U9866 ( n9534,n9611,n9520 );
   nor U9867 ( n9613,n9614,n9615 );
   nand U9868 ( n9615,n9616,n9617 );
   nand U9869 ( n9617,n9400,n9618 );
   nand U9870 ( n9616,instqueue_reg_13__7_,n9619 );
   nor U9871 ( n9614,n9404,n9620 );
   nor U9872 ( n9612,n9621,n9622 );
   nor U9873 ( n9622,n7828,n9623 );
   nor U9874 ( n9621,n8768,n9624 );
   nor U9875 ( n9626,n9627,n9628 );
   nand U9876 ( n9628,n9629,n9630 );
   nand U9877 ( n9630,n9417,n9618 );
   nand U9878 ( n9629,instqueue_reg_13__6_,n9619 );
   nor U9879 ( n9627,n9418,n9620 );
   nor U9880 ( n9625,n9631,n9632 );
   nor U9881 ( n9632,n7826,n9623 );
   nor U9882 ( n9631,n8770,n9624 );
   nor U9883 ( n9634,n9635,n9636 );
   nand U9884 ( n9636,n9637,n9638 );
   nand U9885 ( n9638,n9429,n9618 );
   nand U9886 ( n9637,instqueue_reg_13__5_,n9619 );
   nor U9887 ( n9635,n9430,n9620 );
   nor U9888 ( n9633,n9639,n9640 );
   nor U9889 ( n9640,n7824,n9623 );
   nor U9890 ( n9639,n8772,n9624 );
   nor U9891 ( n9642,n9643,n9644 );
   nand U9892 ( n9644,n9645,n9646 );
   nand U9893 ( n9646,n9441,n9618 );
   nand U9894 ( n9645,instqueue_reg_13__4_,n9619 );
   nor U9895 ( n9643,n9442,n9620 );
   nor U9896 ( n9641,n9647,n9648 );
   nor U9897 ( n9648,n7822,n9623 );
   nor U9898 ( n9647,n8776,n9624 );
   nor U9899 ( n9650,n9651,n9652 );
   nand U9900 ( n9652,n9653,n9654 );
   nand U9901 ( n9654,n9453,n9618 );
   nand U9902 ( n9653,instqueue_reg_13__3_,n9619 );
   nor U9903 ( n9651,n9454,n9620 );
   nor U9904 ( n9649,n9655,n9656 );
   nor U9905 ( n9656,n7823,n9623 );
   nor U9906 ( n9655,n8780,n9624 );
   nor U9907 ( n9658,n9659,n9660 );
   nand U9908 ( n9660,n9661,n9662 );
   nand U9909 ( n9662,n9465,n9618 );
   nand U9910 ( n9661,instqueue_reg_13__2_,n9619 );
   nor U9911 ( n9659,n9466,n9620 );
   nor U9912 ( n9657,n9663,n9664 );
   nor U9913 ( n9664,n7825,n9623 );
   nor U9914 ( n9663,n8786,n9624 );
   nor U9915 ( n9666,n9667,n9668 );
   nand U9916 ( n9668,n9669,n9670 );
   nand U9917 ( n9670,n9477,n9618 );
   nand U9918 ( n9669,instqueue_reg_13__1_,n9619 );
   nor U9919 ( n9667,n9478,n9620 );
   nor U9920 ( n9665,n9671,n9672 );
   nor U9921 ( n9672,n7827,n9623 );
   nor U9922 ( n9671,n8793,n9624 );
   nor U9923 ( n9674,n9675,n9676 );
   nand U9924 ( n9676,n9677,n9678 );
   nand U9925 ( n9678,n9489,n9618 );
   nand U9926 ( n9618,n9679,n9680 );
   nand U9927 ( n9680,state2_reg_2_,n9681 );
   nand U9928 ( n9679,n9682,n9493 );
   nand U9929 ( n9677,instqueue_reg_13__0_,n9619 );
   nand U9930 ( n9619,n9683,n9684 );
   nand U9931 ( n9684,state2_reg_3_,n9624 );
   nor U9932 ( n9683,n9685,n9686 );
   nor U9933 ( n9686,n9687,n9688 );
   nand U9934 ( n9688,n9689,n9502 );
   nand U9935 ( n9689,n9503,n9690 );
   nand U9936 ( n9690,n9623,n9620 );
   and U9937 ( n9687,n9682,n9505 );
   nand U9938 ( n9682,n9624,n9691 );
   nand U9939 ( n9691,n9692,n9507 );
   nor U9940 ( n9685,n8871,n9681 );
   nand U9941 ( n9681,n9624,n9693 );
   nand U9942 ( n9693,n9694,n9510 );
   nor U9943 ( n9675,n9512,n9620 );
   nand U9944 ( n9620,n9695,n9513 );
   nor U9945 ( n9673,n9696,n9697 );
   nor U9946 ( n9697,n8767,n9623 );
   nand U9947 ( n9623,n8924,n9610 );
   nor U9948 ( n9696,n8814,n9624 );
   nand U9949 ( n9624,n9698,n9520 );
   nor U9950 ( n9700,n9701,n9702 );
   nand U9951 ( n9702,n9703,n9704 );
   nand U9952 ( n9704,n9400,n9705 );
   nand U9953 ( n9703,instqueue_reg_12__7_,n9706 );
   nor U9954 ( n9701,n9404,n9707 );
   nor U9955 ( n9699,n9708,n9709 );
   nor U9956 ( n9709,n9408,n9710 );
   nor U9957 ( n9708,n9410,n9711 );
   nor U9958 ( n9713,n9714,n9715 );
   nand U9959 ( n9715,n9716,n9717 );
   nand U9960 ( n9717,n9417,n9705 );
   nand U9961 ( n9716,instqueue_reg_12__6_,n9706 );
   nor U9962 ( n9714,n9418,n9707 );
   nor U9963 ( n9712,n9718,n9719 );
   nor U9964 ( n9719,n9421,n9710 );
   nor U9965 ( n9718,n9422,n9711 );
   nor U9966 ( n9721,n9722,n9723 );
   nand U9967 ( n9723,n9724,n9725 );
   nand U9968 ( n9725,n9429,n9705 );
   nand U9969 ( n9724,instqueue_reg_12__5_,n9706 );
   nor U9970 ( n9722,n9430,n9707 );
   nor U9971 ( n9720,n9726,n9727 );
   nor U9972 ( n9727,n9433,n9710 );
   nor U9973 ( n9726,n9434,n9711 );
   nor U9974 ( n9729,n9730,n9731 );
   nand U9975 ( n9731,n9732,n9733 );
   nand U9976 ( n9733,n9441,n9705 );
   nand U9977 ( n9732,instqueue_reg_12__4_,n9706 );
   nor U9978 ( n9730,n9442,n9707 );
   nor U9979 ( n9728,n9734,n9735 );
   nor U9980 ( n9735,n9445,n9710 );
   nor U9981 ( n9734,n9446,n9711 );
   nor U9982 ( n9737,n9738,n9739 );
   nand U9983 ( n9739,n9740,n9741 );
   nand U9984 ( n9741,n9453,n9705 );
   nand U9985 ( n9740,instqueue_reg_12__3_,n9706 );
   nor U9986 ( n9738,n9454,n9707 );
   nor U9987 ( n9736,n9742,n9743 );
   nor U9988 ( n9743,n9457,n9710 );
   nor U9989 ( n9742,n9458,n9711 );
   nor U9990 ( n9745,n9746,n9747 );
   nand U9991 ( n9747,n9748,n9749 );
   nand U9992 ( n9749,n9465,n9705 );
   nand U9993 ( n9748,instqueue_reg_12__2_,n9706 );
   nor U9994 ( n9746,n9466,n9707 );
   nor U9995 ( n9744,n9750,n9751 );
   nor U9996 ( n9751,n9469,n9710 );
   nor U9997 ( n9750,n9470,n9711 );
   nor U9998 ( n9753,n9754,n9755 );
   nand U9999 ( n9755,n9756,n9757 );
   nand U10000 ( n9757,n9477,n9705 );
   nand U10001 ( n9756,instqueue_reg_12__1_,n9706 );
   nor U10002 ( n9754,n9478,n9707 );
   nor U10003 ( n9752,n9758,n9759 );
   nor U10004 ( n9759,n9481,n9710 );
   nor U10005 ( n9758,n9482,n9711 );
   nor U10006 ( n9761,n9762,n9763 );
   nand U10007 ( n9763,n9764,n9765 );
   nand U10008 ( n9765,n9489,n9705 );
   nand U10009 ( n9705,n9766,n9767 );
   nand U10010 ( n9767,n9694,n9591 );
   nand U10011 ( n9766,n9768,n9493 );
   nand U10012 ( n9764,instqueue_reg_12__0_,n9706 );
   nand U10013 ( n9706,n9769,n9770 );
   nand U10014 ( n9770,state2_reg_3_,n9711 );
   nor U10015 ( n9769,n9771,n9772 );
   nor U10016 ( n9772,n9773,n9774 );
   and U10017 ( n9774,n9768,n9505 );
   nand U10018 ( n9768,n9711,n9775 );
   nand U10019 ( n9775,n9507,n8920 );
   nor U10020 ( n9507,n8947,n8933 );
   nor U10021 ( n9773,n9776,n9777 );
   and U10022 ( n9776,n9707,n9710 );
   nor U10023 ( n9771,n9778,n8789 );
   nor U10024 ( n9778,n9605,n9779 );
   nor U10025 ( n9762,n9512,n9707 );
   nand U10026 ( n9707,n9780,n9513 );
   nor U10027 ( n9513,n9781,n9782 );
   nor U10028 ( n9760,n9783,n9784 );
   nor U10029 ( n9784,n9517,n9710 );
   nand U10030 ( n9710,n9785,n9610 );
   nor U10031 ( n9610,n9786,n8954 );
   nor U10032 ( n9783,n9519,n9711 );
   nand U10033 ( n9711,n9787,n9520 );
   nor U10034 ( n9520,n9354,n9788 );
   nor U10035 ( n9790,n9791,n9792 );
   nand U10036 ( n9792,n9793,n9794 );
   nand U10037 ( n9794,n9400,n9795 );
   nand U10038 ( n9793,instqueue_reg_11__7_,n9796 );
   nor U10039 ( n9791,n9404,n9797 );
   nor U10040 ( n9789,n9798,n9799 );
   nor U10041 ( n9799,n9408,n9800 );
   nor U10042 ( n9798,n9410,n9801 );
   nor U10043 ( n9803,n9804,n9805 );
   nand U10044 ( n9805,n9806,n9807 );
   nand U10045 ( n9807,n9417,n9795 );
   nand U10046 ( n9806,instqueue_reg_11__6_,n9796 );
   nor U10047 ( n9804,n9418,n9797 );
   nor U10048 ( n9802,n9808,n9809 );
   nor U10049 ( n9809,n9421,n9800 );
   nor U10050 ( n9808,n9422,n9801 );
   nor U10051 ( n9811,n9812,n9813 );
   nand U10052 ( n9813,n9814,n9815 );
   nand U10053 ( n9815,n9429,n9795 );
   nand U10054 ( n9814,instqueue_reg_11__5_,n9796 );
   nor U10055 ( n9812,n9430,n9797 );
   nor U10056 ( n9810,n9816,n9817 );
   nor U10057 ( n9817,n9433,n9800 );
   nor U10058 ( n9816,n9434,n9801 );
   nor U10059 ( n9819,n9820,n9821 );
   nand U10060 ( n9821,n9822,n9823 );
   nand U10061 ( n9823,n9441,n9795 );
   nand U10062 ( n9822,instqueue_reg_11__4_,n9796 );
   nor U10063 ( n9820,n9442,n9797 );
   nor U10064 ( n9818,n9824,n9825 );
   nor U10065 ( n9825,n9445,n9800 );
   nor U10066 ( n9824,n9446,n9801 );
   nor U10067 ( n9827,n9828,n9829 );
   nand U10068 ( n9829,n9830,n9831 );
   nand U10069 ( n9831,n9453,n9795 );
   nand U10070 ( n9830,instqueue_reg_11__3_,n9796 );
   nor U10071 ( n9828,n9454,n9797 );
   nor U10072 ( n9826,n9832,n9833 );
   nor U10073 ( n9833,n9457,n9800 );
   nor U10074 ( n9832,n9458,n9801 );
   nor U10075 ( n9835,n9836,n9837 );
   nand U10076 ( n9837,n9838,n9839 );
   nand U10077 ( n9839,n9465,n9795 );
   nand U10078 ( n9838,instqueue_reg_11__2_,n9796 );
   nor U10079 ( n9836,n9466,n9797 );
   nor U10080 ( n9834,n9840,n9841 );
   nor U10081 ( n9841,n9469,n9800 );
   nor U10082 ( n9840,n9470,n9801 );
   nor U10083 ( n9843,n9844,n9845 );
   nand U10084 ( n9845,n9846,n9847 );
   nand U10085 ( n9847,n9477,n9795 );
   nand U10086 ( n9846,instqueue_reg_11__1_,n9796 );
   nor U10087 ( n9844,n9478,n9797 );
   nor U10088 ( n9842,n9848,n9849 );
   nor U10089 ( n9849,n9481,n9800 );
   nor U10090 ( n9848,n9482,n9801 );
   nor U10091 ( n9851,n9852,n9853 );
   nand U10092 ( n9853,n9854,n9855 );
   nand U10093 ( n9855,n9489,n9795 );
   nand U10094 ( n9795,n9856,n9857 );
   nand U10095 ( n9857,state2_reg_2_,n9858 );
   nand U10096 ( n9856,n9859,n9493 );
   nand U10097 ( n9854,instqueue_reg_11__0_,n9796 );
   nand U10098 ( n9796,n9860,n9861 );
   nand U10099 ( n9861,state2_reg_3_,n9801 );
   nor U10100 ( n9860,n9862,n9863 );
   nor U10101 ( n9863,n9864,n9865 );
   nand U10102 ( n9865,n9866,n9502 );
   nand U10103 ( n9866,n9503,n9867 );
   nand U10104 ( n9867,n9800,n9797 );
   and U10105 ( n9864,n9859,n9505 );
   nand U10106 ( n9859,n9801,n9868 );
   nand U10107 ( n9868,n9869,n9508 );
   nor U10108 ( n9862,n8789,n9858 );
   nand U10109 ( n9858,n9801,n9870 );
   nand U10110 ( n9870,n9871,n9511 );
   nor U10111 ( n9852,n9512,n9797 );
   nand U10112 ( n9797,n9872,n9514 );
   nor U10113 ( n9850,n9873,n9874 );
   nor U10114 ( n9874,n9517,n9800 );
   nand U10115 ( n9800,n9875,n8938 );
   nor U10116 ( n9873,n9519,n9801 );
   nand U10117 ( n9801,n9876,n9521 );
   nor U10118 ( n9878,n9879,n9880 );
   nand U10119 ( n9880,n9881,n9882 );
   nand U10120 ( n9882,n9400,n9883 );
   nand U10121 ( n9881,instqueue_reg_10__7_,n9884 );
   nor U10122 ( n9879,n9404,n9885 );
   nor U10123 ( n9877,n9886,n9887 );
   nor U10124 ( n9887,n9408,n9888 );
   nor U10125 ( n9886,n9410,n9889 );
   nor U10126 ( n9891,n9892,n9893 );
   nand U10127 ( n9893,n9894,n9895 );
   nand U10128 ( n9895,n9417,n9883 );
   nand U10129 ( n9894,instqueue_reg_10__6_,n9884 );
   nor U10130 ( n9892,n9418,n9885 );
   nor U10131 ( n9890,n9896,n9897 );
   nor U10132 ( n9897,n9421,n9888 );
   nor U10133 ( n9896,n9422,n9889 );
   nor U10134 ( n9899,n9900,n9901 );
   nand U10135 ( n9901,n9902,n9903 );
   nand U10136 ( n9903,n9429,n9883 );
   nand U10137 ( n9902,instqueue_reg_10__5_,n9884 );
   nor U10138 ( n9900,n9430,n9885 );
   nor U10139 ( n9898,n9904,n9905 );
   nor U10140 ( n9905,n9433,n9888 );
   nor U10141 ( n9904,n9434,n9889 );
   nor U10142 ( n9907,n9908,n9909 );
   nand U10143 ( n9909,n9910,n9911 );
   nand U10144 ( n9911,n9441,n9883 );
   nand U10145 ( n9910,instqueue_reg_10__4_,n9884 );
   nor U10146 ( n9908,n9442,n9885 );
   nor U10147 ( n9906,n9912,n9913 );
   nor U10148 ( n9913,n9445,n9888 );
   nor U10149 ( n9912,n9446,n9889 );
   nor U10150 ( n9915,n9916,n9917 );
   nand U10151 ( n9917,n9918,n9919 );
   nand U10152 ( n9919,n9453,n9883 );
   nand U10153 ( n9918,instqueue_reg_10__3_,n9884 );
   nor U10154 ( n9916,n9454,n9885 );
   nor U10155 ( n9914,n9920,n9921 );
   nor U10156 ( n9921,n9457,n9888 );
   nor U10157 ( n9920,n9458,n9889 );
   nor U10158 ( n9923,n9924,n9925 );
   nand U10159 ( n9925,n9926,n9927 );
   nand U10160 ( n9927,n9465,n9883 );
   nand U10161 ( n9926,instqueue_reg_10__2_,n9884 );
   nor U10162 ( n9924,n9466,n9885 );
   nor U10163 ( n9922,n9928,n9929 );
   nor U10164 ( n9929,n9469,n9888 );
   nor U10165 ( n9928,n9470,n9889 );
   nor U10166 ( n9931,n9932,n9933 );
   nand U10167 ( n9933,n9934,n9935 );
   nand U10168 ( n9935,n9477,n9883 );
   nand U10169 ( n9934,instqueue_reg_10__1_,n9884 );
   nor U10170 ( n9932,n9478,n9885 );
   nor U10171 ( n9930,n9936,n9937 );
   nor U10172 ( n9937,n9481,n9888 );
   nor U10173 ( n9936,n9482,n9889 );
   nor U10174 ( n9939,n9940,n9941 );
   nand U10175 ( n9941,n9942,n9943 );
   nand U10176 ( n9943,n9489,n9883 );
   nand U10177 ( n9883,n9944,n9945 );
   nand U10178 ( n9945,n9946,n9511 );
   not U10179 ( n9511,n9606 );
   nand U10180 ( n9944,n9947,n9493 );
   not U10181 ( n9947,n9948 );
   nand U10182 ( n9942,instqueue_reg_10__0_,n9884 );
   nand U10183 ( n9884,n9949,n9950 );
   nand U10184 ( n9950,state2_reg_3_,n9889 );
   nor U10185 ( n9949,n9951,n9952 );
   nor U10186 ( n9952,n9953,n9954 );
   nand U10187 ( n9954,n9955,n9502 );
   nand U10188 ( n9955,n9503,n9956 );
   nand U10189 ( n9956,n9888,n9885 );
   nor U10190 ( n9953,n9948,n9602 );
   nand U10191 ( n9948,n9869,n9603 );
   nor U10192 ( n9951,n9957,n8871 );
   nor U10193 ( n9957,n9606,n9958 );
   nand U10194 ( n9606,n9959,n9960 );
   nor U10195 ( n9940,n9512,n9885 );
   nand U10196 ( n9885,n9872,n9607 );
   nor U10197 ( n9938,n9961,n9962 );
   nor U10198 ( n9962,n9517,n9888 );
   nand U10199 ( n9888,n9875,n8923 );
   nor U10200 ( n9961,n9519,n9889 );
   nand U10201 ( n9889,n9876,n9611 );
   nor U10202 ( n9964,n9965,n9966 );
   nand U10203 ( n9966,n9967,n9968 );
   nand U10204 ( n9968,n9400,n9969 );
   nand U10205 ( n9967,instqueue_reg_9__7_,n9970 );
   nor U10206 ( n9965,n9404,n9971 );
   nor U10207 ( n9963,n9972,n9973 );
   nor U10208 ( n9973,n7828,n9974 );
   nor U10209 ( n9972,n8768,n9975 );
   nor U10210 ( n9977,n9978,n9979 );
   nand U10211 ( n9979,n9980,n9981 );
   nand U10212 ( n9981,n9417,n9969 );
   nand U10213 ( n9980,instqueue_reg_9__6_,n9970 );
   nor U10214 ( n9978,n9418,n9971 );
   nor U10215 ( n9976,n9982,n9983 );
   nor U10216 ( n9983,n7826,n9974 );
   nor U10217 ( n9982,n8770,n9975 );
   nor U10218 ( n9985,n9986,n9987 );
   nand U10219 ( n9987,n9988,n9989 );
   nand U10220 ( n9989,n9429,n9969 );
   nand U10221 ( n9988,instqueue_reg_9__5_,n9970 );
   nor U10222 ( n9986,n9430,n9971 );
   nor U10223 ( n9984,n9990,n9991 );
   nor U10224 ( n9991,n7824,n9974 );
   nor U10225 ( n9990,n8772,n9975 );
   nor U10226 ( n9993,n9994,n9995 );
   nand U10227 ( n9995,n9996,n9997 );
   nand U10228 ( n9997,n9441,n9969 );
   nand U10229 ( n9996,instqueue_reg_9__4_,n9970 );
   nor U10230 ( n9994,n9442,n9971 );
   nor U10231 ( n9992,n9998,n9999 );
   nor U10232 ( n9999,n7822,n9974 );
   nor U10233 ( n9998,n8776,n9975 );
   nor U10234 ( n10001,n10002,n10003 );
   nand U10235 ( n10003,n10004,n10005 );
   nand U10236 ( n10005,n9453,n9969 );
   nand U10237 ( n10004,instqueue_reg_9__3_,n9970 );
   nor U10238 ( n10002,n9454,n9971 );
   nor U10239 ( n10000,n10006,n10007 );
   nor U10240 ( n10007,n7823,n9974 );
   nor U10241 ( n10006,n8780,n9975 );
   nor U10242 ( n10009,n10010,n10011 );
   nand U10243 ( n10011,n10012,n10013 );
   nand U10244 ( n10013,n9465,n9969 );
   nand U10245 ( n10012,instqueue_reg_9__2_,n9970 );
   nor U10246 ( n10010,n9466,n9971 );
   nor U10247 ( n10008,n10014,n10015 );
   nor U10248 ( n10015,n7825,n9974 );
   nor U10249 ( n10014,n8786,n9975 );
   nor U10250 ( n10017,n10018,n10019 );
   nand U10251 ( n10019,n10020,n10021 );
   nand U10252 ( n10021,n9477,n9969 );
   nand U10253 ( n10020,instqueue_reg_9__1_,n9970 );
   nor U10254 ( n10018,n9478,n9971 );
   nor U10255 ( n10016,n10022,n10023 );
   nor U10256 ( n10023,n7827,n9974 );
   nor U10257 ( n10022,n8793,n9975 );
   nor U10258 ( n10025,n10026,n10027 );
   nand U10259 ( n10027,n10028,n10029 );
   nand U10260 ( n10029,n9489,n9969 );
   nand U10261 ( n9969,n10030,n10031 );
   nand U10262 ( n10031,state2_reg_2_,n10032 );
   nand U10263 ( n10030,n10033,n9493 );
   nand U10264 ( n10028,instqueue_reg_9__0_,n9970 );
   nand U10265 ( n9970,n10034,n10035 );
   nand U10266 ( n10035,state2_reg_3_,n9975 );
   nor U10267 ( n10034,n10036,n10037 );
   nor U10268 ( n10037,n10038,n10039 );
   nand U10269 ( n10039,n10040,n9502 );
   nand U10270 ( n10040,n9503,n10041 );
   nand U10271 ( n10041,n9974,n9971 );
   and U10272 ( n10038,n10033,n9505 );
   nand U10273 ( n10033,n9975,n10042 );
   nand U10274 ( n10042,n9869,n9692 );
   nor U10275 ( n10036,n8790,n10032 );
   nand U10276 ( n10032,n9975,n10043 );
   nand U10277 ( n10043,n9871,n9694 );
   nor U10278 ( n10026,n9512,n9971 );
   nand U10279 ( n9971,n9872,n9695 );
   nor U10280 ( n10024,n10044,n10045 );
   nor U10281 ( n10045,n8767,n9974 );
   nand U10282 ( n9974,n9875,n8924 );
   nor U10283 ( n10044,n8814,n9975 );
   nand U10284 ( n9975,n9876,n9698 );
   nor U10285 ( n10047,n10048,n10049 );
   nand U10286 ( n10049,n10050,n10051 );
   nand U10287 ( n10051,n9400,n10052 );
   nand U10288 ( n10050,instqueue_reg_8__7_,n10053 );
   nor U10289 ( n10048,n8769,n10054 );
   nor U10290 ( n10046,n10055,n10056 );
   nor U10291 ( n10056,n7828,n10057 );
   nor U10292 ( n10055,n8768,n10058 );
   nor U10293 ( n10060,n10061,n10062 );
   nand U10294 ( n10062,n10063,n10064 );
   nand U10295 ( n10064,n9417,n10052 );
   nand U10296 ( n10063,instqueue_reg_8__6_,n10053 );
   nor U10297 ( n10061,n8771,n10054 );
   nor U10298 ( n10059,n10065,n10066 );
   nor U10299 ( n10066,n7826,n10057 );
   nor U10300 ( n10065,n8770,n10058 );
   nor U10301 ( n10068,n10069,n10070 );
   nand U10302 ( n10070,n10071,n10072 );
   nand U10303 ( n10072,n9429,n10052 );
   nand U10304 ( n10071,instqueue_reg_8__5_,n10053 );
   nor U10305 ( n10069,n8773,n10054 );
   nor U10306 ( n10067,n10073,n10074 );
   nor U10307 ( n10074,n7824,n10057 );
   nor U10308 ( n10073,n8772,n10058 );
   nor U10309 ( n10076,n10077,n10078 );
   nand U10310 ( n10078,n10079,n10080 );
   nand U10311 ( n10080,n9441,n10052 );
   nand U10312 ( n10079,instqueue_reg_8__4_,n10053 );
   nor U10313 ( n10077,n8777,n10054 );
   nor U10314 ( n10075,n10081,n10082 );
   nor U10315 ( n10082,n7822,n10057 );
   nor U10316 ( n10081,n8776,n10058 );
   nor U10317 ( n10084,n10085,n10086 );
   nand U10318 ( n10086,n10087,n10088 );
   nand U10319 ( n10088,n9453,n10052 );
   nand U10320 ( n10087,instqueue_reg_8__3_,n10053 );
   nor U10321 ( n10085,n8781,n10054 );
   nor U10322 ( n10083,n10089,n10090 );
   nor U10323 ( n10090,n7823,n10057 );
   nor U10324 ( n10089,n8780,n10058 );
   nor U10325 ( n10092,n10093,n10094 );
   nand U10326 ( n10094,n10095,n10096 );
   nand U10327 ( n10096,n9465,n10052 );
   nand U10328 ( n10095,instqueue_reg_8__2_,n10053 );
   nor U10329 ( n10093,n8787,n10054 );
   nor U10330 ( n10091,n10097,n10098 );
   nor U10331 ( n10098,n7825,n10057 );
   nor U10332 ( n10097,n8786,n10058 );
   nor U10333 ( n10100,n10101,n10102 );
   nand U10334 ( n10102,n10103,n10104 );
   nand U10335 ( n10104,n9477,n10052 );
   nand U10336 ( n10103,instqueue_reg_8__1_,n10053 );
   nor U10337 ( n10101,n8794,n10054 );
   nor U10338 ( n10099,n10105,n10106 );
   nor U10339 ( n10106,n7827,n10057 );
   nor U10340 ( n10105,n8793,n10058 );
   nor U10341 ( n10108,n10109,n10110 );
   nand U10342 ( n10110,n10111,n10112 );
   nand U10343 ( n10112,n9489,n10052 );
   nand U10344 ( n10052,n10113,n10114 );
   nand U10345 ( n10114,n9946,n9694 );
   not U10346 ( n9694,n9779 );
   nand U10347 ( n10113,n10115,n9493 );
   nand U10348 ( n10111,instqueue_reg_8__0_,n10053 );
   nand U10349 ( n10053,n10116,n10117 );
   nand U10350 ( n10117,state2_reg_3_,n10058 );
   nor U10351 ( n10116,n10118,n10119 );
   nor U10352 ( n10119,n10120,n10121 );
   and U10353 ( n10121,n10115,n9505 );
   nand U10354 ( n10115,n10058,n10122 );
   nand U10355 ( n10122,n9869,n8920 );
   nor U10356 ( n9869,n10123,n8947 );
   nor U10357 ( n10120,n10124,n9777 );
   and U10358 ( n10124,n10054,n10057 );
   nor U10359 ( n10118,n10125,n8789 );
   nor U10360 ( n10125,n9779,n9958 );
   nand U10361 ( n9779,n10126,n9959 );
   nor U10362 ( n10109,n8815,n10054 );
   nand U10363 ( n10054,n9872,n9780 );
   nor U10364 ( n10107,n10127,n10128 );
   nor U10365 ( n10128,n8767,n10057 );
   nand U10366 ( n10057,n9875,n9785 );
   nor U10367 ( n9875,n8937,n8954 );
   nor U10368 ( n10127,n8814,n10058 );
   nand U10369 ( n10058,n9876,n9787 );
   nor U10370 ( n10130,n10131,n10132 );
   nand U10371 ( n10132,n10133,n10134 );
   nand U10372 ( n10134,n9400,n10135 );
   nand U10373 ( n10133,instqueue_reg_7__7_,n10136 );
   nor U10374 ( n10131,n9408,n8952 );
   nor U10375 ( n10129,n10137,n10138 );
   nor U10376 ( n10138,n9404,n10139 );
   nor U10377 ( n10137,n9410,n10140 );
   nor U10378 ( n10142,n10143,n10144 );
   nand U10379 ( n10144,n10145,n10146 );
   nand U10380 ( n10146,n9417,n10135 );
   nand U10381 ( n10145,instqueue_reg_7__6_,n10136 );
   nor U10382 ( n10143,n9421,n8952 );
   nor U10383 ( n10141,n10147,n10148 );
   nor U10384 ( n10148,n9418,n10139 );
   nor U10385 ( n10147,n9422,n10140 );
   nor U10386 ( n10150,n10151,n10152 );
   nand U10387 ( n10152,n10153,n10154 );
   nand U10388 ( n10154,n9429,n10135 );
   nand U10389 ( n10153,instqueue_reg_7__5_,n10136 );
   nor U10390 ( n10151,n9433,n8952 );
   nor U10391 ( n10149,n10155,n10156 );
   nor U10392 ( n10156,n9430,n10139 );
   nor U10393 ( n10155,n9434,n10140 );
   nor U10394 ( n10158,n10159,n10160 );
   nand U10395 ( n10160,n10161,n10162 );
   nand U10396 ( n10162,n9441,n10135 );
   nand U10397 ( n10161,instqueue_reg_7__4_,n10136 );
   nor U10398 ( n10159,n9445,n8952 );
   nor U10399 ( n10157,n10163,n10164 );
   nor U10400 ( n10164,n9442,n10139 );
   nor U10401 ( n10163,n9446,n10140 );
   nor U10402 ( n10166,n10167,n10168 );
   nand U10403 ( n10168,n10169,n10170 );
   nand U10404 ( n10170,n9453,n10135 );
   nand U10405 ( n10169,instqueue_reg_7__3_,n10136 );
   nor U10406 ( n10167,n9457,n8952 );
   nor U10407 ( n10165,n10171,n10172 );
   nor U10408 ( n10172,n9454,n10139 );
   nor U10409 ( n10171,n9458,n10140 );
   nor U10410 ( n10174,n10175,n10176 );
   nand U10411 ( n10176,n10177,n10178 );
   nand U10412 ( n10178,n9465,n10135 );
   nand U10413 ( n10177,instqueue_reg_7__2_,n10136 );
   nor U10414 ( n10175,n9469,n8952 );
   nor U10415 ( n10173,n10179,n10180 );
   nor U10416 ( n10180,n9466,n10139 );
   nor U10417 ( n10179,n9470,n10140 );
   nor U10418 ( n10182,n10183,n10184 );
   nand U10419 ( n10184,n10185,n10186 );
   nand U10420 ( n10186,n9477,n10135 );
   nand U10421 ( n10185,instqueue_reg_7__1_,n10136 );
   nor U10422 ( n10183,n9481,n8952 );
   nor U10423 ( n10181,n10187,n10188 );
   nor U10424 ( n10188,n9478,n10139 );
   nor U10425 ( n10187,n9482,n10140 );
   nor U10426 ( n10190,n10191,n10192 );
   nand U10427 ( n10192,n10193,n10194 );
   nand U10428 ( n10194,n9489,n10135 );
   nand U10429 ( n10135,n10195,n10196 );
   nand U10430 ( n10196,state2_reg_2_,n10197 );
   nand U10431 ( n10195,n10198,n9493 );
   nand U10432 ( n10193,instqueue_reg_7__0_,n10136 );
   nand U10433 ( n10136,n10199,n10200 );
   nor U10434 ( n10200,n10201,n10202 );
   nor U10435 ( n10202,n8871,n10197 );
   nand U10436 ( n10197,n10140,n10203 );
   nand U10437 ( n10203,n10204,n9510 );
   nor U10438 ( n10201,n10198,n10205 );
   nand U10439 ( n10205,n10206,n10207 );
   not U10440 ( n10207,n10208 );
   nand U10441 ( n10206,n10209,n10210 );
   nand U10442 ( n10210,n10139,n8952 );
   nand U10443 ( n10198,n10140,n10211 );
   nand U10444 ( n10211,n10212,n9508 );
   nor U10445 ( n10199,n10213,n9602 );
   nor U10446 ( n10213,n10214,n9018 );
   nor U10447 ( n10191,n9517,n8952 );
   nand U10448 ( n8952,n8953,n8954 );
   not U10449 ( n8954,n9518 );
   not U10450 ( n8953,n8936 );
   nand U10451 ( n8936,n8938,n8937 );
   nor U10452 ( n10189,n10215,n10216 );
   nor U10453 ( n10216,n9512,n10139 );
   nor U10454 ( n10215,n9519,n10140 );
   nor U10455 ( n10218,n10219,n10220 );
   nand U10456 ( n10220,n10221,n10222 );
   nand U10457 ( n10222,n9400,n10223 );
   nand U10458 ( n10221,instqueue_reg_6__7_,n10224 );
   nor U10459 ( n10219,n9404,n10225 );
   nor U10460 ( n10217,n10226,n10227 );
   nor U10461 ( n10227,n7828,n10228 );
   nor U10462 ( n10226,n8768,n10229 );
   nor U10463 ( n10231,n10232,n10233 );
   nand U10464 ( n10233,n10234,n10235 );
   nand U10465 ( n10235,n9417,n10223 );
   nand U10466 ( n10234,instqueue_reg_6__6_,n10224 );
   nor U10467 ( n10232,n9418,n10225 );
   nor U10468 ( n10230,n10236,n10237 );
   nor U10469 ( n10237,n7826,n10228 );
   nor U10470 ( n10236,n8770,n10229 );
   nor U10471 ( n10239,n10240,n10241 );
   nand U10472 ( n10241,n10242,n10243 );
   nand U10473 ( n10243,n9429,n10223 );
   nand U10474 ( n10242,instqueue_reg_6__5_,n10224 );
   nor U10475 ( n10240,n9430,n10225 );
   nor U10476 ( n10238,n10244,n10245 );
   nor U10477 ( n10245,n7824,n10228 );
   nor U10478 ( n10244,n8772,n10229 );
   nor U10479 ( n10247,n10248,n10249 );
   nand U10480 ( n10249,n10250,n10251 );
   nand U10481 ( n10251,n9441,n10223 );
   nand U10482 ( n10250,instqueue_reg_6__4_,n10224 );
   nor U10483 ( n10248,n9442,n10225 );
   nor U10484 ( n10246,n10252,n10253 );
   nor U10485 ( n10253,n7822,n10228 );
   nor U10486 ( n10252,n8776,n10229 );
   nor U10487 ( n10255,n10256,n10257 );
   nand U10488 ( n10257,n10258,n10259 );
   nand U10489 ( n10259,n9453,n10223 );
   nand U10490 ( n10258,instqueue_reg_6__3_,n10224 );
   nor U10491 ( n10256,n9454,n10225 );
   nor U10492 ( n10254,n10260,n10261 );
   nor U10493 ( n10261,n7823,n10228 );
   nor U10494 ( n10260,n8780,n10229 );
   nor U10495 ( n10263,n10264,n10265 );
   nand U10496 ( n10265,n10266,n10267 );
   nand U10497 ( n10267,n9465,n10223 );
   nand U10498 ( n10266,instqueue_reg_6__2_,n10224 );
   nor U10499 ( n10264,n9466,n10225 );
   nor U10500 ( n10262,n10268,n10269 );
   nor U10501 ( n10269,n7825,n10228 );
   nor U10502 ( n10268,n8786,n10229 );
   nor U10503 ( n10271,n10272,n10273 );
   nand U10504 ( n10273,n10274,n10275 );
   nand U10505 ( n10275,n9477,n10223 );
   nand U10506 ( n10274,instqueue_reg_6__1_,n10224 );
   nor U10507 ( n10272,n9478,n10225 );
   nor U10508 ( n10270,n10276,n10277 );
   nor U10509 ( n10277,n7827,n10228 );
   nor U10510 ( n10276,n8793,n10229 );
   nor U10511 ( n10279,n10280,n10281 );
   nand U10512 ( n10281,n10282,n10283 );
   nand U10513 ( n10283,n9489,n10223 );
   nand U10514 ( n10223,n10284,n10285 );
   nand U10515 ( n10285,n10204,n9591 );
   nand U10516 ( n10284,n10286,n9493 );
   not U10517 ( n10286,n10287 );
   nand U10518 ( n10282,instqueue_reg_6__0_,n10224 );
   nand U10519 ( n10224,n10288,n10289 );
   nand U10520 ( n10289,state2_reg_3_,n10229 );
   nor U10521 ( n10288,n10290,n10291 );
   nor U10522 ( n10291,n10292,n10293 );
   nand U10523 ( n10293,n10294,n9502 );
   nand U10524 ( n10294,n9503,n10295 );
   nand U10525 ( n10295,n10228,n10225 );
   nor U10526 ( n10292,n10287,n9602 );
   nand U10527 ( n10287,n10212,n9603 );
   nor U10528 ( n10290,n10296,n8790 );
   nor U10529 ( n10296,n9605,n10297 );
   nor U10530 ( n10280,n9512,n10225 );
   nand U10531 ( n10225,n9607,n10298 );
   nor U10532 ( n10278,n10299,n10300 );
   nor U10533 ( n10300,n8767,n10228 );
   nand U10534 ( n10228,n10301,n8923 );
   nor U10535 ( n10299,n8814,n10229 );
   nand U10536 ( n10229,n9611,n10302 );
   nor U10537 ( n10304,n10305,n10306 );
   nand U10538 ( n10306,n10307,n10308 );
   nand U10539 ( n10308,n9400,n10309 );
   nand U10540 ( n10307,instqueue_reg_5__7_,n10310 );
   nor U10541 ( n10305,n8769,n10311 );
   nor U10542 ( n10303,n10312,n10313 );
   nor U10543 ( n10313,n9408,n10314 );
   nor U10544 ( n10312,n9410,n10315 );
   nor U10545 ( n10317,n10318,n10319 );
   nand U10546 ( n10319,n10320,n10321 );
   nand U10547 ( n10321,n9417,n10309 );
   nand U10548 ( n10320,instqueue_reg_5__6_,n10310 );
   nor U10549 ( n10318,n8771,n10311 );
   nor U10550 ( n10316,n10322,n10323 );
   nor U10551 ( n10323,n9421,n10314 );
   nor U10552 ( n10322,n9422,n10315 );
   nor U10553 ( n10325,n10326,n10327 );
   nand U10554 ( n10327,n10328,n10329 );
   nand U10555 ( n10329,n9429,n10309 );
   nand U10556 ( n10328,instqueue_reg_5__5_,n10310 );
   nor U10557 ( n10326,n8773,n10311 );
   nor U10558 ( n10324,n10330,n10331 );
   nor U10559 ( n10331,n9433,n10314 );
   nor U10560 ( n10330,n9434,n10315 );
   nor U10561 ( n10333,n10334,n10335 );
   nand U10562 ( n10335,n10336,n10337 );
   nand U10563 ( n10337,n9441,n10309 );
   nand U10564 ( n10336,instqueue_reg_5__4_,n10310 );
   nor U10565 ( n10334,n8777,n10311 );
   nor U10566 ( n10332,n10338,n10339 );
   nor U10567 ( n10339,n9445,n10314 );
   nor U10568 ( n10338,n9446,n10315 );
   nor U10569 ( n10341,n10342,n10343 );
   nand U10570 ( n10343,n10344,n10345 );
   nand U10571 ( n10345,n9453,n10309 );
   nand U10572 ( n10344,instqueue_reg_5__3_,n10310 );
   nor U10573 ( n10342,n8781,n10311 );
   nor U10574 ( n10340,n10346,n10347 );
   nor U10575 ( n10347,n9457,n10314 );
   nor U10576 ( n10346,n9458,n10315 );
   nor U10577 ( n10349,n10350,n10351 );
   nand U10578 ( n10351,n10352,n10353 );
   nand U10579 ( n10353,n9465,n10309 );
   nand U10580 ( n10352,instqueue_reg_5__2_,n10310 );
   nor U10581 ( n10350,n8787,n10311 );
   nor U10582 ( n10348,n10354,n10355 );
   nor U10583 ( n10355,n9469,n10314 );
   nor U10584 ( n10354,n9470,n10315 );
   nor U10585 ( n10357,n10358,n10359 );
   nand U10586 ( n10359,n10360,n10361 );
   nand U10587 ( n10361,n9477,n10309 );
   nand U10588 ( n10360,instqueue_reg_5__1_,n10310 );
   nor U10589 ( n10358,n8794,n10311 );
   nor U10590 ( n10356,n10362,n10363 );
   nor U10591 ( n10363,n9481,n10314 );
   nor U10592 ( n10362,n9482,n10315 );
   nor U10593 ( n10365,n10366,n10367 );
   nand U10594 ( n10367,n10368,n10369 );
   nand U10595 ( n10369,n9489,n10309 );
   nand U10596 ( n10309,n10370,n10371 );
   nand U10597 ( n10371,state2_reg_2_,n10372 );
   nand U10598 ( n10370,n10373,n9493 );
   nand U10599 ( n10368,instqueue_reg_5__0_,n10310 );
   nand U10600 ( n10310,n10374,n10375 );
   nand U10601 ( n10375,state2_reg_3_,n10315 );
   nor U10602 ( n10374,n10376,n10377 );
   nor U10603 ( n10377,n10378,n10379 );
   nand U10604 ( n10379,n10380,n9502 );
   nand U10605 ( n10380,n9503,n10381 );
   nand U10606 ( n10381,n10314,n10311 );
   and U10607 ( n10378,n10373,n9505 );
   nand U10608 ( n10373,n10315,n10382 );
   nand U10609 ( n10382,n10212,n9692 );
   nor U10610 ( n10376,n8871,n10372 );
   nand U10611 ( n10372,n10315,n10383 );
   nand U10612 ( n10383,n10384,n9510 );
   nor U10613 ( n9510,n9605,instqueuewr_addr_reg_0_ );
   nor U10614 ( n10366,n8815,n10311 );
   nand U10615 ( n10311,n9695,n10298 );
   nor U10616 ( n10364,n10385,n10386 );
   nor U10617 ( n10386,n9517,n10314 );
   nand U10618 ( n10314,n10301,n8924 );
   nor U10619 ( n10385,n9519,n10315 );
   nand U10620 ( n10315,n9698,n10302 );
   nor U10621 ( n10388,n10389,n10390 );
   nand U10622 ( n10390,n10391,n10392 );
   nand U10623 ( n10392,n9400,n10393 );
   nand U10624 ( n10391,instqueue_reg_4__7_,n10394 );
   nor U10625 ( n10389,n8769,n10395 );
   nor U10626 ( n10387,n10396,n10397 );
   nor U10627 ( n10397,n9408,n10398 );
   nor U10628 ( n10396,n9410,n10399 );
   nor U10629 ( n10401,n10402,n10403 );
   nand U10630 ( n10403,n10404,n10405 );
   nand U10631 ( n10405,n9417,n10393 );
   nand U10632 ( n10404,instqueue_reg_4__6_,n10394 );
   nor U10633 ( n10402,n8771,n10395 );
   nor U10634 ( n10400,n10406,n10407 );
   nor U10635 ( n10407,n9421,n10398 );
   nor U10636 ( n10406,n9422,n10399 );
   nor U10637 ( n10409,n10410,n10411 );
   nand U10638 ( n10411,n10412,n10413 );
   nand U10639 ( n10413,n9429,n10393 );
   nand U10640 ( n10412,instqueue_reg_4__5_,n10394 );
   nor U10641 ( n10410,n8773,n10395 );
   nor U10642 ( n10408,n10414,n10415 );
   nor U10643 ( n10415,n9433,n10398 );
   nor U10644 ( n10414,n9434,n10399 );
   nor U10645 ( n10417,n10418,n10419 );
   nand U10646 ( n10419,n10420,n10421 );
   nand U10647 ( n10421,n9441,n10393 );
   nand U10648 ( n10420,instqueue_reg_4__4_,n10394 );
   nor U10649 ( n10418,n8777,n10395 );
   nor U10650 ( n10416,n10422,n10423 );
   nor U10651 ( n10423,n9445,n10398 );
   nor U10652 ( n10422,n9446,n10399 );
   nor U10653 ( n10425,n10426,n10427 );
   nand U10654 ( n10427,n10428,n10429 );
   nand U10655 ( n10429,n9453,n10393 );
   nand U10656 ( n10428,instqueue_reg_4__3_,n10394 );
   nor U10657 ( n10426,n8781,n10395 );
   nor U10658 ( n10424,n10430,n10431 );
   nor U10659 ( n10431,n9457,n10398 );
   nor U10660 ( n10430,n9458,n10399 );
   nor U10661 ( n10433,n10434,n10435 );
   nand U10662 ( n10435,n10436,n10437 );
   nand U10663 ( n10437,n9465,n10393 );
   nand U10664 ( n10436,instqueue_reg_4__2_,n10394 );
   nor U10665 ( n10434,n8787,n10395 );
   nor U10666 ( n10432,n10438,n10439 );
   nor U10667 ( n10439,n9469,n10398 );
   nor U10668 ( n10438,n9470,n10399 );
   nor U10669 ( n10441,n10442,n10443 );
   nand U10670 ( n10443,n10444,n10445 );
   nand U10671 ( n10445,n9477,n10393 );
   nand U10672 ( n10444,instqueue_reg_4__1_,n10394 );
   nor U10673 ( n10442,n8794,n10395 );
   nor U10674 ( n10440,n10446,n10447 );
   nor U10675 ( n10447,n9481,n10398 );
   nor U10676 ( n10446,n9482,n10399 );
   nor U10677 ( n10449,n10450,n10451 );
   nand U10678 ( n10451,n10452,n10453 );
   nand U10679 ( n10453,n9489,n10393 );
   nand U10680 ( n10393,n10454,n10455 );
   nand U10681 ( n10455,n10384,n9591 );
   nor U10682 ( n9591,n8790,n9605 );
   nand U10683 ( n10454,n10456,n9493 );
   not U10684 ( n10456,n10457 );
   nand U10685 ( n10452,instqueue_reg_4__0_,n10394 );
   nand U10686 ( n10394,n10458,n10459 );
   nand U10687 ( n10459,state2_reg_3_,n10399 );
   nor U10688 ( n10458,n10460,n10461 );
   nor U10689 ( n10461,n10462,n10463 );
   nand U10690 ( n10463,n10464,n9502 );
   nand U10691 ( n10464,n9503,n10465 );
   nand U10692 ( n10465,n10398,n10395 );
   nor U10693 ( n10462,n10457,n9602 );
   nand U10694 ( n10457,n10212,n8920 );
   nor U10695 ( n10212,n8933,n10466 );
   nor U10696 ( n10460,n10467,n8789 );
   nor U10697 ( n10467,n9605,n10468 );
   nor U10698 ( n10450,n8815,n10395 );
   nand U10699 ( n10395,n9780,n10298 );
   nor U10700 ( n10448,n10469,n10470 );
   nor U10701 ( n10470,n9517,n10398 );
   nand U10702 ( n10398,n10301,n9785 );
   nor U10703 ( n10301,n9518,n9786 );
   not U10704 ( n9786,n8937 );
   nor U10705 ( n10469,n9519,n10399 );
   nand U10706 ( n10399,n9787,n10302 );
   nor U10707 ( n10472,n10473,n10474 );
   nand U10708 ( n10474,n10475,n10476 );
   nand U10709 ( n10476,n9400,n10477 );
   nand U10710 ( n10475,instqueue_reg_3__7_,n10478 );
   nor U10711 ( n10473,n8769,n10479 );
   nor U10712 ( n10471,n10480,n10481 );
   nor U10713 ( n10481,n9408,n10482 );
   nor U10714 ( n10480,n9410,n10483 );
   nor U10715 ( n10485,n10486,n10487 );
   nand U10716 ( n10487,n10488,n10489 );
   nand U10717 ( n10489,n9417,n10477 );
   nand U10718 ( n10488,instqueue_reg_3__6_,n10478 );
   nor U10719 ( n10486,n8771,n10479 );
   nor U10720 ( n10484,n10490,n10491 );
   nor U10721 ( n10491,n9421,n10482 );
   nor U10722 ( n10490,n9422,n10483 );
   nor U10723 ( n10493,n10494,n10495 );
   nand U10724 ( n10495,n10496,n10497 );
   nand U10725 ( n10497,n9429,n10477 );
   nand U10726 ( n10496,instqueue_reg_3__5_,n10478 );
   nor U10727 ( n10494,n8773,n10479 );
   nor U10728 ( n10492,n10498,n10499 );
   nor U10729 ( n10499,n9433,n10482 );
   nor U10730 ( n10498,n9434,n10483 );
   nor U10731 ( n10501,n10502,n10503 );
   nand U10732 ( n10503,n10504,n10505 );
   nand U10733 ( n10505,n9441,n10477 );
   nand U10734 ( n10504,instqueue_reg_3__4_,n10478 );
   nor U10735 ( n10502,n8777,n10479 );
   nor U10736 ( n10500,n10506,n10507 );
   nor U10737 ( n10507,n9445,n10482 );
   nor U10738 ( n10506,n9446,n10483 );
   nor U10739 ( n10509,n10510,n10511 );
   nand U10740 ( n10511,n10512,n10513 );
   nand U10741 ( n10513,n9453,n10477 );
   nand U10742 ( n10512,instqueue_reg_3__3_,n10478 );
   nor U10743 ( n10510,n8781,n10479 );
   nor U10744 ( n10508,n10514,n10515 );
   nor U10745 ( n10515,n9457,n10482 );
   nor U10746 ( n10514,n9458,n10483 );
   nor U10747 ( n10517,n10518,n10519 );
   nand U10748 ( n10519,n10520,n10521 );
   nand U10749 ( n10521,n9465,n10477 );
   nand U10750 ( n10520,instqueue_reg_3__2_,n10478 );
   nor U10751 ( n10518,n8787,n10479 );
   nor U10752 ( n10516,n10522,n10523 );
   nor U10753 ( n10523,n9469,n10482 );
   nor U10754 ( n10522,n9470,n10483 );
   nor U10755 ( n10525,n10526,n10527 );
   nand U10756 ( n10527,n10528,n10529 );
   nand U10757 ( n10529,n9477,n10477 );
   nand U10758 ( n10528,instqueue_reg_3__1_,n10478 );
   nor U10759 ( n10526,n8794,n10479 );
   nor U10760 ( n10524,n10530,n10531 );
   nor U10761 ( n10531,n9481,n10482 );
   nor U10762 ( n10530,n9482,n10483 );
   nor U10763 ( n10533,n10534,n10535 );
   nand U10764 ( n10535,n10536,n10537 );
   nand U10765 ( n10537,n9489,n10477 );
   nand U10766 ( n10477,n10538,n10539 );
   nand U10767 ( n10539,state2_reg_2_,n10540 );
   nand U10768 ( n10538,n10541,n9493 );
   nand U10769 ( n10536,instqueue_reg_3__0_,n10478 );
   nand U10770 ( n10478,n10542,n10543 );
   nand U10771 ( n10543,state2_reg_3_,n10483 );
   nor U10772 ( n10542,n10544,n10545 );
   nor U10773 ( n10545,n10546,n10547 );
   nand U10774 ( n10547,n10548,n9502 );
   nand U10775 ( n10548,n9503,n10549 );
   nand U10776 ( n10549,n10482,n10479 );
   and U10777 ( n10546,n10541,n9505 );
   nand U10778 ( n10541,n10483,n10550 );
   nand U10779 ( n10550,n10551,n9508 );
   nor U10780 ( n9508,n8910,n8920 );
   nor U10781 ( n10544,n8789,n10540 );
   nand U10782 ( n10540,n10483,n10552 );
   nand U10783 ( n10552,n10204,n9871 );
   nor U10784 ( n10534,n8815,n10479 );
   nand U10785 ( n10479,n10553,n9514 );
   nor U10786 ( n10532,n10554,n10555 );
   nor U10787 ( n10555,n9517,n10482 );
   nand U10788 ( n10482,n10556,n8938 );
   nor U10789 ( n8938,n8905,n10557 );
   nor U10790 ( n10554,n9519,n10483 );
   nand U10791 ( n10483,n10558,n9521 );
   nor U10792 ( n10560,n10561,n10562 );
   nand U10793 ( n10562,n10563,n10564 );
   nand U10794 ( n10564,n9400,n10565 );
   nand U10795 ( n10563,instqueue_reg_2__7_,n10566 );
   nor U10796 ( n10561,n8769,n10567 );
   nor U10797 ( n10559,n10568,n10569 );
   nor U10798 ( n10569,n9408,n10570 );
   nor U10799 ( n10568,n9410,n10571 );
   nor U10800 ( n10573,n10574,n10575 );
   nand U10801 ( n10575,n10576,n10577 );
   nand U10802 ( n10577,n9417,n10565 );
   nand U10803 ( n10576,instqueue_reg_2__6_,n10566 );
   nor U10804 ( n10574,n8771,n10567 );
   nor U10805 ( n10572,n10578,n10579 );
   nor U10806 ( n10579,n9421,n10570 );
   nor U10807 ( n10578,n9422,n10571 );
   nor U10808 ( n10581,n10582,n10583 );
   nand U10809 ( n10583,n10584,n10585 );
   nand U10810 ( n10585,n9429,n10565 );
   nand U10811 ( n10584,instqueue_reg_2__5_,n10566 );
   nor U10812 ( n10582,n8773,n10567 );
   nor U10813 ( n10580,n10586,n10587 );
   nor U10814 ( n10587,n9433,n10570 );
   nor U10815 ( n10586,n9434,n10571 );
   nor U10816 ( n10589,n10590,n10591 );
   nand U10817 ( n10591,n10592,n10593 );
   nand U10818 ( n10593,n9441,n10565 );
   nand U10819 ( n10592,instqueue_reg_2__4_,n10566 );
   nor U10820 ( n10590,n8777,n10567 );
   nor U10821 ( n10588,n10594,n10595 );
   nor U10822 ( n10595,n9445,n10570 );
   nor U10823 ( n10594,n9446,n10571 );
   nor U10824 ( n10597,n10598,n10599 );
   nand U10825 ( n10599,n10600,n10601 );
   nand U10826 ( n10601,n9453,n10565 );
   nand U10827 ( n10600,instqueue_reg_2__3_,n10566 );
   nor U10828 ( n10598,n8781,n10567 );
   nor U10829 ( n10596,n10602,n10603 );
   nor U10830 ( n10603,n9457,n10570 );
   nor U10831 ( n10602,n9458,n10571 );
   nor U10832 ( n10605,n10606,n10607 );
   nand U10833 ( n10607,n10608,n10609 );
   nand U10834 ( n10609,n9465,n10565 );
   nand U10835 ( n10608,instqueue_reg_2__2_,n10566 );
   nor U10836 ( n10606,n8787,n10567 );
   nor U10837 ( n10604,n10610,n10611 );
   nor U10838 ( n10611,n9469,n10570 );
   nor U10839 ( n10610,n9470,n10571 );
   nor U10840 ( n10613,n10614,n10615 );
   nand U10841 ( n10615,n10616,n10617 );
   nand U10842 ( n10617,n9477,n10565 );
   nand U10843 ( n10616,instqueue_reg_2__1_,n10566 );
   nor U10844 ( n10614,n8794,n10567 );
   nor U10845 ( n10612,n10618,n10619 );
   nor U10846 ( n10619,n9481,n10570 );
   nor U10847 ( n10618,n9482,n10571 );
   nor U10848 ( n10621,n10622,n10623 );
   nand U10849 ( n10623,n10624,n10625 );
   nand U10850 ( n10625,n9489,n10565 );
   nand U10851 ( n10565,n10626,n10627 );
   nand U10852 ( n10627,n10204,n9946 );
   not U10853 ( n10204,n10297 );
   nand U10854 ( n10626,n10628,n9493 );
   not U10855 ( n10628,n10629 );
   nand U10856 ( n10624,instqueue_reg_2__0_,n10566 );
   nand U10857 ( n10566,n10630,n10631 );
   nand U10858 ( n10631,state2_reg_3_,n10571 );
   nor U10859 ( n10630,n10632,n10633 );
   nor U10860 ( n10633,n10634,n10635 );
   nand U10861 ( n10635,n10636,n9502 );
   nand U10862 ( n10636,n9503,n10637 );
   nand U10863 ( n10637,n10570,n10567 );
   nor U10864 ( n10634,n10629,n9602 );
   nand U10865 ( n10629,n10551,n9603 );
   nor U10866 ( n10632,n10638,n8790 );
   nor U10867 ( n10638,n9958,n10297 );
   nand U10868 ( n10297,n10639,n9960 );
   not U10869 ( n9960,n10126 );
   nor U10870 ( n10622,n8815,n10567 );
   nand U10871 ( n10567,n10553,n9607 );
   nor U10872 ( n10620,n10640,n10641 );
   nor U10873 ( n10641,n9517,n10570 );
   nand U10874 ( n10570,n10556,n8923 );
   nor U10875 ( n8923,n10642,n10557 );
   nor U10876 ( n10640,n9519,n10571 );
   nand U10877 ( n10571,n10558,n9611 );
   nor U10878 ( n10644,n10645,n10646 );
   nand U10879 ( n10646,n10647,n10648 );
   nand U10880 ( n10648,n9400,n10649 );
   not U10881 ( n9400,n10650 );
   nand U10882 ( n10647,instqueue_reg_1__7_,n10651 );
   nor U10883 ( n10645,n8769,n10652 );
   nor U10884 ( n10643,n10653,n10654 );
   nor U10885 ( n10654,n9408,n10655 );
   nor U10886 ( n10653,n9410,n10656 );
   nor U10887 ( n10658,n10659,n10660 );
   nand U10888 ( n10660,n10661,n10662 );
   nand U10889 ( n10662,n9417,n10649 );
   not U10890 ( n9417,n10663 );
   nand U10891 ( n10661,instqueue_reg_1__6_,n10651 );
   nor U10892 ( n10659,n8771,n10652 );
   nor U10893 ( n10657,n10664,n10665 );
   nor U10894 ( n10665,n9421,n10655 );
   nor U10895 ( n10664,n9422,n10656 );
   nor U10896 ( n10667,n10668,n10669 );
   nand U10897 ( n10669,n10670,n10671 );
   nand U10898 ( n10671,n9429,n10649 );
   not U10899 ( n9429,n10672 );
   nand U10900 ( n10670,instqueue_reg_1__5_,n10651 );
   nor U10901 ( n10668,n8773,n10652 );
   nor U10902 ( n10666,n10673,n10674 );
   nor U10903 ( n10674,n9433,n10655 );
   nor U10904 ( n10673,n9434,n10656 );
   nor U10905 ( n10676,n10677,n10678 );
   nand U10906 ( n10678,n10679,n10680 );
   nand U10907 ( n10680,n9441,n10649 );
   not U10908 ( n9441,n10681 );
   nand U10909 ( n10679,instqueue_reg_1__4_,n10651 );
   nor U10910 ( n10677,n8777,n10652 );
   nor U10911 ( n10675,n10682,n10683 );
   nor U10912 ( n10683,n9445,n10655 );
   nor U10913 ( n10682,n9446,n10656 );
   nor U10914 ( n10685,n10686,n10687 );
   nand U10915 ( n10687,n10688,n10689 );
   nand U10916 ( n10689,n9453,n10649 );
   not U10917 ( n9453,n10690 );
   nand U10918 ( n10688,instqueue_reg_1__3_,n10651 );
   nor U10919 ( n10686,n8781,n10652 );
   nor U10920 ( n10684,n10691,n10692 );
   nor U10921 ( n10692,n9457,n10655 );
   nor U10922 ( n10691,n9458,n10656 );
   nor U10923 ( n10694,n10695,n10696 );
   nand U10924 ( n10696,n10697,n10698 );
   nand U10925 ( n10698,n9465,n10649 );
   not U10926 ( n9465,n10699 );
   nand U10927 ( n10697,instqueue_reg_1__2_,n10651 );
   nor U10928 ( n10695,n8787,n10652 );
   nor U10929 ( n10693,n10700,n10701 );
   nor U10930 ( n10701,n9469,n10655 );
   nor U10931 ( n10700,n9470,n10656 );
   nor U10932 ( n10703,n10704,n10705 );
   nand U10933 ( n10705,n10706,n10707 );
   nand U10934 ( n10707,n9477,n10649 );
   not U10935 ( n9477,n10708 );
   nand U10936 ( n10706,instqueue_reg_1__1_,n10651 );
   nor U10937 ( n10704,n8794,n10652 );
   nor U10938 ( n10702,n10709,n10710 );
   nor U10939 ( n10710,n9481,n10655 );
   nor U10940 ( n10709,n9482,n10656 );
   nor U10941 ( n10712,n10713,n10714 );
   nand U10942 ( n10714,n10715,n10716 );
   nand U10943 ( n10716,n9489,n10649 );
   nand U10944 ( n10649,n10717,n10718 );
   nand U10945 ( n10718,state2_reg_2_,n10719 );
   nand U10946 ( n10717,n10720,n9493 );
   not U10947 ( n9489,n10721 );
   nand U10948 ( n10715,instqueue_reg_1__0_,n10651 );
   nand U10949 ( n10651,n10722,n10723 );
   nand U10950 ( n10723,state2_reg_3_,n10656 );
   nor U10951 ( n10722,n10724,n10725 );
   nor U10952 ( n10725,n10726,n10727 );
   nand U10953 ( n10727,n10728,n9502 );
   nand U10954 ( n10728,n9503,n10729 );
   nand U10955 ( n10729,n10655,n10652 );
   and U10956 ( n10726,n10720,n9505 );
   nand U10957 ( n10720,n10656,n10730 );
   nand U10958 ( n10730,n10551,n9692 );
   nor U10959 ( n9692,n8910,n9603 );
   nor U10960 ( n10724,n8789,n10719 );
   nand U10961 ( n10719,n10656,n10731 );
   nand U10962 ( n10731,n10384,n9871 );
   nor U10963 ( n9871,n9958,instqueuewr_addr_reg_0_ );
   nor U10964 ( n10713,n8815,n10652 );
   nand U10965 ( n10652,n10553,n9695 );
   nor U10966 ( n10711,n10732,n10733 );
   nor U10967 ( n10733,n9517,n10655 );
   nand U10968 ( n10655,n10556,n8924 );
   nor U10969 ( n8924,n10734,n8905 );
   nor U10970 ( n10732,n9519,n10656 );
   nand U10971 ( n10656,n10558,n9698 );
   nor U10972 ( n10736,n10737,n10738 );
   nand U10973 ( n10738,n10739,n10740 );
   or U10974 ( n10740,n10741,n7828 );
   nand U10975 ( n9408,datai_31_,n10742 );
   or U10976 ( n10739,n10743,n8768 );
   nand U10977 ( n9410,n10744,n10745 );
   nor U10978 ( n10737,n9404,n10746 );
   nand U10979 ( n9404,datai_23_,n10742 );
   nor U10980 ( n10735,n10747,n10748 );
   nor U10981 ( n10748,n10749,n10750 );
   nor U10982 ( n10747,n10751,n10650 );
   nand U10983 ( n10650,datai_7_,n9505 );
   nor U10984 ( n10753,n10754,n10755 );
   nand U10985 ( n10755,n10756,n10757 );
   or U10986 ( n10757,n10741,n7826 );
   nand U10987 ( n9421,datai_30_,n10742 );
   or U10988 ( n10756,n10743,n8770 );
   nand U10989 ( n9422,n10744,n10758 );
   nor U10990 ( n10754,n9418,n10746 );
   nand U10991 ( n9418,datai_22_,n10742 );
   nor U10992 ( n10752,n10759,n10760 );
   nor U10993 ( n10760,n10749,n10761 );
   nor U10994 ( n10759,n10751,n10663 );
   nand U10995 ( n10663,datai_6_,n9505 );
   nor U10996 ( n10763,n10764,n10765 );
   nand U10997 ( n10765,n10766,n10767 );
   or U10998 ( n10767,n10741,n7824 );
   nand U10999 ( n9433,datai_29_,n10742 );
   or U11000 ( n10766,n10743,n8772 );
   nand U11001 ( n9434,n10744,n10768 );
   nor U11002 ( n10764,n9430,n10746 );
   nand U11003 ( n9430,datai_21_,n10742 );
   nor U11004 ( n10762,n10769,n10770 );
   nor U11005 ( n10770,n10749,n10771 );
   nor U11006 ( n10769,n10751,n10672 );
   nand U11007 ( n10672,datai_5_,n9505 );
   nor U11008 ( n10773,n10774,n10775 );
   nand U11009 ( n10775,n10776,n10777 );
   or U11010 ( n10777,n10741,n7822 );
   nand U11011 ( n9445,datai_28_,n10742 );
   or U11012 ( n10776,n10743,n8776 );
   nand U11013 ( n9446,n10744,n10778 );
   nor U11014 ( n10774,n9442,n10746 );
   nand U11015 ( n9442,datai_20_,n10742 );
   nor U11016 ( n10772,n10779,n10780 );
   nor U11017 ( n10780,n10749,n10781 );
   nor U11018 ( n10779,n10751,n10681 );
   nand U11019 ( n10681,datai_4_,n9505 );
   nor U11020 ( n10783,n10784,n10785 );
   nand U11021 ( n10785,n10786,n10787 );
   or U11022 ( n10787,n10741,n7823 );
   nand U11023 ( n9457,datai_27_,n10742 );
   or U11024 ( n10786,n10743,n8780 );
   nand U11025 ( n9458,n10744,n10788 );
   nor U11026 ( n10784,n9454,n10746 );
   nand U11027 ( n9454,datai_19_,n10742 );
   nor U11028 ( n10782,n10789,n10790 );
   nor U11029 ( n10790,n10749,n10791 );
   nor U11030 ( n10789,n10751,n10690 );
   nand U11031 ( n10690,datai_3_,n9505 );
   nor U11032 ( n10793,n10794,n10795 );
   nand U11033 ( n10795,n10796,n10797 );
   or U11034 ( n10797,n10741,n7825 );
   nand U11035 ( n9469,datai_26_,n10742 );
   or U11036 ( n10796,n10743,n8786 );
   nand U11037 ( n9470,n10744,n10798 );
   nor U11038 ( n10794,n9466,n10746 );
   nand U11039 ( n9466,datai_18_,n10742 );
   nor U11040 ( n10792,n10799,n10800 );
   nor U11041 ( n10800,n10749,n10801 );
   nor U11042 ( n10799,n10751,n10699 );
   nand U11043 ( n10699,datai_2_,n9505 );
   nor U11044 ( n10803,n10804,n10805 );
   nand U11045 ( n10805,n10806,n10807 );
   or U11046 ( n10807,n10741,n7827 );
   nand U11047 ( n9481,datai_25_,n10742 );
   or U11048 ( n10806,n10743,n8793 );
   nand U11049 ( n9482,n10744,n10808 );
   nor U11050 ( n10804,n9478,n10746 );
   nand U11051 ( n9478,datai_17_,n10742 );
   nor U11052 ( n10802,n10809,n10810 );
   nor U11053 ( n10810,n10749,n10811 );
   nor U11054 ( n10809,n10751,n10708 );
   nand U11055 ( n10708,datai_1_,n9505 );
   nor U11056 ( n10813,n10814,n10815 );
   nand U11057 ( n10815,n10816,n10817 );
   or U11058 ( n10817,n10741,n8767 );
   nand U11059 ( n9517,datai_24_,n10742 );
   or U11060 ( n10816,n10743,n8814 );
   nand U11061 ( n9519,n10744,n10818 );
   nor U11062 ( n10744,n9602,n9018 );
   nor U11063 ( n10814,n9512,n10746 );
   nand U11064 ( n9512,datai_16_,n10742 );
   nor U11065 ( n10812,n10819,n10820 );
   nor U11066 ( n10820,n10751,n10721 );
   nand U11067 ( n10721,datai_0_,n9505 );
   and U11068 ( n10751,n10821,n10822 );
   nand U11069 ( n10822,n10384,n9946 );
   nor U11070 ( n9946,n9958,n8871 );
   not U11071 ( n10384,n10468 );
   nand U11072 ( n10821,n9493,n10823 );
   not U11073 ( n10823,n10824 );
   nand U11074 ( n9493,n10209,n8922 );
   nor U11075 ( n10819,n10749,n10825 );
   and U11076 ( n10749,n10826,n10827 );
   nand U11077 ( n10827,state2_reg_3_,n10743 );
   nand U11078 ( n10743,n10558,n9787 );
   nor U11079 ( n9787,instqueuewr_addr_reg_1_,instqueuewr_addr_reg_0_ );
   nor U11080 ( n10558,instqueuewr_addr_reg_3_,instqueuewr_addr_reg_2_ );
   nor U11081 ( n10826,n10828,n10829 );
   nor U11082 ( n10829,n10830,n10831 );
   nand U11083 ( n10831,n10832,n9502 );
   nand U11084 ( n9502,n10208,n9505 );
   nor U11085 ( n10208,n8916,n10742 );
   nor U11086 ( n10742,n9602,n8922 );
   nand U11087 ( n8922,statebs16_reg,n8857 );
   not U11088 ( n8916,n10209 );
   nand U11089 ( n10832,n9503,n10833 );
   nand U11090 ( n10833,n10741,n10746 );
   nand U11091 ( n10746,n10553,n9780 );
   nor U11092 ( n9780,n8905,n8917 );
   nor U11093 ( n10553,n8930,n8944 );
   nand U11094 ( n10741,n10556,n9785 );
   nor U11095 ( n9785,n10734,n10642 );
   not U11096 ( n10734,n10557 );
   nor U11097 ( n10557,n9607,n9695 );
   nor U11098 ( n9695,n8917,n10642 );
   nor U11099 ( n9607,n8905,n10834 );
   nor U11100 ( n10556,n9518,n8937 );
   xor U11101 ( n8937,n9514,n8930 );
   nand U11102 ( n9518,n10835,n10836 );
   or U11103 ( n10836,n9781,n9514 );
   nor U11104 ( n10835,n9872,n10837 );
   not U11105 ( n10837,n10139 );
   nand U11106 ( n10139,n10298,n9514 );
   nor U11107 ( n9514,n10834,n10642 );
   nor U11108 ( n10298,n8944,n9782 );
   nor U11109 ( n9872,n9781,n8930 );
   not U11110 ( n9503,n9777 );
   nand U11111 ( n9777,n9505,n10209 );
   nand U11112 ( n10209,n8857,n10838 );
   nor U11113 ( n10830,n10824,n9602 );
   nand U11114 ( n10824,n10551,n8920 );
   nor U11115 ( n10551,n10123,n10466 );
   nor U11116 ( n10828,n10839,n8790 );
   nor U11117 ( n10839,n9958,n10468 );
   nand U11118 ( n10468,n10639,n10126 );
   and U11119 ( u3019,instqueuewr_addr_reg_4_,n8900 );
   not U11120 ( n8900,n8902 );
   nand U11121 ( n8902,n10840,n10841 );
   nand U11122 ( n10841,n10842,n8908 );
   nand U11123 ( n8908,n9373,n10843 );
   nand U11124 ( n10843,n10844,n9375 );
   nand U11125 ( n9375,n10845,n10846 );
   nand U11126 ( n10846,n10847,instqueuerd_addr_reg_3_ );
   nand U11127 ( n10845,n9368,n8948 );
   nand U11128 ( n9368,n10848,n10849 );
   nand U11129 ( n10849,n9014,instqueuerd_addr_reg_3_ );
   nand U11130 ( n10848,n9004,n9340 );
   nand U11131 ( n9004,n10850,n10851 );
   nor U11132 ( n10851,n10852,n10853 );
   nor U11133 ( n10853,n10854,n10855 );
   nor U11134 ( n10852,n10856,n10857 );
   nor U11135 ( n10856,n10858,n10859 );
   nor U11136 ( n10859,instqueuerd_addr_reg_3_,n10860 );
   nor U11137 ( n10860,n10861,n10862 );
   nor U11138 ( n10858,n10861,n10863 );
   nand U11139 ( n10863,n10862,n10864 );
   nor U11140 ( n10850,n10865,n10866 );
   nor U11141 ( n10866,n9350,n10867 );
   nor U11142 ( n10865,n9364,n8947 );
   not U11143 ( n8947,n10466 );
   and U11144 ( n10844,n10868,n9376 );
   nand U11145 ( n9376,n10869,n10870 );
   nand U11146 ( n10870,n10871,n9327 );
   nand U11147 ( n9327,n9014,n10864 );
   nor U11148 ( n10871,state2_reg_1_,n9328 );
   and U11149 ( n9328,n8992,n9340 );
   and U11150 ( n8992,n10872,n10873 );
   nor U11151 ( n10873,n10874,n10875 );
   nor U11152 ( n10875,n10857,n8989 );
   nor U11153 ( n10857,n10876,n10877 );
   nor U11154 ( n10874,n10878,n10855 );
   nand U11155 ( n10855,n10879,n10880 );
   nor U11156 ( n10879,n10808,n10881 );
   nor U11157 ( n10872,n10882,n10883 );
   nor U11158 ( n10883,n10884,n9350 );
   nor U11159 ( n10882,n9364,n8933 );
   not U11160 ( n9364,n9349 );
   nand U11161 ( n9349,n10885,n10886 );
   nor U11162 ( n10886,n10887,n10888 );
   nand U11163 ( n10888,n10889,n10890 );
   not U11164 ( n10887,n10891 );
   nor U11165 ( n10885,n10892,n10893 );
   nand U11166 ( n10893,n10894,n10745 );
   nand U11167 ( n10869,n10847,instqueuerd_addr_reg_2_ );
   and U11168 ( n9373,n10895,n10896 );
   nand U11169 ( n10896,n10897,n8948 );
   nand U11170 ( n10897,n9009,n10898 );
   nand U11171 ( n10898,n9014,instqueuerd_addr_reg_4_ );
   not U11172 ( n9014,n9340 );
   nand U11173 ( n9340,n10899,n10900 );
   nor U11174 ( n10900,n10901,n10902 );
   nand U11175 ( n10902,n10903,n10904 );
   nand U11176 ( n10903,n10905,n9391 );
   nor U11177 ( n10905,n10906,n10798 );
   nor U11178 ( n10901,ready_n,n10907 );
   nor U11179 ( n10907,n10908,n10909 );
   nor U11180 ( n10909,n9380,n10889 );
   nor U11181 ( n10908,n9393,n10910 );
   nor U11182 ( n10910,n10911,n10912 );
   nor U11183 ( n10911,n10913,n8867 );
   nor U11184 ( n10913,n8961,n10914 );
   nor U11185 ( n10899,n10915,n10916 );
   nand U11186 ( n10916,n10917,n10918 );
   nand U11187 ( n10918,n10876,n9384 );
   nand U11188 ( n9009,n9379,n10919 );
   nand U11189 ( n10895,n10847,instqueuerd_addr_reg_4_ );
   nor U11190 ( n10847,n8948,flush_reg );
   nor U11191 ( n10840,n9012,n9505 );
   not U11192 ( n9505,n9602 );
   nand U11193 ( n9602,n8821,n10920 );
   nand U11194 ( n10920,n10921,n9273 );
   nand U11195 ( n9273,state2_reg_1_,n8789 );
   nor U11196 ( n10921,n9275,n8969 );
   nor U11197 ( n8969,n9018,n9393 );
   and U11198 ( n9012,flush_reg,n10842 );
   not U11199 ( n10842,n9295 );
   nand U11200 ( n9295,n9020,state2_reg_0_ );
   nor U11201 ( n10923,n10924,n10925 );
   nor U11202 ( n10925,n8889,n10926 );
   nor U11203 ( n10924,n8812,n10928 );
   nor U11204 ( n10922,n10929,n10930 );
   nand U11205 ( n10930,n10931,n10932 );
   nand U11206 ( n10931,instaddrpointer_reg_0_,n10933 );
   nand U11207 ( n10933,n10934,n8800 );
   nor U11208 ( n10929,n8751,n10936 );
   nor U11209 ( n10938,n10939,n10940 );
   nand U11210 ( n10940,n10941,n10942 );
   or U11211 ( n10941,n10943,n8812 );
   nor U11212 ( n10939,n9192,n10926 );
   nor U11213 ( n10937,n10944,n10945 );
   nand U11214 ( n10945,n10946,n10947 );
   nand U11215 ( n10947,instaddrpointer_reg_1_,n10948 );
   nand U11216 ( n10948,n10934,n10932 );
   nand U11217 ( n10932,n10949,n8965 );
   nand U11218 ( n10946,n10950,n8996 );
   nor U11219 ( n10950,n8792,n8965 );
   nor U11220 ( n10944,n8752,n10952 );
   nor U11221 ( n10954,n10955,n10956 );
   nand U11222 ( n10956,n10957,n10958 );
   nand U11223 ( n10958,n10959,n10960 );
   nand U11224 ( n10960,n10961,n10962 );
   nand U11225 ( n10957,n10963,n8779 );
   nor U11226 ( n10955,n9187,n8739 );
   nor U11227 ( n10953,n10965,n10966 );
   nand U11228 ( n10966,n10967,n10968 );
   nand U11229 ( n10968,instaddrpointer_reg_2_,n10969 );
   nand U11230 ( n10969,n10970,n10971 );
   nand U11231 ( n10971,n10972,n10973 );
   nor U11232 ( n10970,n10974,n10975 );
   nand U11233 ( n10967,n10976,n10977 );
   nor U11234 ( n10976,n10978,n8996 );
   nor U11235 ( n10978,n10979,n10980 );
   nor U11236 ( n10979,n8965,n8775 );
   nor U11237 ( n10965,n8754,n10982 );
   nor U11238 ( n10984,n10985,n10986 );
   nor U11239 ( n10986,n9182,n8740 );
   nor U11240 ( n10985,n10987,n10988 );
   nand U11241 ( n10988,n10989,n8779 );
   nor U11242 ( n10983,n10990,n10991 );
   nand U11243 ( n10991,n10992,n10993 );
   nand U11244 ( n10993,instaddrpointer_reg_3_,n10994 );
   nand U11245 ( n10994,n10995,n10996 );
   nor U11246 ( n10995,n10975,n10997 );
   nor U11247 ( n10997,instaddrpointer_reg_2_,n8800 );
   not U11248 ( n10975,n10942 );
   nand U11249 ( n10942,n10980,n8996 );
   nand U11250 ( n10992,n10998,n10999 );
   nand U11251 ( n10998,n11000,n11001 );
   nand U11252 ( n11001,n11002,instaddrpointer_reg_2_ );
   nor U11253 ( n11002,n8996,n8800 );
   not U11254 ( n11000,n11003 );
   nor U11255 ( n10990,n8754,n11004 );
   nor U11256 ( n11006,n11007,n11008 );
   nor U11257 ( n11008,n9177,n10926 );
   nor U11258 ( n11007,n11009,n11010 );
   nand U11259 ( n11010,n11011,n8779 );
   nor U11260 ( n11005,n11012,n11013 );
   nand U11261 ( n11013,n11014,n11015 );
   nand U11262 ( n11015,instaddrpointer_reg_4_,n11016 );
   nand U11263 ( n11016,n11017,n10996 );
   and U11264 ( n10996,n11018,n11019 );
   nand U11265 ( n11019,n11020,n10959 );
   nor U11266 ( n11018,n10974,n11021 );
   nor U11267 ( n11021,n11022,n10981 );
   nor U11268 ( n11017,n11023,n11024 );
   nor U11269 ( n11024,instaddrpointer_reg_3_,n10951 );
   nor U11270 ( n11023,n11025,n8800 );
   nand U11271 ( n11014,n11026,n11027 );
   nand U11272 ( n11026,n11028,n11029 );
   nand U11273 ( n11029,instaddrpointer_reg_3_,n11003 );
   nand U11274 ( n11003,n11030,n11031 );
   nand U11275 ( n11031,n11022,n10972 );
   not U11276 ( n11022,n10962 );
   nand U11277 ( n11030,n10959,n10961 );
   nand U11278 ( n11028,n11025,n8817 );
   nor U11279 ( n11012,n8751,n11032 );
   nor U11280 ( n11034,n11035,n11036 );
   nor U11281 ( n11036,n9172,n8739 );
   and U11282 ( n11035,n10964,n11037 );
   nor U11283 ( n11033,n11038,n11039 );
   nand U11284 ( n11039,n11040,n11041 );
   nand U11285 ( n11041,instaddrpointer_reg_5_,n11042 );
   nand U11286 ( n11042,n11043,n11044 );
   nand U11287 ( n11044,n10980,n11045 );
   nand U11288 ( n11040,n11046,n11047 );
   nand U11289 ( n11046,n11048,n11049 );
   or U11290 ( n11049,n11045,n10935 );
   not U11291 ( n11048,n11050 );
   nor U11292 ( n11038,n8751,n11051 );
   nor U11293 ( n11053,n11054,n11055 );
   nor U11294 ( n11055,n9167,n8740 );
   and U11295 ( n11054,n8779,n11056 );
   nor U11296 ( n11052,n11057,n11058 );
   nand U11297 ( n11058,n11059,n11060 );
   nand U11298 ( n11060,instaddrpointer_reg_6_,n11061 );
   nand U11299 ( n11061,n11062,n11043 );
   and U11300 ( n11043,n11063,n11064 );
   nand U11301 ( n11064,n10959,n11065 );
   nor U11302 ( n11063,n10974,n11066 );
   nor U11303 ( n11066,n11067,n8775 );
   nor U11304 ( n11062,n11068,n11069 );
   nor U11305 ( n11069,instaddrpointer_reg_5_,n10951 );
   nor U11306 ( n11068,n11070,n10935 );
   nand U11307 ( n11059,n11071,n11072 );
   not U11308 ( n11072,instaddrpointer_reg_6_ );
   nand U11309 ( n11071,n11073,n11074 );
   nand U11310 ( n11074,instaddrpointer_reg_5_,n11050 );
   nand U11311 ( n11050,n11075,n11076 );
   nand U11312 ( n11076,n11067,n10972 );
   not U11313 ( n11067,n11077 );
   or U11314 ( n11075,n11065,n11078 );
   nand U11315 ( n11073,n11070,n8817 );
   nor U11316 ( n11057,n8753,n11079 );
   nor U11317 ( n11081,n11082,n11083 );
   nor U11318 ( n11083,n9162,n10926 );
   and U11319 ( n11082,n10964,n11084 );
   nor U11320 ( n11080,n11085,n11086 );
   nand U11321 ( n11086,n11087,n11088 );
   nand U11322 ( n11088,instaddrpointer_reg_7_,n11089 );
   nand U11323 ( n11089,n11090,n11091 );
   nand U11324 ( n11091,n10980,n11092 );
   nand U11325 ( n11087,n11093,n11094 );
   nand U11326 ( n11093,n11095,n11096 );
   or U11327 ( n11096,n11092,n10935 );
   not U11328 ( n11095,n11097 );
   nor U11329 ( n11085,n8753,n11098 );
   nor U11330 ( n11100,n11101,n11102 );
   nor U11331 ( n11102,n9157,n8739 );
   nor U11332 ( n11101,n10927,n11103 );
   nor U11333 ( n11099,n11104,n11105 );
   nand U11334 ( n11105,n11106,n11107 );
   nand U11335 ( n11107,instaddrpointer_reg_8_,n11108 );
   nand U11336 ( n11108,n11109,n11090 );
   and U11337 ( n11090,n11110,n11111 );
   nand U11338 ( n11111,n10959,n11112 );
   nor U11339 ( n11110,n8816,n11113 );
   nor U11340 ( n11113,n11114,n10981 );
   nor U11341 ( n11109,n11115,n11116 );
   nor U11342 ( n11116,instaddrpointer_reg_7_,n10951 );
   nor U11343 ( n11115,n11117,n10935 );
   nand U11344 ( n11106,n11118,n11119 );
   nand U11345 ( n11118,n11120,n11121 );
   nand U11346 ( n11121,instaddrpointer_reg_7_,n11097 );
   nand U11347 ( n11097,n11122,n11123 );
   nand U11348 ( n11123,n11114,n10972 );
   not U11349 ( n11114,n11124 );
   or U11350 ( n11122,n11112,n11078 );
   nand U11351 ( n11120,n11117,n8817 );
   nor U11352 ( n11104,n8752,n11125 );
   nor U11353 ( n11127,n11128,n11129 );
   nor U11354 ( n11129,n9152,n8740 );
   and U11355 ( n11128,n10964,n11130 );
   nor U11356 ( n11126,n11131,n11132 );
   nand U11357 ( n11132,n11133,n11134 );
   nand U11358 ( n11134,instaddrpointer_reg_9_,n11135 );
   nand U11359 ( n11135,n11136,n11137 );
   nand U11360 ( n11137,n10980,n11138 );
   nand U11361 ( n11133,n11139,n11140 );
   nand U11362 ( n11139,n11141,n11142 );
   or U11363 ( n11142,n11138,n8800 );
   not U11364 ( n11141,n11143 );
   nor U11365 ( n11131,n8752,n11144 );
   nor U11366 ( n11146,n11147,n11148 );
   nor U11367 ( n11148,n9147,n10926 );
   nor U11368 ( n11147,n8812,n11149 );
   nor U11369 ( n11145,n11150,n11151 );
   nand U11370 ( n11151,n11152,n11153 );
   nand U11371 ( n11153,instaddrpointer_reg_10_,n11154 );
   nand U11372 ( n11154,n11155,n11136 );
   and U11373 ( n11136,n11156,n11157 );
   nand U11374 ( n11157,n10959,n11158 );
   nor U11375 ( n11156,n10974,n11159 );
   nor U11376 ( n11159,n11160,n10981 );
   nor U11377 ( n11155,n11161,n11162 );
   nor U11378 ( n11162,instaddrpointer_reg_9_,n10951 );
   nor U11379 ( n11161,n11163,n8800 );
   nand U11380 ( n11152,n11164,n11165 );
   nand U11381 ( n11164,n11166,n11167 );
   nand U11382 ( n11167,instaddrpointer_reg_9_,n11143 );
   nand U11383 ( n11143,n11168,n11169 );
   nand U11384 ( n11169,n11160,n10972 );
   not U11385 ( n11160,n11170 );
   or U11386 ( n11168,n11158,n11078 );
   nand U11387 ( n11166,n11163,n8817 );
   nor U11388 ( n11150,n8754,n11171 );
   nor U11389 ( n11173,n11174,n11175 );
   nor U11390 ( n11175,n9142,n8739 );
   and U11391 ( n11174,n10964,n11176 );
   nor U11392 ( n11172,n11177,n11178 );
   nand U11393 ( n11178,n11179,n11180 );
   nand U11394 ( n11180,instaddrpointer_reg_11_,n11181 );
   nand U11395 ( n11181,n11182,n11183 );
   nand U11396 ( n11183,n10980,n11184 );
   nand U11397 ( n11179,n11185,n11186 );
   nand U11398 ( n11185,n11187,n11188 );
   or U11399 ( n11188,n11184,n8800 );
   not U11400 ( n11187,n11189 );
   nor U11401 ( n11177,n8754,n11190 );
   nor U11402 ( n11192,n11193,n11194 );
   nor U11403 ( n11194,n9137,n8740 );
   nor U11404 ( n11193,n8812,n11195 );
   nor U11405 ( n11191,n11196,n11197 );
   nand U11406 ( n11197,n11198,n11199 );
   nand U11407 ( n11199,instaddrpointer_reg_12_,n11200 );
   nand U11408 ( n11200,n11201,n11182 );
   and U11409 ( n11182,n11202,n11203 );
   nand U11410 ( n11203,n10959,n11204 );
   nor U11411 ( n11202,n10974,n11205 );
   nor U11412 ( n11205,n11206,n10981 );
   nor U11413 ( n11201,n11207,n11208 );
   nor U11414 ( n11208,instaddrpointer_reg_11_,n10951 );
   nor U11415 ( n11207,n11209,n10935 );
   nand U11416 ( n11198,n11210,n11211 );
   nand U11417 ( n11210,n11212,n11213 );
   nand U11418 ( n11213,instaddrpointer_reg_11_,n11189 );
   nand U11419 ( n11189,n11214,n11215 );
   nand U11420 ( n11215,n11206,n10972 );
   not U11421 ( n11206,n11216 );
   or U11422 ( n11214,n11204,n11078 );
   nand U11423 ( n11212,n11209,n8817 );
   nor U11424 ( n11196,n8752,n11217 );
   nor U11425 ( n11219,n11220,n11221 );
   nor U11426 ( n11221,n9132,n8739 );
   nor U11427 ( n11220,n10927,n11222 );
   nor U11428 ( n11218,n11223,n11224 );
   nand U11429 ( n11224,n11225,n11226 );
   nand U11430 ( n11226,instaddrpointer_reg_13_,n11227 );
   nand U11431 ( n11227,n11228,n11229 );
   nand U11432 ( n11229,n10980,n11230 );
   nand U11433 ( n11225,n11231,n11232 );
   nand U11434 ( n11231,n11233,n11234 );
   or U11435 ( n11234,n11230,n10935 );
   not U11436 ( n11233,n11235 );
   nor U11437 ( n11223,n8753,n11236 );
   nor U11438 ( n11238,n11239,n11240 );
   nor U11439 ( n11240,n9127,n10926 );
   nor U11440 ( n11239,n10927,n11241 );
   nor U11441 ( n11237,n11242,n11243 );
   nand U11442 ( n11243,n11244,n11245 );
   nand U11443 ( n11245,instaddrpointer_reg_14_,n11246 );
   nand U11444 ( n11246,n11247,n11228 );
   and U11445 ( n11228,n11248,n11249 );
   nand U11446 ( n11249,n10959,n11250 );
   nor U11447 ( n11248,n10974,n11251 );
   nor U11448 ( n11251,n11252,n10981 );
   nor U11449 ( n11247,n11253,n11254 );
   nor U11450 ( n11254,instaddrpointer_reg_13_,n10951 );
   nor U11451 ( n11253,n11255,n10935 );
   nand U11452 ( n11244,n11256,n11257 );
   nand U11453 ( n11256,n11258,n11259 );
   nand U11454 ( n11259,instaddrpointer_reg_13_,n11235 );
   nand U11455 ( n11235,n11260,n11261 );
   nand U11456 ( n11261,n11252,n10972 );
   not U11457 ( n11252,n11262 );
   or U11458 ( n11260,n11250,n11078 );
   nand U11459 ( n11258,n11255,n8817 );
   nor U11460 ( n11242,n8753,n11263 );
   nor U11461 ( n11265,n11266,n11267 );
   nor U11462 ( n11267,n9122,n8740 );
   nor U11463 ( n11266,n10927,n11268 );
   nor U11464 ( n11264,n11269,n11270 );
   nand U11465 ( n11270,n11271,n11272 );
   nand U11466 ( n11272,instaddrpointer_reg_15_,n11273 );
   nand U11467 ( n11273,n11274,n11275 );
   nand U11468 ( n11275,n10980,n11276 );
   nand U11469 ( n11271,n11277,n11278 );
   nand U11470 ( n11277,n11279,n11280 );
   or U11471 ( n11280,n11276,n10935 );
   not U11472 ( n11279,n11281 );
   nor U11473 ( n11269,n8751,n11282 );
   nor U11474 ( n11284,n11285,n11286 );
   nor U11475 ( n11286,n9117,n8739 );
   nor U11476 ( n11285,n10927,n11287 );
   nor U11477 ( n11283,n11288,n11289 );
   nand U11478 ( n11289,n11290,n11291 );
   nand U11479 ( n11291,instaddrpointer_reg_16_,n11292 );
   nand U11480 ( n11292,n11293,n11274 );
   and U11481 ( n11274,n11294,n11295 );
   nand U11482 ( n11295,n10959,n11296 );
   nor U11483 ( n11294,n10974,n11297 );
   nor U11484 ( n11297,n11298,n10981 );
   nor U11485 ( n11293,n11299,n11300 );
   nor U11486 ( n11300,instaddrpointer_reg_15_,n10951 );
   nor U11487 ( n11299,n11301,n10935 );
   nand U11488 ( n11290,n11302,n11303 );
   not U11489 ( n11303,instaddrpointer_reg_16_ );
   nand U11490 ( n11302,n11304,n11305 );
   nand U11491 ( n11305,instaddrpointer_reg_15_,n11281 );
   nand U11492 ( n11281,n11306,n11307 );
   nand U11493 ( n11307,n11298,n10972 );
   not U11494 ( n11298,n11308 );
   or U11495 ( n11306,n11296,n11078 );
   nand U11496 ( n11304,n11301,n8817 );
   nor U11497 ( n11288,n8751,n11309 );
   nor U11498 ( n11311,n11312,n11313 );
   nor U11499 ( n11313,n9112,n10926 );
   and U11500 ( n11312,n10964,n11314 );
   nor U11501 ( n11310,n11315,n11316 );
   nand U11502 ( n11316,n11317,n11318 );
   nand U11503 ( n11318,instaddrpointer_reg_17_,n11319 );
   nand U11504 ( n11319,n11320,n11321 );
   nand U11505 ( n11321,n10980,n11322 );
   nand U11506 ( n11317,n11323,n11324 );
   nand U11507 ( n11323,n11325,n11326 );
   or U11508 ( n11326,n11322,n8800 );
   not U11509 ( n11325,n11327 );
   nor U11510 ( n11315,n8754,n11328 );
   nor U11511 ( n11330,n11331,n11332 );
   nor U11512 ( n11332,n9107,n8740 );
   and U11513 ( n11331,n10964,n11333 );
   nor U11514 ( n11329,n11334,n11335 );
   nand U11515 ( n11335,n11336,n11337 );
   nand U11516 ( n11337,instaddrpointer_reg_18_,n11338 );
   nand U11517 ( n11338,n11339,n11320 );
   and U11518 ( n11320,n11340,n11341 );
   nand U11519 ( n11341,n10959,n11342 );
   nor U11520 ( n11340,n10974,n11343 );
   nor U11521 ( n11343,n11344,n10981 );
   nor U11522 ( n11339,n11345,n11346 );
   nor U11523 ( n11346,instaddrpointer_reg_17_,n10951 );
   nor U11524 ( n11345,n11347,n8800 );
   nand U11525 ( n11336,n11348,n11349 );
   nand U11526 ( n11348,n11350,n11351 );
   nand U11527 ( n11351,instaddrpointer_reg_17_,n11327 );
   nand U11528 ( n11327,n11352,n11353 );
   nand U11529 ( n11353,n11344,n10972 );
   not U11530 ( n11344,n11354 );
   or U11531 ( n11352,n11342,n11078 );
   nand U11532 ( n11350,n11347,n10980 );
   nor U11533 ( n11334,n8754,n11355 );
   nor U11534 ( n11357,n11358,n11359 );
   nor U11535 ( n11359,n9102,n8739 );
   nor U11536 ( n11358,n10927,n11360 );
   nor U11537 ( n11356,n11361,n11362 );
   nand U11538 ( n11362,n11363,n11364 );
   nand U11539 ( n11364,instaddrpointer_reg_19_,n11365 );
   nand U11540 ( n11365,n11366,n11367 );
   nand U11541 ( n11367,n10980,n11368 );
   nand U11542 ( n11363,n11369,n11370 );
   nand U11543 ( n11369,n11371,n11372 );
   or U11544 ( n11372,n11368,n8800 );
   not U11545 ( n11371,n11373 );
   nor U11546 ( n11361,n8752,n11374 );
   nor U11547 ( n11376,n11377,n11378 );
   nor U11548 ( n11378,n9097,n10926 );
   nor U11549 ( n11377,n11379,n11380 );
   nand U11550 ( n11380,n11381,n8779 );
   nor U11551 ( n11375,n11382,n11383 );
   nand U11552 ( n11383,n11384,n11385 );
   nand U11553 ( n11385,instaddrpointer_reg_20_,n11386 );
   nand U11554 ( n11386,n11387,n11366 );
   and U11555 ( n11366,n11388,n11389 );
   nand U11556 ( n11389,n10959,n11390 );
   nor U11557 ( n11388,n10974,n11391 );
   nor U11558 ( n11391,n11392,n10981 );
   nor U11559 ( n11387,n11393,n11394 );
   nor U11560 ( n11394,instaddrpointer_reg_19_,n10951 );
   nor U11561 ( n11393,n11395,n10935 );
   nand U11562 ( n11384,n11396,n11397 );
   nand U11563 ( n11396,n11398,n11399 );
   nand U11564 ( n11399,instaddrpointer_reg_19_,n11373 );
   nand U11565 ( n11373,n11400,n11401 );
   nand U11566 ( n11401,n11392,n10972 );
   not U11567 ( n11392,n11402 );
   or U11568 ( n11400,n11390,n11078 );
   nand U11569 ( n11398,n11395,n8817 );
   nor U11570 ( n11382,n8752,n11403 );
   nor U11571 ( n11405,n11406,n11407 );
   nor U11572 ( n11407,n9092,n8739 );
   and U11573 ( n11406,n10964,n11408 );
   nor U11574 ( n11404,n11409,n11410 );
   nand U11575 ( n11410,n11411,n11412 );
   nand U11576 ( n11412,instaddrpointer_reg_21_,n11413 );
   nand U11577 ( n11413,n11414,n11415 );
   nand U11578 ( n11415,n10980,n11416 );
   nand U11579 ( n11411,n11417,n11418 );
   nand U11580 ( n11417,n11419,n11420 );
   or U11581 ( n11420,n11416,n8800 );
   not U11582 ( n11419,n11421 );
   nor U11583 ( n11409,n8751,n11422 );
   nor U11584 ( n11424,n11425,n11426 );
   nor U11585 ( n11426,n9087,n8740 );
   and U11586 ( n11425,n8779,n11427 );
   nor U11587 ( n11423,n11428,n11429 );
   nand U11588 ( n11429,n11430,n11431 );
   nand U11589 ( n11431,instaddrpointer_reg_22_,n11432 );
   nand U11590 ( n11432,n11433,n11414 );
   and U11591 ( n11414,n11434,n11435 );
   nand U11592 ( n11435,n10959,n11436 );
   nor U11593 ( n11434,n10974,n11437 );
   nor U11594 ( n11437,n11438,n10981 );
   nor U11595 ( n11433,n11439,n11440 );
   nor U11596 ( n11440,instaddrpointer_reg_21_,n10951 );
   nor U11597 ( n11439,n11441,n8800 );
   nand U11598 ( n11430,n11442,n11443 );
   nand U11599 ( n11442,n11444,n11445 );
   nand U11600 ( n11445,instaddrpointer_reg_21_,n11421 );
   nand U11601 ( n11421,n11446,n11447 );
   nand U11602 ( n11447,n11438,n10972 );
   or U11603 ( n11446,n11436,n11078 );
   nand U11604 ( n11444,n11441,n8817 );
   nor U11605 ( n11428,n8753,n11448 );
   nor U11606 ( n11450,n11451,n11452 );
   nor U11607 ( n11452,n9082,n10926 );
   and U11608 ( n11451,n10964,n11453 );
   nor U11609 ( n11449,n11454,n11455 );
   nand U11610 ( n11455,n11456,n11457 );
   nand U11611 ( n11457,instaddrpointer_reg_23_,n11458 );
   nand U11612 ( n11458,n11459,n11460 );
   nand U11613 ( n11460,n10980,n11461 );
   nand U11614 ( n11456,n11462,n11463 );
   nand U11615 ( n11462,n11464,n11465 );
   or U11616 ( n11465,n11461,n10935 );
   not U11617 ( n11464,n11466 );
   nor U11618 ( n11454,n8753,n11467 );
   nor U11619 ( n11469,n11470,n11471 );
   nor U11620 ( n11471,n9077,n8739 );
   and U11621 ( n11470,n10964,n11472 );
   nor U11622 ( n11468,n11473,n11474 );
   nand U11623 ( n11474,n11475,n11476 );
   nand U11624 ( n11476,instaddrpointer_reg_24_,n11477 );
   nand U11625 ( n11477,n11478,n11459 );
   and U11626 ( n11459,n11479,n11480 );
   nand U11627 ( n11480,n10959,n11481 );
   nor U11628 ( n11479,n8816,n11482 );
   nor U11629 ( n11482,n11483,n10981 );
   nor U11630 ( n11478,n11484,n11485 );
   nor U11631 ( n11485,instaddrpointer_reg_23_,n10951 );
   nor U11632 ( n11484,n11486,n10935 );
   nand U11633 ( n11475,n11487,n11488 );
   nand U11634 ( n11487,n11489,n11490 );
   nand U11635 ( n11490,instaddrpointer_reg_23_,n11466 );
   nand U11636 ( n11466,n11491,n11492 );
   nand U11637 ( n11492,n11483,n10972 );
   not U11638 ( n11483,n11493 );
   nand U11639 ( n11491,n11494,n10959 );
   nand U11640 ( n11489,n11486,n8817 );
   nor U11641 ( n11473,n8752,n11495 );
   nor U11642 ( n11497,n11498,n11499 );
   nor U11643 ( n11499,n9072,n8740 );
   and U11644 ( n11498,n10964,n11500 );
   nor U11645 ( n11496,n11501,n11502 );
   nand U11646 ( n11502,n11503,n11504 );
   nand U11647 ( n11504,instaddrpointer_reg_25_,n11505 );
   nand U11648 ( n11505,n11506,n11507 );
   nand U11649 ( n11507,n10980,n11508 );
   nand U11650 ( n11503,n11509,n11510 );
   nand U11651 ( n11509,n11511,n11512 );
   or U11652 ( n11512,n11508,n8800 );
   not U11653 ( n11511,n11513 );
   nor U11654 ( n11501,n8752,n11514 );
   nor U11655 ( n11516,n11517,n11518 );
   nor U11656 ( n11518,n9067,n10926 );
   nor U11657 ( n11517,n10927,n11519 );
   nor U11658 ( n11515,n11520,n11521 );
   nand U11659 ( n11521,n11522,n11523 );
   nand U11660 ( n11523,instaddrpointer_reg_26_,n11524 );
   nand U11661 ( n11524,n11525,n11506 );
   and U11662 ( n11506,n11526,n11527 );
   nand U11663 ( n11527,n10959,n11528 );
   nor U11664 ( n11526,n8816,n11529 );
   nor U11665 ( n11529,n11530,n10981 );
   nor U11666 ( n11525,n11531,n11532 );
   nor U11667 ( n11532,instaddrpointer_reg_25_,n10951 );
   nor U11668 ( n11531,n11533,n10935 );
   nand U11669 ( n11522,n11534,n11535 );
   nand U11670 ( n11534,n11536,n11537 );
   nand U11671 ( n11537,instaddrpointer_reg_25_,n11513 );
   nand U11672 ( n11513,n11538,n11539 );
   nand U11673 ( n11539,n11530,n10972 );
   not U11674 ( n11530,n11540 );
   or U11675 ( n11538,n11528,n11078 );
   nand U11676 ( n11536,n11533,n8817 );
   nor U11677 ( n11520,n8754,n11541 );
   nor U11678 ( n11543,n11544,n11545 );
   nor U11679 ( n11545,n9062,n8739 );
   and U11680 ( n11544,n10964,n11546 );
   nor U11681 ( n11542,n11547,n11548 );
   nand U11682 ( n11548,n11549,n11550 );
   nand U11683 ( n11550,instaddrpointer_reg_27_,n11551 );
   nand U11684 ( n11551,n11552,n11553 );
   nand U11685 ( n11553,n10980,n11554 );
   nand U11686 ( n11549,n11555,n11556 );
   nand U11687 ( n11555,n11557,n11558 );
   or U11688 ( n11558,n11554,n10935 );
   nor U11689 ( n11547,n8754,n11559 );
   nor U11690 ( n11561,n11562,n11563 );
   nor U11691 ( n11563,n9057,n8740 );
   nor U11692 ( n11562,n10927,n11564 );
   nor U11693 ( n11560,n11565,n11566 );
   nand U11694 ( n11566,n11567,n11568 );
   nand U11695 ( n11568,instaddrpointer_reg_28_,n11569 );
   nand U11696 ( n11569,n11570,n11552 );
   and U11697 ( n11552,n11571,n11572 );
   nand U11698 ( n11572,n10959,n11573 );
   not U11699 ( n10959,n11078 );
   nor U11700 ( n11571,n8816,n11574 );
   nor U11701 ( n11574,n11575,n10981 );
   nor U11702 ( n11570,n11576,n11577 );
   nor U11703 ( n11577,instaddrpointer_reg_27_,n10951 );
   nor U11704 ( n11576,n11578,n8800 );
   nand U11705 ( n11567,n11579,n11580 );
   nand U11706 ( n11579,n11581,n11582 );
   nand U11707 ( n11582,instaddrpointer_reg_27_,n11583 );
   nand U11708 ( n11581,n11578,n8817 );
   not U11709 ( n10980,n8800 );
   nor U11710 ( n11565,n8751,n11584 );
   nor U11711 ( n11586,n11587,n11588 );
   nor U11712 ( n11588,n9052,n10926 );
   and U11713 ( n11587,n10964,n11589 );
   nor U11714 ( n11585,n11590,n11591 );
   nand U11715 ( n11591,n11592,n11593 );
   nand U11716 ( n11593,instaddrpointer_reg_29_,n11594 );
   nand U11717 ( n11592,n11595,n11596 );
   nor U11718 ( n11590,n8751,n11597 );
   nor U11719 ( n11599,n11600,n11601 );
   nor U11720 ( n11601,n9047,n8739 );
   nor U11721 ( n11600,n10927,n11602 );
   nor U11722 ( n11598,n11603,n11604 );
   nand U11723 ( n11604,n11605,n11606 );
   or U11724 ( n11606,n11607,instaddrpointer_reg_30_ );
   or U11725 ( n11605,n11608,n11609 );
   nor U11726 ( n11603,n8753,n11610 );
   nor U11727 ( n11612,n11613,n11614 );
   nor U11728 ( n11614,n9045,n8740 );
   nand U11729 ( n10926,n8789,n10934 );
   nor U11730 ( n11613,n8812,n11615 );
   not U11731 ( n10927,n10964 );
   nand U11732 ( n10964,n11616,n11617 );
   nand U11733 ( n11617,n11618,n10778 );
   nand U11734 ( n11616,n11619,n11620 );
   nand U11735 ( n11620,n11621,n11622 );
   nor U11736 ( n11622,n9379,n10912 );
   not U11737 ( n9379,n10889 );
   nor U11738 ( n11621,n10876,n11623 );
   nor U11739 ( n11623,n11624,n11625 );
   nand U11740 ( n11625,n11626,n11627 );
   nand U11741 ( n11626,n11628,n11629 );
   nand U11742 ( n11629,n8757,n10818 );
   nand U11743 ( n11628,n8874,n10788 );
   not U11744 ( n11624,n9390 );
   not U11745 ( n10876,n9387 );
   nand U11746 ( n9387,n11630,n9367 );
   nor U11747 ( n11630,n11631,n11632 );
   nor U11748 ( n11611,n11633,n11634 );
   nand U11749 ( n11634,n11635,n11636 );
   nand U11750 ( n11636,instaddrpointer_reg_31_,n11637 );
   nand U11751 ( n11637,n11609,n11638 );
   nand U11752 ( n11638,n11639,n11608 );
   nor U11753 ( n11609,n11594,n11640 );
   and U11754 ( n11640,n11639,n11596 );
   nand U11755 ( n11639,n10951,n10935 );
   not U11756 ( n10951,n10949 );
   nand U11757 ( n10949,n11078,n8775 );
   nand U11758 ( n11594,n11641,n11642 );
   nor U11759 ( n11642,n8816,n11643 );
   nor U11760 ( n11643,n11644,n8800 );
   and U11761 ( n11644,instaddrpointer_reg_28_,n11578 );
   nor U11762 ( n11641,n11645,n11646 );
   nor U11763 ( n11646,n11647,n10981 );
   nor U11764 ( n11647,n11648,n11649 );
   nor U11765 ( n11645,n11650,n11078 );
   nor U11766 ( n11650,n11573,n11649 );
   nand U11767 ( n11635,n11651,n8997 );
   nor U11768 ( n11651,n11608,n11607 );
   nand U11769 ( n11607,instaddrpointer_reg_29_,n11595 );
   nand U11770 ( n11595,n11652,n11653 );
   nand U11771 ( n11653,n11654,n11578 );
   nor U11772 ( n11578,n11554,n11556 );
   nand U11773 ( n11554,n11533,instaddrpointer_reg_26_ );
   nor U11774 ( n11533,n11508,n11510 );
   nand U11775 ( n11508,n11486,instaddrpointer_reg_24_ );
   nor U11776 ( n11486,n11461,n11463 );
   nand U11777 ( n11461,n11441,instaddrpointer_reg_22_ );
   nor U11778 ( n11441,n11416,n11418 );
   nand U11779 ( n11416,n11395,instaddrpointer_reg_20_ );
   nor U11780 ( n11395,n11368,n11370 );
   nand U11781 ( n11368,n11347,instaddrpointer_reg_18_ );
   nor U11782 ( n11347,n11322,n11324 );
   nand U11783 ( n11322,n11301,instaddrpointer_reg_16_ );
   nor U11784 ( n11301,n11276,n11278 );
   nand U11785 ( n11276,n11255,instaddrpointer_reg_14_ );
   nor U11786 ( n11255,n11230,n11232 );
   nand U11787 ( n11230,n11209,instaddrpointer_reg_12_ );
   nor U11788 ( n11209,n11184,n11186 );
   nand U11789 ( n11184,n11163,instaddrpointer_reg_10_ );
   nor U11790 ( n11163,n11138,n11140 );
   nand U11791 ( n11138,n11117,instaddrpointer_reg_8_ );
   nor U11792 ( n11117,n11092,n11094 );
   nand U11793 ( n11092,n11070,instaddrpointer_reg_6_ );
   nor U11794 ( n11070,n11045,n11047 );
   nand U11795 ( n11045,n11025,instaddrpointer_reg_4_ );
   and U11796 ( n11025,n11655,instaddrpointer_reg_3_ );
   nor U11797 ( n11655,n8996,n10977 );
   nor U11798 ( n11654,n10935,n11580 );
   nand U11799 ( n10935,n11619,n8961 );
   or U11800 ( n11652,n11649,n11557 );
   not U11801 ( n11557,n11583 );
   nand U11802 ( n11583,n11656,n11657 );
   nand U11803 ( n11657,n11575,n10972 );
   not U11804 ( n10972,n10981 );
   nand U11805 ( n10981,n11619,n11658 );
   nand U11806 ( n11658,n11659,n11660 );
   nor U11807 ( n11660,n11661,n11662 );
   nor U11808 ( n11662,n10758,n11663 );
   nor U11809 ( n11659,n11664,n10892 );
   nand U11810 ( n10892,n11665,n11666 );
   nor U11811 ( n11666,n11667,n11668 );
   nand U11812 ( n11668,n11669,n11670 );
   nand U11813 ( n11667,n11671,n10904 );
   nand U11814 ( n10904,n11672,n10818 );
   nor U11815 ( n11665,n11673,n11674 );
   nand U11816 ( n11674,n11675,n11676 );
   nand U11817 ( n11676,n11677,n10808 );
   nand U11818 ( n11677,n11663,n11678 );
   nand U11819 ( n11678,n11679,n10798 );
   nand U11820 ( n11675,n10818,n10798 );
   nor U11821 ( n11673,n11680,n8758 );
   nor U11822 ( n11664,n10818,n10894 );
   not U11823 ( n11575,n11648 );
   nand U11824 ( n11648,n11681,instaddrpointer_reg_26_ );
   nor U11825 ( n11681,n11510,n11540 );
   nand U11826 ( n11540,n11682,instaddrpointer_reg_24_ );
   nor U11827 ( n11682,n11463,n11493 );
   nand U11828 ( n11493,n11683,n11438 );
   and U11829 ( n11438,n11684,instaddrpointer_reg_20_ );
   nor U11830 ( n11684,n11370,n11402 );
   nand U11831 ( n11402,n11685,instaddrpointer_reg_18_ );
   nor U11832 ( n11685,n11324,n11354 );
   nand U11833 ( n11354,n11686,instaddrpointer_reg_16_ );
   nor U11834 ( n11686,n11278,n11308 );
   nand U11835 ( n11308,n11687,instaddrpointer_reg_14_ );
   nor U11836 ( n11687,n11232,n11262 );
   nand U11837 ( n11262,n11688,instaddrpointer_reg_12_ );
   nor U11838 ( n11688,n11186,n11216 );
   nand U11839 ( n11216,n11689,instaddrpointer_reg_10_ );
   nor U11840 ( n11689,n11140,n11170 );
   nand U11841 ( n11170,n11690,instaddrpointer_reg_8_ );
   nor U11842 ( n11690,n11094,n11124 );
   nand U11843 ( n11124,n11691,instaddrpointer_reg_6_ );
   nor U11844 ( n11691,n11047,n11077 );
   nand U11845 ( n11077,n11692,instaddrpointer_reg_4_ );
   nor U11846 ( n11692,n10999,n10962 );
   nand U11847 ( n10962,instaddrpointer_reg_2_,n8998 );
   not U11848 ( n8998,n10973 );
   or U11849 ( n11656,n11573,n11078 );
   nand U11850 ( n11078,n11619,n10877 );
   nand U11851 ( n11573,n11693,instaddrpointer_reg_26_ );
   nor U11852 ( n11693,n11510,n11528 );
   nand U11853 ( n11528,n11694,instaddrpointer_reg_24_ );
   nor U11854 ( n11694,n11463,n11481 );
   not U11855 ( n11481,n11494 );
   nor U11856 ( n11494,n11695,n11436 );
   nand U11857 ( n11436,n11696,instaddrpointer_reg_20_ );
   nor U11858 ( n11696,n11370,n11390 );
   nand U11859 ( n11390,n11697,instaddrpointer_reg_18_ );
   nor U11860 ( n11697,n11324,n11342 );
   nand U11861 ( n11342,n11698,instaddrpointer_reg_16_ );
   nor U11862 ( n11698,n11278,n11296 );
   nand U11863 ( n11296,n11699,instaddrpointer_reg_14_ );
   nor U11864 ( n11699,n11232,n11250 );
   nand U11865 ( n11250,n11700,instaddrpointer_reg_12_ );
   nor U11866 ( n11700,n11186,n11204 );
   nand U11867 ( n11204,n11701,instaddrpointer_reg_10_ );
   nor U11868 ( n11701,n11140,n11158 );
   nand U11869 ( n11158,n11702,instaddrpointer_reg_8_ );
   nor U11870 ( n11702,n11094,n11112 );
   nand U11871 ( n11112,n11703,instaddrpointer_reg_6_ );
   nor U11872 ( n11703,n11047,n11065 );
   nand U11873 ( n11065,n11704,instaddrpointer_reg_4_ );
   nor U11874 ( n11704,n11020,n10999 );
   not U11875 ( n11020,n10961 );
   nand U11876 ( n10961,n10977,n10973 );
   nand U11877 ( n10973,instaddrpointer_reg_1_,instaddrpointer_reg_0_ );
   not U11878 ( n11047,instaddrpointer_reg_5_ );
   not U11879 ( n11094,instaddrpointer_reg_7_ );
   not U11880 ( n11186,instaddrpointer_reg_11_ );
   nand U11881 ( n11649,instaddrpointer_reg_28_,instaddrpointer_reg_27_ );
   nor U11882 ( n11633,n8753,n11705 );
   nand U11883 ( n11707,n11618,n11708 );
   and U11884 ( n11618,n11709,n11710 );
   nor U11885 ( n11709,n8816,n10891 );
   nand U11886 ( n10891,n11711,n10880 );
   not U11887 ( n10880,n11663 );
   nor U11888 ( n11711,n10808,n10768 );
   nand U11889 ( n11706,n11619,n11712 );
   nor U11890 ( n11619,n8871,n8816 );
   not U11891 ( n10974,n10934 );
   nand U11892 ( n10934,n11713,n11714 );
   nor U11893 ( n11714,n11715,n11716 );
   nor U11894 ( n11716,n11717,n9015 );
   nor U11895 ( n11717,n11718,n10915 );
   nand U11896 ( n10915,n11719,n11670 );
   nand U11897 ( n11670,n8874,n11720 );
   nand U11898 ( n11720,n11721,n11722 );
   nor U11899 ( n11719,n11723,n11724 );
   nor U11900 ( n11724,n11627,n11725 );
   nor U11901 ( n11725,n10818,n11726 );
   nor U11902 ( n11723,n11727,n10798 );
   nor U11903 ( n11727,n11728,n11729 );
   nand U11904 ( n11729,n11730,n10788 );
   nand U11905 ( n11730,n9391,n10881 );
   and U11906 ( n11718,n9367,n11731 );
   nor U11907 ( n11715,n11732,n11733 );
   nand U11908 ( n11733,n9275,n11722 );
   nor U11909 ( n11713,n11734,n11735 );
   nand U11910 ( n11735,n11736,n11737 );
   nand U11911 ( n11737,n11738,n10798 );
   nor U11912 ( n11738,n11739,n11740 );
   nand U11913 ( n11740,n9287,n11741 );
   nand U11914 ( n11739,n11742,n8862 );
   nand U11915 ( n11742,n8867,n10808 );
   nand U11916 ( n11736,n11743,n11627 );
   nor U11917 ( n11743,n11744,n11745 );
   nor U11918 ( n11744,n11746,n11747 );
   nand U11919 ( n11747,n10818,n11748 );
   nor U11920 ( n11746,n10890,n11749 );
   nand U11921 ( n11749,n11750,n8862 );
   nand U11922 ( n11750,n10906,n8867 );
   nor U11923 ( n11752,n11753,n11754 );
   nor U11924 ( n11754,n10928,n8788 );
   xor U11925 ( n10928,n11756,instaddrpointer_reg_0_ );
   nor U11926 ( n11753,n11757,n11758 );
   nor U11927 ( n11757,n11759,n8806 );
   nor U11928 ( n11751,n11760,n11761 );
   nor U11929 ( n11761,n8889,n11762 );
   not U11930 ( n8889,reip_reg_0_ );
   nor U11931 ( n11760,n11763,n11764 );
   nor U11932 ( n11766,n11767,n11768 );
   nor U11933 ( n11768,n11764,n11769 );
   nor U11934 ( n11767,n10943,n8788 );
   xor U11935 ( n10943,n11770,n11771 );
   nand U11936 ( n11771,n11772,n11773 );
   not U11937 ( n11772,n11774 );
   nor U11938 ( n11770,n11756,n8965 );
   nor U11939 ( n11765,n11775,n11776 );
   nand U11940 ( n11776,n11777,n11778 );
   nand U11941 ( n11778,n11759,n11779 );
   nand U11942 ( n11777,n8806,phyaddrpointer_reg_1_ );
   nor U11943 ( n11775,n9192,n11762 );
   nor U11944 ( n11781,n11782,n11783 );
   nand U11945 ( n11783,n11784,n11785 );
   nand U11946 ( n11785,n11786,n10963 );
   xor U11947 ( n10963,n11787,n11788 );
   xor U11948 ( n11788,n11789,n10977 );
   nand U11949 ( n11784,n11790,n11791 );
   nor U11950 ( n11782,n8828,n11793 );
   nor U11951 ( n11780,n11794,n11795 );
   nor U11952 ( n11795,n8808,n11796 );
   nor U11953 ( n11794,n9187,n8737 );
   nor U11954 ( n11798,n11799,n11800 );
   nand U11955 ( n11800,n11801,n11802 );
   nand U11956 ( n11802,n11803,n11786 );
   nor U11957 ( n11803,n11804,n10987 );
   and U11958 ( n10987,n11805,n11806 );
   not U11959 ( n11804,n10989 );
   nand U11960 ( n10989,n11807,n11808 );
   xor U11961 ( n11808,n11809,n10999 );
   nor U11962 ( n11807,n11810,n11811 );
   nor U11963 ( n11811,n11789,n10977 );
   not U11964 ( n11810,n11812 );
   nand U11965 ( n11801,n11813,n8820 );
   and U11966 ( n11799,n11814,n11759 );
   nor U11967 ( n11797,n11815,n11816 );
   nor U11968 ( n11816,n8808,n11817 );
   nor U11969 ( n11815,n9182,n8738 );
   nor U11970 ( n11819,n11820,n11821 );
   nand U11971 ( n11821,n11822,n11823 );
   nand U11972 ( n11823,n11824,n11786 );
   nor U11973 ( n11824,n11825,n11009 );
   nor U11974 ( n11009,n11826,n11827 );
   and U11975 ( n11827,instaddrpointer_reg_4_,n11828 );
   not U11976 ( n11825,n11011 );
   nand U11977 ( n11011,n11829,n11830 );
   xor U11978 ( n11830,n11828,n11027 );
   not U11979 ( n11027,instaddrpointer_reg_4_ );
   nor U11980 ( n11829,n11805,n11831 );
   nor U11981 ( n11831,n11832,n10999 );
   not U11982 ( n11805,n11833 );
   nand U11983 ( n11822,n11834,n11790 );
   nor U11984 ( n11820,n8827,n11835 );
   nor U11985 ( n11818,n11836,n11837 );
   nor U11986 ( n11837,n8810,n11838 );
   nor U11987 ( n11836,n9177,n11762 );
   nor U11988 ( n11840,n11841,n11842 );
   nand U11989 ( n11842,n11843,n11844 );
   nand U11990 ( n11844,n11786,n11037 );
   xor U11991 ( n11037,n11845,n11846 );
   and U11992 ( n11845,n11847,n11848 );
   nand U11993 ( n11843,n11790,n11849 );
   nor U11994 ( n11841,n11850,n11792 );
   nor U11995 ( n11839,n11851,n11852 );
   nor U11996 ( n11852,n8810,n11853 );
   nor U11997 ( n11851,n9172,n8737 );
   nor U11998 ( n11855,n11856,n11857 );
   nand U11999 ( n11857,n11858,n11859 );
   nand U12000 ( n11859,n11786,n11056 );
   xor U12001 ( n11056,n11860,n11861 );
   and U12002 ( n11860,n11862,n11863 );
   nand U12003 ( n11858,n11864,n11790 );
   nor U12004 ( n11856,n11792,n11865 );
   nor U12005 ( n11854,n11866,n11867 );
   nor U12006 ( n11867,n8810,n11868 );
   nor U12007 ( n11866,n9167,n8738 );
   nor U12008 ( n11870,n11871,n11872 );
   nand U12009 ( n11872,n11873,n11874 );
   nand U12010 ( n11874,n11786,n11084 );
   xor U12011 ( n11084,n11875,n11876 );
   nand U12012 ( n11876,n11862,n11877 );
   nor U12013 ( n11875,n11878,n11879 );
   nand U12014 ( n11873,n11880,n11790 );
   and U12015 ( n11871,n11881,n11759 );
   nor U12016 ( n11869,n11882,n11883 );
   nor U12017 ( n11883,n8807,n11884 );
   nor U12018 ( n11882,n9162,n11762 );
   nor U12019 ( n11886,n11887,n11888 );
   nand U12020 ( n11888,n11889,n11890 );
   or U12021 ( n11890,n11755,n11103 );
   nand U12022 ( n11103,n11891,n11892 );
   nand U12023 ( n11892,n11893,n11894 );
   nor U12024 ( n11891,n11895,n11896 );
   nor U12025 ( n11896,instaddrpointer_reg_8_,n11897 );
   nor U12026 ( n11897,n11898,n11893 );
   not U12027 ( n11893,n11899 );
   nor U12028 ( n11898,n11900,n11901 );
   nor U12029 ( n11895,n11119,n11902 );
   nand U12030 ( n11902,n11903,n11901 );
   nand U12031 ( n11889,n11790,n11904 );
   nor U12032 ( n11887,n11792,n11905 );
   nor U12033 ( n11885,n11906,n11907 );
   nor U12034 ( n11907,n8810,n11908 );
   nor U12035 ( n11906,n9157,n8737 );
   nor U12036 ( n11910,n11911,n11912 );
   nand U12037 ( n11912,n11913,n11914 );
   nand U12038 ( n11914,n11786,n11130 );
   xor U12039 ( n11130,n11915,n11916 );
   and U12040 ( n11915,n11917,n11918 );
   nand U12041 ( n11913,n11919,n8820 );
   nor U12042 ( n11911,n11920,n8828 );
   nor U12043 ( n11909,n11921,n11922 );
   nor U12044 ( n11922,n8807,n11923 );
   nor U12045 ( n11921,n9152,n8738 );
   nor U12046 ( n11925,n11926,n11927 );
   nand U12047 ( n11927,n11928,n11929 );
   or U12048 ( n11929,n8788,n11149 );
   nand U12049 ( n11149,n11930,n11931 );
   nand U12050 ( n11931,n11932,n11933 );
   nand U12051 ( n11933,n11934,n11935 );
   nand U12052 ( n11930,n11936,n11935 );
   nand U12053 ( n11928,n11937,n11790 );
   nor U12054 ( n11926,n8827,n11938 );
   nor U12055 ( n11924,n11939,n11940 );
   nor U12056 ( n11940,n8809,n11941 );
   nor U12057 ( n11939,n9147,n11762 );
   nor U12058 ( n11943,n11944,n11945 );
   nand U12059 ( n11945,n11946,n11947 );
   nand U12060 ( n11947,n11786,n11176 );
   xor U12061 ( n11176,n11948,n11949 );
   nand U12062 ( n11949,n11935,n11950 );
   not U12063 ( n11950,n11936 );
   nor U12064 ( n11936,n11951,n11932 );
   nor U12065 ( n11948,n11952,n11953 );
   not U12066 ( n11952,n11954 );
   nand U12067 ( n11946,n11955,n8820 );
   and U12068 ( n11944,n11956,n11759 );
   nor U12069 ( n11942,n11957,n11958 );
   nor U12070 ( n11958,n8809,n11959 );
   nor U12071 ( n11957,n9142,n8737 );
   nor U12072 ( n11961,n11962,n11963 );
   nand U12073 ( n11963,n11964,n11965 );
   or U12074 ( n11965,n11755,n11195 );
   nand U12075 ( n11195,n11966,n11967 );
   nand U12076 ( n11967,n11968,n11969 );
   nand U12077 ( n11969,n11970,n11971 );
   not U12078 ( n11968,n11972 );
   nand U12079 ( n11966,n11973,n11970 );
   not U12080 ( n11973,n11974 );
   nand U12081 ( n11964,n11790,n11975 );
   nor U12082 ( n11962,n8828,n11976 );
   nor U12083 ( n11960,n11977,n11978 );
   nor U12084 ( n11978,n8807,n11979 );
   nor U12085 ( n11977,n9137,n8738 );
   nor U12086 ( n11981,n11982,n11983 );
   nand U12087 ( n11983,n11984,n11985 );
   or U12088 ( n11985,n11755,n11222 );
   xor U12089 ( n11222,n11986,n11987 );
   nand U12090 ( n11987,n11988,n11989 );
   nand U12091 ( n11984,n11790,n11990 );
   and U12092 ( n11982,n11991,n11759 );
   not U12093 ( n11759,n8828 );
   nor U12094 ( n11980,n11992,n11993 );
   nor U12095 ( n11993,n8810,n11994 );
   nor U12096 ( n11992,n9132,n8737 );
   nor U12097 ( n11996,n11997,n11998 );
   nand U12098 ( n11998,n11999,n12000 );
   or U12099 ( n12000,n11755,n11241 );
   xor U12100 ( n11241,n12001,n12002 );
   nand U12101 ( n12002,n12003,n12004 );
   nand U12102 ( n11999,n12005,n8820 );
   nor U12103 ( n11997,n8827,n12006 );
   nor U12104 ( n11995,n12007,n12008 );
   nor U12105 ( n12008,n8808,n12009 );
   nor U12106 ( n12007,n9127,n11762 );
   nor U12107 ( n12011,n12012,n12013 );
   nand U12108 ( n12013,n12014,n12015 );
   or U12109 ( n12015,n11755,n11268 );
   xor U12110 ( n11268,n12016,n12017 );
   nand U12111 ( n12017,n12018,n12019 );
   nand U12112 ( n12014,n12020,n8820 );
   nor U12113 ( n12012,n8827,n12021 );
   nor U12114 ( n12010,n12022,n12023 );
   nor U12115 ( n12023,n8808,n12024 );
   nor U12116 ( n12022,n9122,n8738 );
   nor U12117 ( n12026,n12027,n12028 );
   nand U12118 ( n12028,n12029,n12030 );
   or U12119 ( n12030,n8788,n11287 );
   xor U12120 ( n11287,n12031,n12032 );
   nand U12121 ( n12032,n12033,n12034 );
   nand U12122 ( n12029,n12035,n8820 );
   nor U12123 ( n12027,n8828,n12036 );
   nor U12124 ( n12025,n12037,n12038 );
   nor U12125 ( n12038,n8808,n12039 );
   nor U12126 ( n12037,n9117,n8737 );
   nor U12127 ( n12041,n12042,n12043 );
   nand U12128 ( n12043,n12044,n12045 );
   nand U12129 ( n12045,n11786,n11314 );
   xor U12130 ( n11314,n12046,n12047 );
   nand U12131 ( n12047,n12033,n12048 );
   nand U12132 ( n12048,n12034,n12031 );
   nor U12133 ( n12046,n12049,n12050 );
   nand U12134 ( n12044,n11790,n12051 );
   nor U12135 ( n12042,n8828,n12052 );
   nor U12136 ( n12040,n12053,n12054 );
   nor U12137 ( n12054,n8809,n12055 );
   nor U12138 ( n12053,n9112,n11762 );
   nor U12139 ( n12057,n12058,n12059 );
   nand U12140 ( n12059,n12060,n12061 );
   nand U12141 ( n12061,n11786,n11333 );
   xor U12142 ( n11333,n12062,n12063 );
   xor U12143 ( n12062,n12064,n11349 );
   nand U12144 ( n12060,n12065,n8820 );
   nor U12145 ( n12058,n8828,n12066 );
   nor U12146 ( n12056,n12067,n12068 );
   nor U12147 ( n12068,n8808,n12069 );
   nor U12148 ( n12067,n9107,n8738 );
   nor U12149 ( n12071,n12072,n12073 );
   nand U12150 ( n12073,n12074,n12075 );
   or U12151 ( n12075,n8788,n11360 );
   nand U12152 ( n11360,n12076,n12077 );
   nand U12153 ( n12077,n12078,n12079 );
   nand U12154 ( n12079,n12080,n12081 );
   not U12155 ( n12078,n12082 );
   nand U12156 ( n12076,n12083,n12081 );
   nand U12157 ( n12074,n11790,n12084 );
   nor U12158 ( n12072,n12085,n8827 );
   nor U12159 ( n12070,n12086,n12087 );
   nor U12160 ( n12087,n8807,n12088 );
   nor U12161 ( n12086,n9102,n8737 );
   nor U12162 ( n12090,n12091,n12092 );
   nand U12163 ( n12092,n12093,n12094 );
   nand U12164 ( n12094,n12095,n11786 );
   nor U12165 ( n12095,n12096,n11379 );
   and U12166 ( n11379,n12097,n12098 );
   not U12167 ( n12096,n11381 );
   nand U12168 ( n11381,n12099,n12100 );
   xor U12169 ( n12100,instaddrpointer_reg_20_,n12064 );
   nor U12170 ( n12099,n12101,n12083 );
   nand U12171 ( n12093,n11790,n12102 );
   nor U12172 ( n12091,n8827,n12103 );
   nor U12173 ( n12089,n12104,n12105 );
   nor U12174 ( n12105,n8809,n12106 );
   nor U12175 ( n12104,n9097,n11762 );
   nor U12176 ( n12108,n12109,n12110 );
   nand U12177 ( n12110,n12111,n12112 );
   nand U12178 ( n12112,n11786,n11408 );
   xor U12179 ( n11408,n12113,n12114 );
   nand U12180 ( n12114,n12115,n12098 );
   nand U12181 ( n12098,instaddrpointer_reg_20_,n12116 );
   nor U12182 ( n12113,n12117,n12118 );
   nand U12183 ( n12111,n12119,n8820 );
   nor U12184 ( n12109,n12120,n8828 );
   nor U12185 ( n12107,n12121,n12122 );
   nor U12186 ( n12122,n8809,n12123 );
   nor U12187 ( n12121,n9092,n8737 );
   nor U12188 ( n12125,n12126,n12127 );
   nand U12189 ( n12127,n12128,n12129 );
   nand U12190 ( n12129,n11786,n11427 );
   nand U12191 ( n11427,n12130,n12131 );
   nand U12192 ( n12131,n12132,n12133 );
   nor U12193 ( n12130,n12134,n12135 );
   nor U12194 ( n12135,instaddrpointer_reg_22_,n12136 );
   xor U12195 ( n12136,n12133,n12064 );
   nor U12196 ( n12134,n11443,n12137 );
   or U12197 ( n12137,n12133,n12116 );
   nand U12198 ( n12133,n12138,n12139 );
   or U12199 ( n12139,n12115,n12117 );
   nor U12200 ( n12117,instaddrpointer_reg_21_,n12116 );
   nand U12201 ( n12128,n12140,n8820 );
   nor U12202 ( n12126,n11792,n12141 );
   nor U12203 ( n12124,n12142,n12143 );
   nor U12204 ( n12143,n8808,n12144 );
   nor U12205 ( n12142,n9087,n8738 );
   nor U12206 ( n12146,n12147,n12148 );
   nand U12207 ( n12148,n12149,n12150 );
   nand U12208 ( n12150,n11786,n11453 );
   xor U12209 ( n11453,n12151,n12152 );
   nand U12210 ( n12152,n12138,n12153 );
   nand U12211 ( n12153,n12154,n12155 );
   or U12212 ( n12155,n12132,n12097 );
   nor U12213 ( n12151,n12156,n12157 );
   nand U12214 ( n12149,n11790,n12158 );
   nor U12215 ( n12147,n8827,n12159 );
   nor U12216 ( n12145,n12160,n12161 );
   nor U12217 ( n12161,n8807,n12162 );
   nor U12218 ( n12160,n9082,n11762 );
   nor U12219 ( n12164,n12165,n12166 );
   nand U12220 ( n12166,n12167,n12168 );
   nand U12221 ( n12168,n11786,n11472 );
   xor U12222 ( n11472,n12169,n12170 );
   or U12223 ( n12170,n12171,n12172 );
   and U12224 ( n12169,n12173,n12174 );
   nand U12225 ( n12167,n12175,n8820 );
   nor U12226 ( n12165,n11792,n12176 );
   nor U12227 ( n12163,n12177,n12178 );
   nor U12228 ( n12178,n8809,n12179 );
   nor U12229 ( n12177,n9077,n8737 );
   nor U12230 ( n12181,n12182,n12183 );
   nand U12231 ( n12183,n12184,n12185 );
   nand U12232 ( n12185,n11786,n11500 );
   nand U12233 ( n11500,n12186,n12187 );
   nand U12234 ( n12187,n12188,n12189 );
   not U12235 ( n12188,n12190 );
   nor U12236 ( n12186,n12191,n12192 );
   nor U12237 ( n12192,n11510,n12193 );
   xor U12238 ( n12193,n12189,n12116 );
   nor U12239 ( n12191,instaddrpointer_reg_25_,n12194 );
   or U12240 ( n12194,n12189,n8823 );
   nand U12241 ( n12189,n12195,n12174 );
   not U12242 ( n12174,n12196 );
   nor U12243 ( n12195,n12171,n12197 );
   nor U12244 ( n12197,n12172,n12173 );
   nand U12245 ( n12173,n12198,n12097 );
   not U12246 ( n12097,n12115 );
   nand U12247 ( n12115,n12199,n12200 );
   nand U12248 ( n12200,n12201,n12081 );
   nand U12249 ( n12199,n8823,n11397 );
   nor U12250 ( n12198,n12202,n12157 );
   not U12251 ( n12202,n12154 );
   nand U12252 ( n12154,n8823,n11695 );
   nand U12253 ( n12184,n11790,n12203 );
   nor U12254 ( n12182,n8828,n12204 );
   nor U12255 ( n12180,n12205,n12206 );
   nor U12256 ( n12206,n8809,n12207 );
   nor U12257 ( n12205,n9072,n8738 );
   nor U12258 ( n12209,n12210,n12211 );
   nand U12259 ( n12211,n12212,n12213 );
   or U12260 ( n12213,n11755,n11519 );
   nand U12261 ( n11519,n12214,n12215 );
   nand U12262 ( n12215,n12216,n12217 );
   nand U12263 ( n12217,n12218,n12219 );
   not U12264 ( n12216,n12220 );
   nand U12265 ( n12214,n12221,n12218 );
   nand U12266 ( n12212,n11790,n12222 );
   nor U12267 ( n12210,n11792,n12223 );
   nor U12268 ( n12208,n12224,n12225 );
   nor U12269 ( n12225,n8809,n12226 );
   nor U12270 ( n12224,n9067,n11762 );
   nor U12271 ( n12228,n12229,n12230 );
   nand U12272 ( n12230,n12231,n12232 );
   nand U12273 ( n12232,n11786,n11546 );
   xor U12274 ( n11546,n12233,n12234 );
   nand U12275 ( n12234,n12235,n12236 );
   nor U12276 ( n12233,n12237,n12221 );
   not U12277 ( n12237,n12218 );
   nand U12278 ( n12231,n12238,n8820 );
   nor U12279 ( n12229,n11792,n12239 );
   nor U12280 ( n12227,n12240,n12241 );
   nor U12281 ( n12241,n8807,n12242 );
   nor U12282 ( n12240,n9062,n8737 );
   nor U12283 ( n12244,n12245,n12246 );
   nand U12284 ( n12246,n12247,n12248 );
   or U12285 ( n12248,n8788,n11564 );
   nand U12286 ( n11564,n12249,n12250 );
   nand U12287 ( n12250,n12251,n12252 );
   nand U12288 ( n12252,n12253,n12254 );
   nand U12289 ( n12254,n12255,n12218 );
   nor U12290 ( n12251,n12256,n12257 );
   nand U12291 ( n12249,n12258,n12259 );
   nand U12292 ( n12258,n12260,n12235 );
   nand U12293 ( n12247,n11790,n12261 );
   nor U12294 ( n12245,n11792,n12262 );
   nor U12295 ( n12243,n12263,n12264 );
   nor U12296 ( n12264,n8807,n12265 );
   nor U12297 ( n12263,n9057,n8738 );
   nor U12298 ( n12267,n12268,n12269 );
   nand U12299 ( n12269,n12270,n12271 );
   nand U12300 ( n12271,n11786,n11589 );
   xor U12301 ( n11589,n12272,n12273 );
   nand U12302 ( n12273,n12274,n12260 );
   and U12303 ( n12260,n12218,n12275 );
   nand U12304 ( n12275,n12256,n12253 );
   nor U12305 ( n12274,n12257,n12255 );
   not U12306 ( n12257,n12235 );
   nor U12307 ( n12272,n12276,n12277 );
   not U12308 ( n11786,n8788 );
   nand U12309 ( n12270,n11790,n12278 );
   nor U12310 ( n12268,n12279,n11792 );
   nor U12311 ( n12266,n12280,n12281 );
   nor U12312 ( n12281,n8810,n12282 );
   nor U12313 ( n12280,n9052,n11762 );
   nor U12314 ( n12284,n12285,n12286 );
   nand U12315 ( n12286,n12287,n12288 );
   or U12316 ( n12288,n11755,n11602 );
   nand U12317 ( n11602,n12289,n12290 );
   nand U12318 ( n12290,n12291,n8823 );
   nor U12319 ( n12289,n12292,n12293 );
   nor U12320 ( n12293,n11608,n12294 );
   xor U12321 ( n12294,n12295,n12064 );
   not U12322 ( n11608,instaddrpointer_reg_30_ );
   nor U12323 ( n12292,instaddrpointer_reg_30_,n12296 );
   nand U12324 ( n12296,n12116,n12295 );
   nand U12325 ( n12287,n11790,n12297 );
   nor U12326 ( n12285,n8827,n12298 );
   nor U12327 ( n12283,n12299,n12300 );
   nor U12328 ( n12300,n8810,n12301 );
   nor U12329 ( n12299,n9047,n8737 );
   nor U12330 ( n12303,n12304,n12305 );
   nand U12331 ( n12305,n12306,n12307 );
   nand U12332 ( n12307,n12308,n8820 );
   not U12333 ( n11790,n11764 );
   nand U12334 ( n11764,n12309,statebs16_reg );
   nor U12335 ( n12309,n8806,n8948 );
   or U12336 ( n12306,n11755,n11615 );
   xor U12337 ( n11615,n12310,n12311 );
   nand U12338 ( n12311,n12312,n12313 );
   nand U12339 ( n12313,n12314,n8823 );
   nand U12340 ( n12314,n12315,instaddrpointer_reg_30_ );
   not U12341 ( n12312,n12291 );
   nor U12342 ( n12291,n12295,instaddrpointer_reg_30_ );
   nand U12343 ( n12295,n12316,n12317 );
   nor U12344 ( n12317,n12255,n12318 );
   nand U12345 ( n12318,n12218,n12235 );
   nand U12346 ( n12235,instaddrpointer_reg_27_,n12116 );
   nand U12347 ( n12218,instaddrpointer_reg_26_,n12116 );
   not U12348 ( n12255,n12259 );
   nand U12349 ( n12259,instaddrpointer_reg_28_,n12116 );
   nor U12350 ( n12316,n12276,n12315 );
   and U12351 ( n12315,n12319,n12256 );
   and U12352 ( n12256,n12221,n12236 );
   nand U12353 ( n12236,n11556,n8823 );
   not U12354 ( n11556,instaddrpointer_reg_27_ );
   and U12355 ( n12221,n12220,n12219 );
   nand U12356 ( n12219,n8823,n11535 );
   not U12357 ( n11535,instaddrpointer_reg_26_ );
   nand U12358 ( n12220,n12320,n12321 );
   nor U12359 ( n12321,n12322,n12323 );
   or U12360 ( n12323,n12171,n12101 );
   not U12361 ( n12101,n12081 );
   nand U12362 ( n12081,instaddrpointer_reg_19_,n12116 );
   nor U12363 ( n12171,n11488,n8823 );
   not U12364 ( n11488,instaddrpointer_reg_24_ );
   nor U12365 ( n12322,n12324,n12325 );
   nand U12366 ( n12325,n12083,n12326 );
   nand U12367 ( n12326,n8823,n12327 );
   nand U12368 ( n12327,n11683,instaddrpointer_reg_20_ );
   not U12369 ( n11683,n11695 );
   nand U12370 ( n11695,instaddrpointer_reg_22_,instaddrpointer_reg_21_ );
   not U12371 ( n12083,n12201 );
   nand U12372 ( n12201,n12082,n12080 );
   nand U12373 ( n12080,n8823,n11370 );
   not U12374 ( n11370,instaddrpointer_reg_19_ );
   nand U12375 ( n12082,n12328,n12329 );
   nand U12376 ( n12329,n12063,n12330 );
   nand U12377 ( n12330,n11349,n8823 );
   not U12378 ( n11349,instaddrpointer_reg_18_ );
   nand U12379 ( n12063,n12331,n12332 );
   nand U12380 ( n12332,n12333,n12034 );
   nand U12381 ( n12034,n12334,n12335 );
   nor U12382 ( n12334,instaddrpointer_reg_16_,n12116 );
   nor U12383 ( n12333,n12050,n12336 );
   not U12384 ( n12336,n12031 );
   nand U12385 ( n12031,n12019,n12337 );
   nand U12386 ( n12337,n12018,n12016 );
   nand U12387 ( n12016,n12004,n12338 );
   nand U12388 ( n12338,n12003,n12001 );
   nand U12389 ( n12001,n12339,n11988 );
   nand U12390 ( n11988,n12340,instaddrpointer_reg_13_ );
   and U12391 ( n12340,n12341,n12342 );
   nand U12392 ( n12339,n11989,n11986 );
   nand U12393 ( n11986,n11974,n11970 );
   or U12394 ( n11970,n11211,n12343 );
   nand U12395 ( n11974,n11972,n11971 );
   nand U12396 ( n11971,n12343,n11211 );
   not U12397 ( n11211,instaddrpointer_reg_12_ );
   nand U12398 ( n12343,n12344,n12341 );
   nand U12399 ( n11972,n11954,n12345 );
   nand U12400 ( n12345,n12346,n12347 );
   nand U12401 ( n12347,n11932,n11935 );
   nand U12402 ( n11935,n12348,instaddrpointer_reg_10_ );
   and U12403 ( n12348,n12341,n12349 );
   and U12404 ( n11932,n11918,n12350 );
   nand U12405 ( n12350,n11917,n11916 );
   nand U12406 ( n11916,n11899,n12351 );
   nand U12407 ( n12351,instaddrpointer_reg_8_,n11901 );
   nand U12408 ( n11899,n11900,n12352 );
   nand U12409 ( n12352,n11894,n11119 );
   not U12410 ( n11119,instaddrpointer_reg_8_ );
   not U12411 ( n11894,n11901 );
   nand U12412 ( n11901,n12353,n12354 );
   nand U12413 ( n12354,n12355,n12356 );
   nor U12414 ( n12356,n12357,n12358 );
   nor U12415 ( n12355,n12359,n12360 );
   nand U12416 ( n12353,n12341,n12361 );
   not U12417 ( n11900,n11903 );
   nor U12418 ( n11903,n11878,n12362 );
   nor U12419 ( n12362,n12363,n11879 );
   nor U12420 ( n11879,n12364,instaddrpointer_reg_7_ );
   and U12421 ( n12363,n11862,n11877 );
   nand U12422 ( n11877,n11861,n11863 );
   or U12423 ( n11863,n12365,instaddrpointer_reg_6_ );
   nand U12424 ( n11861,n11848,n12366 );
   nand U12425 ( n12366,n11847,n11846 );
   nand U12426 ( n11846,n12367,n11826 );
   nand U12427 ( n11826,n12368,n12369 );
   nand U12428 ( n12369,n11806,n11833 );
   nand U12429 ( n11833,n12370,n12371 );
   nand U12430 ( n12371,n12372,n11812 );
   nand U12431 ( n11812,n11787,n12373 );
   nand U12432 ( n12373,n11789,n10977 );
   not U12433 ( n10977,instaddrpointer_reg_2_ );
   not U12434 ( n11789,n12374 );
   nand U12435 ( n11787,n11773,n12375 );
   nand U12436 ( n12375,n12376,instaddrpointer_reg_0_ );
   nor U12437 ( n12376,n11756,n11774 );
   nor U12438 ( n11774,n12377,instaddrpointer_reg_1_ );
   and U12439 ( n11756,n12378,n12379 );
   nor U12440 ( n12378,n12380,n12381 );
   nor U12441 ( n12381,n12359,n12382 );
   nor U12442 ( n12380,n10642,n12383 );
   nand U12443 ( n11773,instaddrpointer_reg_1_,n12377 );
   nand U12444 ( n12377,n12384,n12385 );
   nor U12445 ( n12385,n12386,n12387 );
   nor U12446 ( n12387,n12388,n12359 );
   xor U12447 ( n12388,n12382,n12389 );
   nor U12448 ( n12384,n12390,n9392 );
   nor U12449 ( n12390,n12383,n10834 );
   not U12450 ( n10834,n8917 );
   nand U12451 ( n12372,instaddrpointer_reg_2_,n12374 );
   nand U12452 ( n12374,n12391,n12379 );
   nand U12453 ( n12379,n9391,n10788 );
   nor U12454 ( n12391,n12392,n12393 );
   nor U12455 ( n12393,n9782,n12383 );
   nor U12456 ( n12392,n12394,n12359 );
   nor U12457 ( n12394,n12395,n12396 );
   nor U12458 ( n12395,n12397,n12398 );
   nand U12459 ( n12370,n11832,n10999 );
   not U12460 ( n10999,instaddrpointer_reg_3_ );
   not U12461 ( n11832,n11809 );
   nand U12462 ( n11806,instaddrpointer_reg_3_,n11809 );
   nand U12463 ( n11809,n12399,n12400 );
   nand U12464 ( n12400,n8874,n12401 );
   xor U12465 ( n12401,n12402,n12403 );
   nand U12466 ( n12399,n8944,n12341 );
   or U12467 ( n12368,n11828,instaddrpointer_reg_4_ );
   nand U12468 ( n12367,instaddrpointer_reg_4_,n11828 );
   nand U12469 ( n11828,n12404,n12405 );
   or U12470 ( n12405,n12406,n12359 );
   xor U12471 ( n12406,n12407,n12408 );
   nand U12472 ( n12408,n12403,n12402 );
   nand U12473 ( n12404,n12409,n12341 );
   or U12474 ( n11847,n12410,instaddrpointer_reg_5_ );
   nand U12475 ( n11848,instaddrpointer_reg_5_,n12410 );
   nand U12476 ( n12410,n12411,n12412 );
   nand U12477 ( n12412,n12413,n8874 );
   nor U12478 ( n12413,n12414,n12415 );
   nor U12479 ( n12415,n12416,n12417 );
   not U12480 ( n12414,n12360 );
   nand U12481 ( n12411,n12418,n12341 );
   nand U12482 ( n11862,instaddrpointer_reg_6_,n12365 );
   nand U12483 ( n12365,n12419,n12420 );
   nand U12484 ( n12420,n12421,n8874 );
   xor U12485 ( n12421,n12358,n12360 );
   or U12486 ( n12419,n12422,n12383 );
   and U12487 ( n11878,instaddrpointer_reg_7_,n12364 );
   nand U12488 ( n12364,n12423,n12424 );
   nand U12489 ( n12424,n12425,n12426 );
   nor U12490 ( n12425,n12427,n12383 );
   nand U12491 ( n12423,n12428,n8874 );
   xor U12492 ( n12428,n12429,n12430 );
   nor U12493 ( n12429,n12358,n12360 );
   nand U12494 ( n12360,n12416,n12417 );
   and U12495 ( n12416,n12431,n12407 );
   nor U12496 ( n12431,n12432,n12396 );
   not U12497 ( n12396,n12402 );
   nand U12498 ( n12402,n12397,n12398 );
   nand U12499 ( n12398,n12433,n12382 );
   not U12500 ( n12358,n12434 );
   nand U12501 ( n11917,n11140,n12435 );
   nand U12502 ( n12435,n12436,n12341 );
   not U12503 ( n11140,instaddrpointer_reg_9_ );
   nand U12504 ( n11918,n12437,instaddrpointer_reg_9_ );
   nor U12505 ( n12437,n12383,n12438 );
   nor U12506 ( n12346,n11951,n11953 );
   nor U12507 ( n11953,instaddrpointer_reg_11_,n12439 );
   not U12508 ( n11951,n11934 );
   nand U12509 ( n11934,n11165,n12440 );
   nand U12510 ( n12440,n12349,n12341 );
   not U12511 ( n11165,instaddrpointer_reg_10_ );
   nand U12512 ( n11954,instaddrpointer_reg_11_,n12439 );
   and U12513 ( n12439,n12441,n12341 );
   nand U12514 ( n11989,n11232,n12442 );
   nand U12515 ( n12442,n12342,n12341 );
   not U12516 ( n11232,instaddrpointer_reg_13_ );
   nand U12517 ( n12003,n11257,n12443 );
   nand U12518 ( n12443,n12444,n12341 );
   not U12519 ( n11257,instaddrpointer_reg_14_ );
   nand U12520 ( n12004,n12445,instaddrpointer_reg_14_ );
   nor U12521 ( n12445,n12383,n12446 );
   nand U12522 ( n12018,n11278,n12447 );
   nand U12523 ( n12447,n12448,n12341 );
   not U12524 ( n11278,instaddrpointer_reg_15_ );
   nand U12525 ( n12019,n12449,instaddrpointer_reg_15_ );
   and U12526 ( n12449,n12341,n12448 );
   nor U12527 ( n12331,n12049,n12450 );
   nor U12528 ( n12450,n12033,n12050 );
   nor U12529 ( n12050,n12116,instaddrpointer_reg_17_ );
   nand U12530 ( n12033,instaddrpointer_reg_16_,n12451 );
   nand U12531 ( n12451,n12335,n8823 );
   nand U12532 ( n12335,n12452,n12453 );
   nor U12533 ( n12452,n12454,n12383 );
   nor U12534 ( n12049,n11324,n8823 );
   not U12535 ( n11324,instaddrpointer_reg_17_ );
   nand U12536 ( n12328,instaddrpointer_reg_18_,n12116 );
   nand U12537 ( n12324,n12455,n12190 );
   nand U12538 ( n12190,n11510,n8823 );
   nor U12539 ( n12455,n12172,n12157 );
   nor U12540 ( n12157,instaddrpointer_reg_23_,n12116 );
   nor U12541 ( n12172,n12116,instaddrpointer_reg_24_ );
   nor U12542 ( n12320,n12456,n12196 );
   nand U12543 ( n12196,n12457,n12138 );
   nor U12544 ( n12138,n12458,n12118 );
   nor U12545 ( n12118,n11418,n12064 );
   not U12546 ( n11418,instaddrpointer_reg_21_ );
   nor U12547 ( n12458,n11397,n12064 );
   not U12548 ( n11397,instaddrpointer_reg_20_ );
   nor U12549 ( n12457,n12132,n12156 );
   nor U12550 ( n12156,n11463,n8823 );
   not U12551 ( n11463,instaddrpointer_reg_23_ );
   nor U12552 ( n12132,n11443,n8823 );
   not U12553 ( n11443,instaddrpointer_reg_22_ );
   nor U12554 ( n12456,n12064,n11510 );
   not U12555 ( n11510,instaddrpointer_reg_25_ );
   nor U12556 ( n12319,n12277,n12459 );
   not U12557 ( n12459,n12253 );
   nand U12558 ( n12253,n11580,n8823 );
   not U12559 ( n11580,instaddrpointer_reg_28_ );
   nor U12560 ( n12277,n12116,instaddrpointer_reg_29_ );
   not U12561 ( n12116,n12064 );
   nor U12562 ( n12276,n11596,n8823 );
   not U12563 ( n11596,instaddrpointer_reg_29_ );
   xor U12564 ( n12310,n12064,n8997 );
   nand U12565 ( n12064,n12460,n12454 );
   nor U12566 ( n12460,n12453,n12383 );
   nand U12567 ( n11755,state2_reg_0_,n8810 );
   nor U12568 ( n12304,n12461,n8827 );
   nand U12569 ( n11792,n12462,n12463 );
   nor U12570 ( n12463,n7819,n8868 );
   nor U12571 ( n12462,state2_reg_0_,n8806 );
   nor U12572 ( n12302,n12464,n12465 );
   nor U12573 ( n12465,n8808,n12466 );
   nor U12574 ( n12464,n9045,n8738 );
   nand U12575 ( n11762,n8868,n8808 );
   nand U12576 ( n12468,n8857,n8821 );
   and U12577 ( n12467,n12469,n12470 );
   nand U12578 ( n12472,n8799,eax_reg_15_ );
   nor U12579 ( n12471,n12474,n12475 );
   nor U12580 ( n12475,n12476,n12477 );
   nor U12581 ( n12474,n8834,n12478 );
   nand U12582 ( n12480,n12473,eax_reg_14_ );
   nor U12583 ( n12479,n12481,n12482 );
   nor U12584 ( n12481,n8834,n12483 );
   nand U12585 ( n12485,n12473,eax_reg_13_ );
   nor U12586 ( n12484,n12486,n12487 );
   nor U12587 ( n12486,n8836,n12488 );
   nand U12588 ( n12490,n12473,eax_reg_12_ );
   nor U12589 ( n12489,n12491,n12492 );
   nor U12590 ( n12491,n8836,n12493 );
   nand U12591 ( n12495,n12473,eax_reg_11_ );
   nor U12592 ( n12494,n12496,n12497 );
   nor U12593 ( n12496,n8833,n12498 );
   nand U12594 ( n12500,n12473,eax_reg_10_ );
   nor U12595 ( n12499,n12501,n12502 );
   nor U12596 ( n12501,n8833,n12503 );
   nand U12597 ( n12505,n12473,eax_reg_9_ );
   nor U12598 ( n12504,n12506,n12507 );
   nor U12599 ( n12506,n8835,n12508 );
   nand U12600 ( n12510,n12473,eax_reg_8_ );
   nor U12601 ( n12509,n12511,n12512 );
   nor U12602 ( n12511,n8833,n12513 );
   nand U12603 ( n12515,n12473,eax_reg_7_ );
   nor U12604 ( n12514,n12516,n12517 );
   nor U12605 ( n12516,n8835,n12518 );
   nand U12606 ( n12520,n12473,eax_reg_6_ );
   nor U12607 ( n12519,n12521,n12522 );
   nor U12608 ( n12521,n8835,n12523 );
   nand U12609 ( n12525,n12473,eax_reg_5_ );
   nor U12610 ( n12524,n12526,n12527 );
   nor U12611 ( n12526,n8833,n12528 );
   nand U12612 ( n12530,n12473,eax_reg_4_ );
   nor U12613 ( n12529,n12531,n12532 );
   nor U12614 ( n12531,n8834,n12533 );
   nand U12615 ( n12535,n12473,eax_reg_3_ );
   nor U12616 ( n12534,n12536,n12537 );
   nor U12617 ( n12536,n8833,n12538 );
   nand U12618 ( n12540,n12473,eax_reg_2_ );
   nor U12619 ( n12539,n12541,n12542 );
   nor U12620 ( n12541,n8835,n12543 );
   nand U12621 ( n12545,n12473,eax_reg_1_ );
   nor U12622 ( n12544,n12546,n12547 );
   nor U12623 ( n12546,n8835,n12548 );
   nand U12624 ( n12550,n12473,eax_reg_0_ );
   nor U12625 ( n12549,n12551,n12552 );
   nor U12626 ( n12551,n8835,n12553 );
   nand U12627 ( n12555,n12473,eax_reg_30_ );
   nor U12628 ( n12554,n12556,n12482 );
   nor U12629 ( n12482,n12476,n12557 );
   nor U12630 ( n12556,n8834,n12558 );
   nand U12631 ( n12560,n8799,eax_reg_29_ );
   nor U12632 ( n12559,n12561,n12487 );
   nor U12633 ( n12487,n12476,n12562 );
   nor U12634 ( n12561,n8836,n12563 );
   nand U12635 ( n12565,n8799,eax_reg_28_ );
   nor U12636 ( n12564,n12566,n12492 );
   nor U12637 ( n12492,n12476,n12567 );
   nor U12638 ( n12566,n8836,n12568 );
   nand U12639 ( n12570,n8799,eax_reg_27_ );
   nor U12640 ( n12569,n12571,n12497 );
   nor U12641 ( n12497,n12476,n12572 );
   nor U12642 ( n12571,n8834,n12573 );
   nand U12643 ( n12575,n8799,eax_reg_26_ );
   nor U12644 ( n12574,n12576,n12502 );
   nor U12645 ( n12502,n12476,n12577 );
   nor U12646 ( n12576,n8834,n12578 );
   nand U12647 ( n12580,n8799,eax_reg_25_ );
   nor U12648 ( n12579,n12581,n12507 );
   nor U12649 ( n12507,n12476,n12582 );
   nor U12650 ( n12581,n8833,n12583 );
   nand U12651 ( n12585,n8799,eax_reg_24_ );
   nor U12652 ( n12584,n12586,n12512 );
   nor U12653 ( n12512,n12476,n12587 );
   nor U12654 ( n12586,n8835,n12588 );
   nand U12655 ( n12590,n8799,eax_reg_23_ );
   nor U12656 ( n12589,n12591,n12517 );
   nor U12657 ( n12517,n12592,n8785 );
   nor U12658 ( n12591,n8835,n12593 );
   nand U12659 ( n12595,n8799,eax_reg_22_ );
   nor U12660 ( n12594,n12596,n12522 );
   nor U12661 ( n12522,n12597,n8785 );
   nor U12662 ( n12596,n8834,n12598 );
   nand U12663 ( n12600,n8799,eax_reg_21_ );
   nor U12664 ( n12599,n12601,n12527 );
   nor U12665 ( n12527,n12602,n8785 );
   nor U12666 ( n12601,n8834,n12603 );
   nand U12667 ( n12605,n8799,eax_reg_20_ );
   nor U12668 ( n12604,n12606,n12532 );
   nor U12669 ( n12532,n12607,n12476 );
   nor U12670 ( n12606,n8836,n12608 );
   nand U12671 ( n12610,n8799,eax_reg_19_ );
   nor U12672 ( n12609,n12611,n12537 );
   nor U12673 ( n12537,n12612,n12476 );
   nor U12674 ( n12611,n8836,n12613 );
   nand U12675 ( n12615,n8799,eax_reg_18_ );
   nor U12676 ( n12614,n12616,n12542 );
   nor U12677 ( n12542,n12617,n8785 );
   nor U12678 ( n12616,n8833,n12618 );
   nand U12679 ( n12620,n8799,eax_reg_17_ );
   nor U12680 ( n12619,n12621,n12547 );
   nor U12681 ( n12547,n12622,n8785 );
   nor U12682 ( n12621,n8833,n12623 );
   nand U12683 ( n12625,n8799,eax_reg_16_ );
   and U12684 ( n12473,n8836,n10906 );
   nor U12685 ( n12624,n12626,n12552 );
   nor U12686 ( n12552,n12627,n8785 );
   nand U12687 ( n12476,n8834,n10808 );
   nor U12688 ( n12626,n8836,n12628 );
   nor U12689 ( n12630,n9391,n12631 );
   nor U12690 ( n12631,n8874,n8862 );
   nor U12691 ( n12629,n10890,n11745 );
   nand U12692 ( n12633,datao_reg_0_,n8795 );
   nor U12693 ( n12632,n12635,n12636 );
   nor U12694 ( n12636,n12637,n12638 );
   nor U12695 ( n12635,n12553,n8735 );
   not U12696 ( n12553,lword_reg_0_ );
   nand U12697 ( n12641,datao_reg_1_,n8795 );
   nor U12698 ( n12640,n12642,n12643 );
   and U12699 ( n12643,eax_reg_1_,n12644 );
   nor U12700 ( n12642,n12548,n8735 );
   not U12701 ( n12548,lword_reg_1_ );
   nand U12702 ( n12646,datao_reg_2_,n12634 );
   nor U12703 ( n12645,n12647,n12648 );
   nor U12704 ( n12648,n12649,n12638 );
   nor U12705 ( n12647,n12543,n8736 );
   not U12706 ( n12543,lword_reg_2_ );
   nand U12707 ( n12651,datao_reg_3_,n12634 );
   nor U12708 ( n12650,n12652,n12653 );
   nor U12709 ( n12653,n12654,n12638 );
   nor U12710 ( n12652,n12538,n12639 );
   not U12711 ( n12538,lword_reg_3_ );
   nand U12712 ( n12656,datao_reg_4_,n12634 );
   nor U12713 ( n12655,n12657,n12658 );
   nor U12714 ( n12658,n12659,n12638 );
   nor U12715 ( n12657,n12533,n8735 );
   not U12716 ( n12533,lword_reg_4_ );
   nand U12717 ( n12661,datao_reg_5_,n12634 );
   nor U12718 ( n12660,n12662,n12663 );
   nor U12719 ( n12663,n12664,n12638 );
   nor U12720 ( n12662,n12528,n8736 );
   not U12721 ( n12528,lword_reg_5_ );
   nand U12722 ( n12666,datao_reg_6_,n12634 );
   nor U12723 ( n12665,n12667,n12668 );
   nor U12724 ( n12668,n12669,n12638 );
   nor U12725 ( n12667,n12523,n12639 );
   not U12726 ( n12523,lword_reg_6_ );
   nand U12727 ( n12671,datao_reg_7_,n12634 );
   nor U12728 ( n12670,n12672,n12673 );
   nor U12729 ( n12673,n12674,n12638 );
   nor U12730 ( n12672,n12518,n8735 );
   not U12731 ( n12518,lword_reg_7_ );
   nand U12732 ( n12676,datao_reg_8_,n12634 );
   nor U12733 ( n12675,n12677,n12678 );
   and U12734 ( n12678,eax_reg_8_,n12644 );
   nor U12735 ( n12677,n12513,n8736 );
   not U12736 ( n12513,lword_reg_8_ );
   nand U12737 ( n12680,datao_reg_9_,n12634 );
   nor U12738 ( n12679,n12681,n12682 );
   nor U12739 ( n12682,n12683,n12638 );
   nor U12740 ( n12681,n12508,n12639 );
   not U12741 ( n12508,lword_reg_9_ );
   nand U12742 ( n12685,datao_reg_10_,n12634 );
   nor U12743 ( n12684,n12686,n12687 );
   and U12744 ( n12687,eax_reg_10_,n12644 );
   nor U12745 ( n12686,n12503,n8735 );
   not U12746 ( n12503,lword_reg_10_ );
   nand U12747 ( n12689,datao_reg_11_,n12634 );
   nor U12748 ( n12688,n12690,n12691 );
   nor U12749 ( n12691,n12692,n12638 );
   nor U12750 ( n12690,n12498,n8736 );
   not U12751 ( n12498,lword_reg_11_ );
   nand U12752 ( n12694,datao_reg_12_,n12634 );
   nor U12753 ( n12693,n12695,n12696 );
   nor U12754 ( n12696,n12697,n12638 );
   nor U12755 ( n12695,n12493,n12639 );
   not U12756 ( n12493,lword_reg_12_ );
   nand U12757 ( n12699,datao_reg_13_,n12634 );
   nor U12758 ( n12698,n12700,n12701 );
   nor U12759 ( n12701,n12702,n12638 );
   nor U12760 ( n12700,n12488,n8735 );
   not U12761 ( n12488,lword_reg_13_ );
   nand U12762 ( n12704,datao_reg_14_,n12634 );
   nor U12763 ( n12703,n12705,n12706 );
   and U12764 ( n12706,eax_reg_14_,n12644 );
   nor U12765 ( n12705,n12483,n12639 );
   not U12766 ( n12483,lword_reg_14_ );
   nand U12767 ( n12708,datao_reg_15_,n12634 );
   nor U12768 ( n12707,n12709,n12710 );
   and U12769 ( n12710,eax_reg_15_,n12644 );
   nor U12770 ( n12709,n12478,n8736 );
   not U12771 ( n12478,lword_reg_15_ );
   nand U12772 ( n12712,datao_reg_16_,n12634 );
   nor U12773 ( n12711,n12713,n12714 );
   nor U12774 ( n12714,n12715,n12716 );
   nor U12775 ( n12713,n12628,n8735 );
   not U12776 ( n12628,uword_reg_0_ );
   nand U12777 ( n12718,datao_reg_17_,n12634 );
   nor U12778 ( n12717,n12719,n12720 );
   nor U12779 ( n12720,n12721,n8791 );
   nor U12780 ( n12719,n12623,n12639 );
   not U12781 ( n12623,uword_reg_1_ );
   nand U12782 ( n12723,datao_reg_18_,n12634 );
   nor U12783 ( n12722,n12724,n12725 );
   nor U12784 ( n12725,n12726,n8791 );
   nor U12785 ( n12724,n12618,n8736 );
   not U12786 ( n12618,uword_reg_2_ );
   nand U12787 ( n12728,datao_reg_19_,n12634 );
   nor U12788 ( n12727,n12729,n12730 );
   nor U12789 ( n12730,n12731,n8791 );
   nor U12790 ( n12729,n12613,n12639 );
   not U12791 ( n12613,uword_reg_3_ );
   nand U12792 ( n12733,datao_reg_20_,n12634 );
   nor U12793 ( n12732,n12734,n12735 );
   nor U12794 ( n12735,n12736,n12716 );
   nor U12795 ( n12734,n12608,n8735 );
   not U12796 ( n12608,uword_reg_4_ );
   nand U12797 ( n12738,datao_reg_21_,n12634 );
   nor U12798 ( n12737,n12739,n12740 );
   nor U12799 ( n12740,n12741,n12716 );
   nor U12800 ( n12739,n12603,n8736 );
   not U12801 ( n12603,uword_reg_5_ );
   nand U12802 ( n12743,datao_reg_22_,n12634 );
   nor U12803 ( n12742,n12744,n12745 );
   nor U12804 ( n12745,n12746,n12716 );
   nor U12805 ( n12744,n12598,n12639 );
   not U12806 ( n12598,uword_reg_6_ );
   nand U12807 ( n12748,datao_reg_23_,n12634 );
   nor U12808 ( n12747,n12749,n12750 );
   nor U12809 ( n12750,n12751,n12716 );
   nor U12810 ( n12749,n12593,n8735 );
   not U12811 ( n12593,uword_reg_7_ );
   nand U12812 ( n12753,datao_reg_24_,n8795 );
   nor U12813 ( n12752,n12754,n12755 );
   nor U12814 ( n12755,n12756,n12716 );
   nor U12815 ( n12754,n12588,n8736 );
   not U12816 ( n12588,uword_reg_8_ );
   nand U12817 ( n12758,datao_reg_25_,n8795 );
   nor U12818 ( n12757,n12759,n12760 );
   nor U12819 ( n12760,n12761,n12716 );
   nor U12820 ( n12759,n12583,n12639 );
   not U12821 ( n12583,uword_reg_9_ );
   nand U12822 ( n12763,datao_reg_26_,n8795 );
   nor U12823 ( n12762,n12764,n12765 );
   nor U12824 ( n12765,n12766,n12716 );
   nor U12825 ( n12764,n12578,n8735 );
   not U12826 ( n12578,uword_reg_10_ );
   nand U12827 ( n12768,datao_reg_27_,n8795 );
   nor U12828 ( n12767,n12769,n12770 );
   nor U12829 ( n12770,n12771,n12716 );
   nor U12830 ( n12769,n12573,n8736 );
   not U12831 ( n12573,uword_reg_11_ );
   nand U12832 ( n12773,datao_reg_28_,n8795 );
   nor U12833 ( n12772,n12774,n12775 );
   nor U12834 ( n12775,n12776,n12716 );
   nor U12835 ( n12774,n12568,n12639 );
   not U12836 ( n12568,uword_reg_12_ );
   nand U12837 ( n12778,datao_reg_29_,n8795 );
   nor U12838 ( n12777,n12779,n12780 );
   nor U12839 ( n12780,n12781,n12716 );
   nor U12840 ( n12779,n12563,n8735 );
   not U12841 ( n12563,uword_reg_13_ );
   nand U12842 ( n12783,datao_reg_30_,n8795 );
   nor U12843 ( n12782,n12784,n12785 );
   nor U12844 ( n12785,n12786,n12716 );
   nand U12845 ( n12716,n12644,n10818 );
   not U12846 ( n12644,n12638 );
   nand U12847 ( n12638,state2_reg_0_,n12787 );
   nor U12848 ( n12784,n12558,n8736 );
   nand U12849 ( n12639,n8821,n12787 );
   not U12850 ( n12558,uword_reg_14_ );
   not U12851 ( n12634,n12787 );
   nand U12852 ( n12787,n12788,n12789 );
   nand U12853 ( n12789,n12790,n8876 );
   nor U12854 ( n12790,n12791,n11745 );
   nor U12855 ( n12791,n11712,n8961 );
   not U12856 ( n8961,n9350 );
   not U12857 ( n11712,n9311 );
   nand U12858 ( n9311,n8874,n10914 );
   nand U12859 ( n12788,n9020,n8821 );
   not U12860 ( n9020,n8860 );
   nand U12861 ( n8860,state2_reg_1_,state2_reg_2_ );
   nand U12862 ( n12793,n12794,eax_reg_0_ );
   nor U12863 ( n12792,n12795,n12796 );
   nor U12864 ( n12796,n11763,n8730 );
   nor U12865 ( n12795,n12627,n12797 );
   nand U12866 ( n12799,n8813,eax_reg_1_ );
   nor U12867 ( n12798,n12800,n12801 );
   nor U12868 ( n12801,n11769,n8728 );
   nor U12869 ( n12800,n12622,n8783 );
   nand U12870 ( n12803,n8813,eax_reg_2_ );
   nor U12871 ( n12802,n12804,n12805 );
   nor U12872 ( n12805,n12806,n8729 );
   nor U12873 ( n12804,n12617,n8783 );
   nand U12874 ( n12808,n12794,eax_reg_3_ );
   nor U12875 ( n12807,n12809,n12810 );
   nor U12876 ( n12810,n12811,n8730 );
   nor U12877 ( n12809,n12612,n8783 );
   nand U12878 ( n12813,n12794,eax_reg_4_ );
   nor U12879 ( n12812,n12814,n12815 );
   nor U12880 ( n12815,n12816,n8728 );
   nor U12881 ( n12814,n12607,n12797 );
   nand U12882 ( n12818,n12794,eax_reg_5_ );
   nor U12883 ( n12817,n12819,n12820 );
   nor U12884 ( n12820,n12821,n8729 );
   nor U12885 ( n12819,n12602,n12797 );
   nand U12886 ( n12823,n12794,eax_reg_6_ );
   nor U12887 ( n12822,n12824,n12825 );
   nor U12888 ( n12825,n12826,n8730 );
   nor U12889 ( n12824,n12597,n12797 );
   nand U12890 ( n12828,n12794,eax_reg_7_ );
   nor U12891 ( n12827,n12829,n12830 );
   nor U12892 ( n12830,n12831,n8728 );
   nor U12893 ( n12829,n12592,n12797 );
   nand U12894 ( n12833,n12794,eax_reg_8_ );
   nor U12895 ( n12832,n12834,n12835 );
   nor U12896 ( n12835,n12836,n8729 );
   nor U12897 ( n12834,n12587,n12797 );
   nand U12898 ( n12838,n12794,eax_reg_9_ );
   nor U12899 ( n12837,n12839,n12840 );
   nor U12900 ( n12840,n12841,n8730 );
   nor U12901 ( n12839,n12582,n12797 );
   nand U12902 ( n12843,n12794,eax_reg_10_ );
   nor U12903 ( n12842,n12844,n12845 );
   nor U12904 ( n12845,n12846,n8728 );
   nor U12905 ( n12844,n12577,n12797 );
   nand U12906 ( n12848,n8813,eax_reg_11_ );
   nor U12907 ( n12847,n12849,n12850 );
   nor U12908 ( n12850,n12851,n8729 );
   nor U12909 ( n12849,n12572,n12797 );
   nand U12910 ( n12853,n12794,eax_reg_12_ );
   nor U12911 ( n12852,n12854,n12855 );
   nor U12912 ( n12855,n12856,n8730 );
   nor U12913 ( n12854,n12567,n12797 );
   nand U12914 ( n12858,n8813,eax_reg_13_ );
   nor U12915 ( n12857,n12859,n12860 );
   nor U12916 ( n12860,n12861,n8728 );
   nor U12917 ( n12859,n12562,n12797 );
   nand U12918 ( n12863,n12794,eax_reg_14_ );
   nor U12919 ( n12862,n12864,n12865 );
   nor U12920 ( n12865,n12866,n8729 );
   nor U12921 ( n12864,n12557,n8783 );
   nand U12922 ( n12868,n12794,eax_reg_15_ );
   nor U12923 ( n12867,n12869,n12870 );
   nor U12924 ( n12870,n12871,n8730 );
   nor U12925 ( n12869,n12477,n12797 );
   nand U12926 ( n12797,n12872,n7821 );
   nor U12927 ( n12872,n12874,n11661 );
   not U12928 ( n12477,datai_15_ );
   nor U12929 ( n12876,n12877,n12878 );
   nor U12930 ( n12878,n12879,n8728 );
   nor U12931 ( n12877,n12627,n12880 );
   not U12932 ( n12627,datai_0_ );
   nor U12933 ( n12875,n12881,n12882 );
   nor U12934 ( n12882,n12715,n12873 );
   and U12935 ( n12881,datai_16_,n12883 );
   nor U12936 ( n12885,n12886,n12887 );
   nor U12937 ( n12887,n12888,n8729 );
   nor U12938 ( n12886,n12622,n8778 );
   not U12939 ( n12622,datai_1_ );
   nor U12940 ( n12884,n12889,n12890 );
   nor U12941 ( n12890,n12721,n12873 );
   and U12942 ( n12889,datai_17_,n12883 );
   nor U12943 ( n12892,n12893,n12894 );
   nor U12944 ( n12894,n12895,n8730 );
   nor U12945 ( n12893,n12617,n8778 );
   not U12946 ( n12617,datai_2_ );
   nor U12947 ( n12891,n12896,n12897 );
   nor U12948 ( n12897,n12726,n12873 );
   and U12949 ( n12896,datai_18_,n12883 );
   nor U12950 ( n12899,n12900,n12901 );
   nor U12951 ( n12901,n12902,n8728 );
   nor U12952 ( n12900,n12612,n8778 );
   not U12953 ( n12612,datai_3_ );
   nor U12954 ( n12898,n12903,n12904 );
   nor U12955 ( n12904,n12731,n12873 );
   and U12956 ( n12903,datai_19_,n12883 );
   nor U12957 ( n12906,n12907,n12908 );
   nor U12958 ( n12908,n12909,n8729 );
   nor U12959 ( n12907,n12607,n12880 );
   not U12960 ( n12607,datai_4_ );
   nor U12961 ( n12905,n12910,n12911 );
   nor U12962 ( n12911,n12736,n7821 );
   and U12963 ( n12910,datai_20_,n12883 );
   nor U12964 ( n12913,n12914,n12915 );
   nor U12965 ( n12915,n12916,n8730 );
   nor U12966 ( n12914,n12602,n12880 );
   not U12967 ( n12602,datai_5_ );
   nor U12968 ( n12912,n12917,n12918 );
   nor U12969 ( n12918,n12741,n7821 );
   and U12970 ( n12917,datai_21_,n12883 );
   nor U12971 ( n12920,n12921,n12922 );
   nor U12972 ( n12922,n12923,n8728 );
   nor U12973 ( n12921,n12597,n12880 );
   not U12974 ( n12597,datai_6_ );
   nor U12975 ( n12919,n12924,n12925 );
   nor U12976 ( n12925,n12746,n12873 );
   and U12977 ( n12924,datai_22_,n12883 );
   nor U12978 ( n12927,n12928,n12929 );
   nor U12979 ( n12929,n12930,n8729 );
   nor U12980 ( n12928,n12592,n12880 );
   not U12981 ( n12592,datai_7_ );
   nor U12982 ( n12926,n12931,n12932 );
   nor U12983 ( n12932,n12751,n12873 );
   and U12984 ( n12931,datai_23_,n12883 );
   nor U12985 ( n12934,n12935,n12936 );
   nor U12986 ( n12936,n12937,n8730 );
   nor U12987 ( n12935,n12587,n12880 );
   not U12988 ( n12587,datai_8_ );
   nor U12989 ( n12933,n12938,n12939 );
   nor U12990 ( n12939,n12756,n12873 );
   and U12991 ( n12938,datai_24_,n12883 );
   nor U12992 ( n12941,n12942,n12943 );
   nor U12993 ( n12943,n12944,n8728 );
   nor U12994 ( n12942,n12582,n12880 );
   not U12995 ( n12582,datai_9_ );
   nor U12996 ( n12940,n12945,n12946 );
   nor U12997 ( n12946,n12761,n12873 );
   and U12998 ( n12945,datai_25_,n12883 );
   nor U12999 ( n12948,n12949,n12950 );
   nor U13000 ( n12950,n12951,n8729 );
   nor U13001 ( n12949,n12577,n12880 );
   not U13002 ( n12577,datai_10_ );
   nor U13003 ( n12947,n12952,n12953 );
   nor U13004 ( n12953,n12766,n12873 );
   and U13005 ( n12952,datai_26_,n12883 );
   nor U13006 ( n12955,n12956,n12957 );
   nor U13007 ( n12957,n12958,n8730 );
   nor U13008 ( n12956,n12572,n12880 );
   not U13009 ( n12572,datai_11_ );
   nor U13010 ( n12954,n12959,n12960 );
   nor U13011 ( n12960,n12771,n12873 );
   and U13012 ( n12959,datai_27_,n12883 );
   nor U13013 ( n12962,n12963,n12964 );
   nor U13014 ( n12964,n12965,n8728 );
   nor U13015 ( n12963,n12567,n12880 );
   not U13016 ( n12567,datai_12_ );
   nor U13017 ( n12961,n12966,n12967 );
   nor U13018 ( n12967,n12776,n12873 );
   and U13019 ( n12966,datai_28_,n12883 );
   nor U13020 ( n12969,n12970,n12971 );
   nor U13021 ( n12971,n12972,n8729 );
   nor U13022 ( n12970,n12562,n12880 );
   not U13023 ( n12562,datai_13_ );
   nor U13024 ( n12968,n12973,n12974 );
   nor U13025 ( n12974,n12781,n12873 );
   and U13026 ( n12973,datai_29_,n12883 );
   nor U13027 ( n12976,n12977,n12978 );
   nor U13028 ( n12978,n12979,n8729 );
   nand U13029 ( n12980,n10745,n11722 );
   nor U13030 ( n12977,n12557,n12880 );
   nand U13031 ( n12880,n12981,n12386 );
   nor U13032 ( n12981,n11661,n12794 );
   not U13033 ( n12557,datai_14_ );
   nor U13034 ( n12975,n12982,n12983 );
   nor U13035 ( n12983,n12786,n12873 );
   and U13036 ( n12982,datai_30_,n12883 );
   nand U13037 ( n12985,n12883,datai_31_ );
   nor U13038 ( n12883,n11748,n12794 );
   nor U13039 ( n12984,n12986,n12987 );
   and U13040 ( n12987,eax_reg_31_,n8813 );
   nor U13041 ( n12986,n12794,n12988 );
   nand U13042 ( n12988,n11661,n12308 );
   not U13043 ( n12794,n12873 );
   nand U13044 ( n12873,n12989,n12990 );
   nand U13045 ( n12990,n12991,n10912 );
   nor U13046 ( n10912,n10890,n12992 );
   nor U13047 ( n12991,ready_n,n11745 );
   nand U13048 ( n12989,n12993,n12994 );
   nor U13049 ( n12993,n12995,n12996 );
   nor U13050 ( n12995,n12997,n12998 );
   nand U13051 ( n12998,n12999,n13000 );
   nand U13052 ( n12999,n13001,n9367 );
   nor U13053 ( n13001,n9393,n11631 );
   nor U13054 ( n12997,n13002,n13003 );
   nand U13055 ( n13003,n11741,n8862 );
   nand U13056 ( n13005,ebx_reg_0_,n8797 );
   nor U13057 ( n13004,n13007,n13008 );
   nor U13058 ( n13008,n10936,n8726 );
   nor U13059 ( n13007,n11763,n8734 );
   nand U13060 ( n13011,ebx_reg_1_,n8797 );
   nor U13061 ( n13010,n13012,n13013 );
   nor U13062 ( n13013,n10952,n8727 );
   not U13063 ( n10952,n13014 );
   nor U13064 ( n13012,n11769,n8734 );
   nand U13065 ( n13016,ebx_reg_2_,n13006 );
   nor U13066 ( n13015,n13017,n13018 );
   nor U13067 ( n13018,n10982,n8727 );
   not U13068 ( n10982,n13019 );
   nor U13069 ( n13017,n12806,n8732 );
   not U13070 ( n12806,n11791 );
   nand U13071 ( n13021,ebx_reg_3_,n8797 );
   nor U13072 ( n13020,n13022,n13023 );
   nor U13073 ( n13023,n11004,n8726 );
   not U13074 ( n11004,n13024 );
   nor U13075 ( n13022,n12811,n8732 );
   not U13076 ( n12811,n11813 );
   nand U13077 ( n13026,ebx_reg_4_,n13006 );
   nor U13078 ( n13025,n13027,n13028 );
   nor U13079 ( n13028,n11032,n13009 );
   nor U13080 ( n13027,n12816,n8733 );
   not U13081 ( n12816,n11834 );
   nand U13082 ( n13030,ebx_reg_5_,n13006 );
   nor U13083 ( n13029,n13031,n13032 );
   nor U13084 ( n13032,n11051,n8727 );
   not U13085 ( n11051,n13033 );
   nor U13086 ( n13031,n12821,n8733 );
   not U13087 ( n12821,n11849 );
   nand U13088 ( n13035,ebx_reg_6_,n13006 );
   nor U13089 ( n13034,n13036,n13037 );
   nor U13090 ( n13037,n11079,n8726 );
   nor U13091 ( n13036,n12826,n8734 );
   nand U13092 ( n13039,ebx_reg_7_,n13006 );
   nor U13093 ( n13038,n13040,n13041 );
   nor U13094 ( n13041,n11098,n13009 );
   not U13095 ( n11098,n13042 );
   nor U13096 ( n13040,n12831,n8734 );
   nand U13097 ( n13044,ebx_reg_8_,n13006 );
   nor U13098 ( n13043,n13045,n13046 );
   nor U13099 ( n13046,n11125,n8727 );
   nor U13100 ( n13045,n12836,n8732 );
   not U13101 ( n12836,n11904 );
   nand U13102 ( n13048,ebx_reg_9_,n13006 );
   nor U13103 ( n13047,n13049,n13050 );
   nor U13104 ( n13050,n11144,n8726 );
   not U13105 ( n11144,n13051 );
   nor U13106 ( n13049,n12841,n8732 );
   not U13107 ( n12841,n11919 );
   nand U13108 ( n13053,ebx_reg_10_,n13006 );
   nor U13109 ( n13052,n13054,n13055 );
   nor U13110 ( n13055,n11171,n13009 );
   nor U13111 ( n13054,n12846,n8733 );
   not U13112 ( n12846,n11937 );
   nand U13113 ( n13057,ebx_reg_11_,n13006 );
   nor U13114 ( n13056,n13058,n13059 );
   nor U13115 ( n13059,n11190,n8727 );
   not U13116 ( n11190,n13060 );
   nor U13117 ( n13058,n12851,n8733 );
   not U13118 ( n12851,n11955 );
   nand U13119 ( n13062,ebx_reg_12_,n13006 );
   nor U13120 ( n13061,n13063,n13064 );
   nor U13121 ( n13064,n11217,n8726 );
   nor U13122 ( n13063,n12856,n8733 );
   not U13123 ( n12856,n11975 );
   nand U13124 ( n13066,ebx_reg_13_,n13006 );
   nor U13125 ( n13065,n13067,n13068 );
   nor U13126 ( n13068,n11236,n13009 );
   not U13127 ( n11236,n13069 );
   nor U13128 ( n13067,n12861,n8734 );
   nand U13129 ( n13071,ebx_reg_14_,n13006 );
   nor U13130 ( n13070,n13072,n13073 );
   nor U13131 ( n13073,n11263,n13009 );
   nor U13132 ( n13072,n12866,n8734 );
   not U13133 ( n12866,n12005 );
   nand U13134 ( n13075,ebx_reg_15_,n13006 );
   nor U13135 ( n13074,n13076,n13077 );
   nor U13136 ( n13077,n11282,n8726 );
   not U13137 ( n11282,n13078 );
   nor U13138 ( n13076,n12871,n8733 );
   nand U13139 ( n13080,ebx_reg_16_,n13006 );
   nor U13140 ( n13079,n13081,n13082 );
   nor U13141 ( n13082,n11309,n8727 );
   nor U13142 ( n13081,n12879,n8733 );
   nand U13143 ( n13084,ebx_reg_17_,n13006 );
   nor U13144 ( n13083,n13085,n13086 );
   nor U13145 ( n13086,n11328,n13009 );
   not U13146 ( n11328,n13087 );
   nor U13147 ( n13085,n12888,n8732 );
   nand U13148 ( n13089,ebx_reg_18_,n8797 );
   nor U13149 ( n13088,n13090,n13091 );
   nor U13150 ( n13091,n11355,n8726 );
   nor U13151 ( n13090,n12895,n8732 );
   not U13152 ( n12895,n12065 );
   nand U13153 ( n13093,ebx_reg_19_,n8797 );
   nor U13154 ( n13092,n13094,n13095 );
   nor U13155 ( n13095,n11374,n13009 );
   not U13156 ( n11374,n13096 );
   nor U13157 ( n13094,n12902,n8732 );
   not U13158 ( n12902,n12084 );
   nand U13159 ( n13098,ebx_reg_20_,n8797 );
   nor U13160 ( n13097,n13099,n13100 );
   nor U13161 ( n13100,n11403,n8727 );
   nor U13162 ( n13099,n12909,n8733 );
   nand U13163 ( n13102,ebx_reg_21_,n8797 );
   nor U13164 ( n13101,n13103,n13104 );
   nor U13165 ( n13104,n11422,n8726 );
   not U13166 ( n11422,n13105 );
   nor U13167 ( n13103,n12916,n8733 );
   not U13168 ( n12916,n12119 );
   nand U13169 ( n13107,ebx_reg_22_,n8797 );
   nor U13170 ( n13106,n13108,n13109 );
   nor U13171 ( n13109,n11448,n13009 );
   nor U13172 ( n13108,n12923,n8734 );
   nand U13173 ( n13111,ebx_reg_23_,n8797 );
   nor U13174 ( n13110,n13112,n13113 );
   nor U13175 ( n13113,n11467,n8727 );
   not U13176 ( n11467,n13114 );
   nor U13177 ( n13112,n12930,n8734 );
   nand U13178 ( n13116,ebx_reg_24_,n8797 );
   nor U13179 ( n13115,n13117,n13118 );
   nor U13180 ( n13118,n11495,n8726 );
   nor U13181 ( n13117,n12937,n8732 );
   not U13182 ( n12937,n12175 );
   nand U13183 ( n13120,ebx_reg_25_,n8797 );
   nor U13184 ( n13119,n13121,n13122 );
   nor U13185 ( n13122,n11514,n13009 );
   not U13186 ( n11514,n13123 );
   nor U13187 ( n13121,n12944,n8732 );
   not U13188 ( n12944,n12203 );
   nand U13189 ( n13125,ebx_reg_26_,n8797 );
   nor U13190 ( n13124,n13126,n13127 );
   nor U13191 ( n13127,n11541,n8727 );
   nor U13192 ( n13126,n12951,n8733 );
   not U13193 ( n12951,n12222 );
   nand U13194 ( n13129,ebx_reg_27_,n8797 );
   nor U13195 ( n13128,n13130,n13131 );
   nor U13196 ( n13131,n11559,n8726 );
   not U13197 ( n11559,n13132 );
   nor U13198 ( n13130,n12958,n8733 );
   nand U13199 ( n13134,ebx_reg_28_,n8797 );
   nor U13200 ( n13133,n13135,n13136 );
   nor U13201 ( n13136,n11584,n13009 );
   nor U13202 ( n13135,n12965,n8734 );
   nand U13203 ( n13138,ebx_reg_29_,n8797 );
   nor U13204 ( n13137,n13139,n13140 );
   nor U13205 ( n13140,n11597,n8727 );
   not U13206 ( n11597,n13141 );
   nor U13207 ( n13139,n12972,n8734 );
   not U13208 ( n12972,n12278 );
   nand U13209 ( n13143,ebx_reg_30_,n8797 );
   nor U13210 ( n13142,n13144,n13145 );
   nor U13211 ( n13145,n11610,n8726 );
   not U13212 ( n13009,n13146 );
   not U13213 ( n11610,n13147 );
   nor U13214 ( n13144,n12979,n8732 );
   nand U13215 ( n13149,n13146,n13150 );
   nor U13216 ( n13146,n13006,n10745 );
   nand U13217 ( n13148,ebx_reg_31_,n8797 );
   nand U13218 ( n13006,n9287,n13151 );
   nand U13219 ( n13151,n10917,n13152 );
   or U13220 ( n13152,n13000,n12992 );
   nand U13221 ( n13000,n13153,n13154 );
   nor U13222 ( n13154,n10778,n10745 );
   nor U13223 ( n13153,n13155,n13156 );
   nand U13224 ( n10917,n10877,n9393 );
   nor U13225 ( n13158,n13159,n13160 );
   nand U13226 ( n13160,n13161,n13162 );
   nand U13227 ( n13162,phyaddrpointer_reg_0_,n13163 );
   nand U13228 ( n13163,n13164,n8826 );
   nand U13229 ( n13161,reip_reg_0_,n13166 );
   nand U13230 ( n13166,n13167,n8782 );
   nor U13231 ( n13159,n13169,n11763 );
   xor U13232 ( n11763,n8831,n13170 );
   nand U13233 ( n13170,n13171,n13172 );
   nor U13234 ( n13157,n13173,n13174 );
   nand U13235 ( n13174,n13175,n13176 );
   nand U13236 ( n13176,n8824,n13178 );
   not U13237 ( n13178,n10936 );
   xor U13238 ( n10936,n13179,n13180 );
   nand U13239 ( n13175,n13181,n9348 );
   nor U13240 ( n13173,n13182,n13183 );
   nor U13241 ( n13185,n13186,n13187 );
   nand U13242 ( n13187,n13188,n13189 );
   or U13243 ( n13189,n11769,n13169 );
   not U13244 ( n13169,n13190 );
   xor U13245 ( n11769,n13191,n13192 );
   nand U13246 ( n13192,n13193,n13194 );
   nand U13247 ( n13188,n13177,n13014 );
   xor U13248 ( n13014,n13195,n13196 );
   xor U13249 ( n13196,n13197,n13198 );
   nor U13250 ( n13186,n8920,n13199 );
   nor U13251 ( n13184,n13200,n13201 );
   nand U13252 ( n13201,n13202,n13203 );
   nand U13253 ( n13203,n8822,ebx_reg_1_ );
   nor U13254 ( n13202,n13205,n13206 );
   nor U13255 ( n13206,n9192,n13167 );
   nor U13256 ( n13205,reip_reg_1_,n8782 );
   nand U13257 ( n13200,n13207,n13208 );
   nand U13258 ( n13208,n13209,n11779 );
   nand U13259 ( n13207,n8798,phyaddrpointer_reg_1_ );
   nor U13260 ( n13212,n13213,n13214 );
   nand U13261 ( n13214,n13215,n13216 );
   nand U13262 ( n13216,n13181,n10123 );
   nand U13263 ( n13215,n13209,n13217 );
   nand U13264 ( n13213,n13218,n13219 );
   nand U13265 ( n13219,n13190,n11791 );
   nand U13266 ( n11791,n13220,n13221 );
   nand U13267 ( n13221,n13222,n13223 );
   nand U13268 ( n13222,n13224,n13225 );
   or U13269 ( n13220,n13226,n13227 );
   nand U13270 ( n13218,n13177,n13019 );
   xor U13271 ( n13019,n13228,n13229 );
   nor U13272 ( n13211,n13230,n13231 );
   nand U13273 ( n13231,n13232,n13233 );
   nand U13274 ( n13233,n13210,phyaddrpointer_reg_2_ );
   nand U13275 ( n13232,n13204,ebx_reg_2_ );
   nand U13276 ( n13230,n13234,n13235 );
   nand U13277 ( n13235,reip_reg_2_,n13236 );
   nand U13278 ( n13234,n13237,n9187 );
   nor U13279 ( n13237,n9192,n8782 );
   nor U13280 ( n13239,n13240,n13241 );
   nand U13281 ( n13241,n13242,n13243 );
   nand U13282 ( n13243,n13181,n10466 );
   nand U13283 ( n13242,n13209,n11814 );
   nand U13284 ( n13240,n13244,n13245 );
   nand U13285 ( n13245,n11813,n13190 );
   xor U13286 ( n11813,n13246,n13226 );
   nand U13287 ( n13226,n13225,n13247 );
   nand U13288 ( n13247,n13223,n13224 );
   nand U13289 ( n13223,n13193,n13248 );
   nand U13290 ( n13248,n13191,n13194 );
   nand U13291 ( n13191,n13172,n13249 );
   nand U13292 ( n13249,n8831,n13171 );
   nor U13293 ( n13246,n13250,n13251 );
   not U13294 ( n13250,n13252 );
   nand U13295 ( n13244,n13177,n13024 );
   xor U13296 ( n13024,n13253,n13254 );
   nor U13297 ( n13238,n13255,n13256 );
   nand U13298 ( n13256,n13257,n13258 );
   nand U13299 ( n13258,n8798,phyaddrpointer_reg_3_ );
   nand U13300 ( n13257,n8822,ebx_reg_3_ );
   nand U13301 ( n13255,n13259,n13260 );
   nand U13302 ( n13260,reip_reg_3_,n13261 );
   nand U13303 ( n13261,n13262,n13263 );
   nand U13304 ( n13263,n8747,n9187 );
   not U13305 ( n9187,reip_reg_2_ );
   not U13306 ( n13262,n13236 );
   nand U13307 ( n13236,n8774,n13264 );
   nand U13308 ( n13264,n8745,n9192 );
   nand U13309 ( n13259,n13265,n9182 );
   nor U13310 ( n13265,n13168,n13266 );
   nand U13311 ( n13266,reip_reg_2_,reip_reg_1_ );
   nor U13312 ( n13268,n13269,n13270 );
   nand U13313 ( n13270,n13271,n13272 );
   nand U13314 ( n13272,n13177,n13273 );
   not U13315 ( n13273,n11032 );
   nand U13316 ( n11032,n13274,n13275 );
   nand U13317 ( n13274,n13276,n13277 );
   nand U13318 ( n13271,n13181,n10919 );
   not U13319 ( n13181,n13199 );
   nand U13320 ( n13199,n13278,n13279 );
   nand U13321 ( n13269,n13280,n13281 );
   nand U13322 ( n13280,n11834,n13190 );
   xor U13323 ( n11834,n13282,n13283 );
   and U13324 ( n13282,n13284,n13285 );
   nor U13325 ( n13267,n13286,n13287 );
   nand U13326 ( n13287,n13288,n13289 );
   nand U13327 ( n13289,n8822,ebx_reg_4_ );
   nor U13328 ( n13288,n13290,n13291 );
   nor U13329 ( n13291,reip_reg_4_,n13292 );
   nand U13330 ( n13292,n13293,n8747 );
   nor U13331 ( n13290,n13294,n9177 );
   nand U13332 ( n13286,n13295,n13296 );
   nand U13333 ( n13296,n13209,n13297 );
   nand U13334 ( n13295,n8798,phyaddrpointer_reg_4_ );
   nor U13335 ( n13299,n13300,n13301 );
   nand U13336 ( n13301,n13302,n13303 );
   nand U13337 ( n13303,n13177,n13033 );
   xor U13338 ( n13033,n13275,n13304 );
   or U13339 ( n13302,n8826,n11850 );
   nand U13340 ( n13300,n13305,n13281 );
   nand U13341 ( n13305,n13190,n11849 );
   nand U13342 ( n11849,n13306,n13307 );
   nand U13343 ( n13307,n13308,n13309 );
   nand U13344 ( n13308,n13310,n13311 );
   nand U13345 ( n13306,n13312,n13311 );
   not U13346 ( n13312,n13313 );
   nand U13347 ( n13190,n13314,n13315 );
   nand U13348 ( n13315,n13279,n8845 );
   nor U13349 ( n13298,n13316,n13317 );
   nand U13350 ( n13317,n13318,n13319 );
   nand U13351 ( n13319,n8798,phyaddrpointer_reg_5_ );
   nand U13352 ( n13318,n8822,ebx_reg_5_ );
   nand U13353 ( n13316,n13320,n13321 );
   nand U13354 ( n13321,reip_reg_5_,n13322 );
   nand U13355 ( n13322,n13294,n13323 );
   nand U13356 ( n13323,n8747,n9177 );
   and U13357 ( n13294,n13167,n13324 );
   nand U13358 ( n13324,n8746,n13325 );
   nand U13359 ( n13320,n13326,n9172 );
   nor U13360 ( n13326,n13325,n13327 );
   nand U13361 ( n13327,n8746,reip_reg_4_ );
   nor U13362 ( n13329,n13330,n13331 );
   nand U13363 ( n13331,n13332,n13333 );
   nand U13364 ( n13333,n13177,n13334 );
   not U13365 ( n13334,n11079 );
   nand U13366 ( n11079,n13335,n13336 );
   nand U13367 ( n13335,n13337,n13338 );
   or U13368 ( n13332,n8825,n11865 );
   nand U13369 ( n13330,n13339,n13281 );
   nand U13370 ( n13339,n8819,n11864 );
   not U13371 ( n11864,n12826 );
   nand U13372 ( n12826,n13341,n13342 );
   or U13373 ( n13342,n13343,n13344 );
   nor U13374 ( n13328,n13345,n13346 );
   nand U13375 ( n13346,n13347,n13348 );
   nand U13376 ( n13348,n8798,phyaddrpointer_reg_6_ );
   nand U13377 ( n13347,n8822,ebx_reg_6_ );
   nand U13378 ( n13345,n13349,n13350 );
   nand U13379 ( n13350,reip_reg_6_,n13351 );
   nand U13380 ( n13349,n13352,n9167 );
   nor U13381 ( n13352,n8782,n13353 );
   nor U13382 ( n13355,n13356,n13357 );
   nand U13383 ( n13357,n13358,n13359 );
   nand U13384 ( n13359,n13177,n13042 );
   xor U13385 ( n13042,n13360,n13336 );
   nand U13386 ( n13358,n13209,n11881 );
   nand U13387 ( n13356,n13361,n13281 );
   nand U13388 ( n13361,n13340,n11880 );
   not U13389 ( n11880,n12831 );
   nand U13390 ( n12831,n13362,n13363 );
   nand U13391 ( n13363,n13364,n13341 );
   nand U13392 ( n13341,n13344,n13343 );
   nand U13393 ( n13362,n13365,n13344 );
   nand U13394 ( n13344,n13310,n13366 );
   nand U13395 ( n13366,n13309,n13311 );
   not U13396 ( n13365,n13367 );
   nor U13397 ( n13354,n13368,n13369 );
   nand U13398 ( n13369,n13370,n13371 );
   nand U13399 ( n13371,n8798,phyaddrpointer_reg_7_ );
   nand U13400 ( n13370,n8822,ebx_reg_7_ );
   nand U13401 ( n13368,n13372,n13373 );
   nand U13402 ( n13373,reip_reg_7_,n13374 );
   nand U13403 ( n13374,n13375,n13376 );
   nand U13404 ( n13376,n8745,n9167 );
   not U13405 ( n9167,reip_reg_6_ );
   not U13406 ( n13375,n13351 );
   nand U13407 ( n13351,n13167,n13377 );
   nand U13408 ( n13377,n8745,n13353 );
   nand U13409 ( n13372,n13378,n9162 );
   not U13410 ( n9162,reip_reg_7_ );
   nor U13411 ( n13378,n13353,n13379 );
   nand U13412 ( n13379,n8747,reip_reg_6_ );
   nor U13413 ( n13381,n13382,n13383 );
   nand U13414 ( n13383,n13384,n13385 );
   nand U13415 ( n13385,n13177,n13386 );
   not U13416 ( n13386,n11125 );
   nand U13417 ( n11125,n13387,n13388 );
   nand U13418 ( n13387,n13389,n13390 );
   or U13419 ( n13384,n8825,n11905 );
   nand U13420 ( n13382,n13391,n13281 );
   nand U13421 ( n13391,n8819,n11904 );
   xor U13422 ( n11904,n13392,n13393 );
   nor U13423 ( n13380,n13394,n13395 );
   nand U13424 ( n13395,n13396,n13397 );
   nand U13425 ( n13397,n8798,phyaddrpointer_reg_8_ );
   nand U13426 ( n13396,n8822,ebx_reg_8_ );
   nand U13427 ( n13394,n13398,n13399 );
   nand U13428 ( n13399,reip_reg_8_,n13400 );
   nand U13429 ( n13398,n13401,n9157 );
   nor U13430 ( n13401,n13168,n13402 );
   nor U13431 ( n13404,n13405,n13406 );
   nand U13432 ( n13406,n13407,n13408 );
   nand U13433 ( n13408,n13177,n13051 );
   xor U13434 ( n13051,n13409,n13388 );
   or U13435 ( n13407,n13165,n11920 );
   nand U13436 ( n13405,n13410,n13281 );
   nand U13437 ( n13410,n8819,n11919 );
   xor U13438 ( n11919,n13411,n13412 );
   nor U13439 ( n13403,n13413,n13414 );
   nand U13440 ( n13414,n13415,n13416 );
   nand U13441 ( n13416,n8798,phyaddrpointer_reg_9_ );
   nand U13442 ( n13415,n8822,ebx_reg_9_ );
   nand U13443 ( n13413,n13417,n13418 );
   nand U13444 ( n13418,reip_reg_9_,n13419 );
   nand U13445 ( n13419,n13420,n13421 );
   nand U13446 ( n13421,n8747,n9157 );
   not U13447 ( n13420,n13400 );
   nand U13448 ( n13400,n13167,n13422 );
   nand U13449 ( n13422,n8746,n13402 );
   nand U13450 ( n13417,n13423,n9152 );
   nor U13451 ( n13423,n13402,n13424 );
   nand U13452 ( n13424,n8746,reip_reg_8_ );
   not U13453 ( n13402,n13425 );
   nor U13454 ( n13427,n13428,n13429 );
   nand U13455 ( n13429,n13430,n13431 );
   nand U13456 ( n13431,n13177,n13432 );
   not U13457 ( n13432,n11171 );
   nand U13458 ( n11171,n13433,n13434 );
   nand U13459 ( n13433,n13435,n13436 );
   or U13460 ( n13430,n13165,n11938 );
   nand U13461 ( n13428,n13437,n13281 );
   nand U13462 ( n13437,n8819,n11937 );
   xor U13463 ( n11937,n13438,n13439 );
   nor U13464 ( n13426,n13440,n13441 );
   nand U13465 ( n13441,n13442,n13443 );
   nand U13466 ( n13443,n8798,phyaddrpointer_reg_10_ );
   nand U13467 ( n13442,n8822,ebx_reg_10_ );
   nand U13468 ( n13440,n13444,n13445 );
   nand U13469 ( n13445,reip_reg_10_,n13446 );
   nand U13470 ( n13444,n13447,n9147 );
   nor U13471 ( n13447,n8782,n13448 );
   nor U13472 ( n13450,n13451,n13452 );
   nand U13473 ( n13452,n13453,n13454 );
   nand U13474 ( n13454,n13177,n13060 );
   xor U13475 ( n13060,n13455,n13434 );
   nand U13476 ( n13453,n13209,n11956 );
   nand U13477 ( n13451,n13456,n13281 );
   nand U13478 ( n13456,n8819,n11955 );
   xor U13479 ( n11955,n13457,n13458 );
   nor U13480 ( n13457,n13438,n13439 );
   nand U13481 ( n13439,n13459,n13460 );
   nand U13482 ( n13459,n13461,n13411 );
   nor U13483 ( n13449,n13462,n13463 );
   nand U13484 ( n13463,n13464,n13465 );
   nand U13485 ( n13465,n8798,phyaddrpointer_reg_11_ );
   nand U13486 ( n13464,n8822,ebx_reg_11_ );
   nand U13487 ( n13462,n13466,n13467 );
   nand U13488 ( n13467,reip_reg_11_,n13468 );
   nand U13489 ( n13468,n13469,n13470 );
   nand U13490 ( n13470,n8745,n9147 );
   not U13491 ( n9147,reip_reg_10_ );
   not U13492 ( n13469,n13446 );
   nand U13493 ( n13446,n13167,n13471 );
   nand U13494 ( n13471,n8745,n13448 );
   nand U13495 ( n13466,n13472,n9142 );
   not U13496 ( n9142,reip_reg_11_ );
   nor U13497 ( n13472,n13448,n13473 );
   nand U13498 ( n13473,n8747,reip_reg_10_ );
   nor U13499 ( n13475,n13476,n13477 );
   nand U13500 ( n13477,n13478,n13479 );
   nand U13501 ( n13479,n13177,n13480 );
   not U13502 ( n13480,n11217 );
   nand U13503 ( n11217,n13481,n13482 );
   nand U13504 ( n13481,n13483,n13484 );
   nand U13505 ( n13478,n13209,n13485 );
   nand U13506 ( n13476,n13486,n13281 );
   nand U13507 ( n13486,n8819,n11975 );
   xor U13508 ( n11975,n13487,n13488 );
   nor U13509 ( n13474,n13489,n13490 );
   nand U13510 ( n13490,n13491,n13492 );
   nand U13511 ( n13492,n8798,phyaddrpointer_reg_12_ );
   nand U13512 ( n13491,n8822,ebx_reg_12_ );
   nand U13513 ( n13489,n13493,n13494 );
   nand U13514 ( n13494,reip_reg_12_,n13495 );
   nand U13515 ( n13493,n13496,n9137 );
   nor U13516 ( n13496,n8782,n13497 );
   nor U13517 ( n13499,n13500,n13501 );
   nand U13518 ( n13501,n13502,n13503 );
   nand U13519 ( n13503,n13177,n13069 );
   xor U13520 ( n13069,n13504,n13482 );
   nand U13521 ( n13502,n13209,n11991 );
   not U13522 ( n13209,n8826 );
   nand U13523 ( n13500,n13505,n13281 );
   nand U13524 ( n13505,n8819,n11990 );
   not U13525 ( n11990,n12861 );
   xor U13526 ( n12861,n13506,n13507 );
   nor U13527 ( n13498,n13508,n13509 );
   nand U13528 ( n13509,n13510,n13511 );
   nand U13529 ( n13511,n8798,phyaddrpointer_reg_13_ );
   nand U13530 ( n13510,n8822,ebx_reg_13_ );
   nand U13531 ( n13508,n13512,n13513 );
   nand U13532 ( n13513,reip_reg_13_,n13514 );
   nand U13533 ( n13514,n13515,n13516 );
   nand U13534 ( n13516,n8747,n9137 );
   not U13535 ( n13515,n13495 );
   nand U13536 ( n13495,n13167,n13517 );
   nand U13537 ( n13517,n8746,n13497 );
   nand U13538 ( n13512,n13518,n9132 );
   nor U13539 ( n13518,n13497,n13519 );
   nand U13540 ( n13519,n8746,reip_reg_12_ );
   not U13541 ( n13497,n13520 );
   nor U13542 ( n13522,n13523,n13524 );
   nand U13543 ( n13524,n13525,n13526 );
   nand U13544 ( n13526,n13177,n13527 );
   not U13545 ( n13527,n11263 );
   nand U13546 ( n11263,n13528,n13529 );
   nand U13547 ( n13528,n13530,n13531 );
   or U13548 ( n13525,n8825,n12006 );
   nand U13549 ( n13523,n13532,n13281 );
   nand U13550 ( n13532,n8819,n12005 );
   xor U13551 ( n12005,n13533,n13534 );
   nor U13552 ( n13521,n13535,n13536 );
   nand U13553 ( n13536,n13537,n13538 );
   nand U13554 ( n13538,n8798,phyaddrpointer_reg_14_ );
   nand U13555 ( n13537,n8822,ebx_reg_14_ );
   nand U13556 ( n13535,n13539,n13540 );
   nand U13557 ( n13540,reip_reg_14_,n13541 );
   nand U13558 ( n13539,n13542,n9127 );
   nor U13559 ( n13542,n13168,n13543 );
   nor U13560 ( n13545,n13546,n13547 );
   nand U13561 ( n13547,n13548,n13549 );
   nand U13562 ( n13549,n13177,n13078 );
   xor U13563 ( n13078,n13550,n13529 );
   or U13564 ( n13548,n13165,n12021 );
   nand U13565 ( n13546,n13551,n13281 );
   nand U13566 ( n13551,n13340,n12020 );
   not U13567 ( n12020,n12871 );
   xor U13568 ( n12871,n13552,n13553 );
   nand U13569 ( n13553,n13533,n13534 );
   and U13570 ( n13533,n13554,n13506 );
   nand U13571 ( n13554,n13507,n13555 );
   not U13572 ( n13555,n13556 );
   nor U13573 ( n13507,n13557,n13558 );
   and U13574 ( n13557,n13487,n13488 );
   nor U13575 ( n13544,n13559,n13560 );
   nand U13576 ( n13560,n13561,n13562 );
   nand U13577 ( n13562,n8798,phyaddrpointer_reg_15_ );
   nand U13578 ( n13561,n8822,ebx_reg_15_ );
   nand U13579 ( n13559,n13563,n13564 );
   nand U13580 ( n13564,reip_reg_15_,n13565 );
   nand U13581 ( n13565,n13566,n13567 );
   nand U13582 ( n13567,n8745,n9127 );
   not U13583 ( n9127,reip_reg_14_ );
   not U13584 ( n13566,n13541 );
   nand U13585 ( n13541,n13167,n13568 );
   nand U13586 ( n13568,n8745,n13543 );
   nand U13587 ( n13563,n13569,n9122 );
   not U13588 ( n9122,reip_reg_15_ );
   nor U13589 ( n13569,n13543,n13570 );
   nand U13590 ( n13570,n8746,reip_reg_14_ );
   nor U13591 ( n13572,n13573,n13574 );
   nand U13592 ( n13574,n13575,n13576 );
   nand U13593 ( n13576,n8824,n13577 );
   not U13594 ( n13577,n11309 );
   nand U13595 ( n11309,n13578,n13579 );
   nand U13596 ( n13578,n13580,n13581 );
   or U13597 ( n13575,n8826,n12036 );
   nand U13598 ( n13573,n13582,n13281 );
   nand U13599 ( n13582,n13340,n12035 );
   not U13600 ( n12035,n12879 );
   nand U13601 ( n12879,n13583,n13584 );
   nand U13602 ( n13584,n13585,n13586 );
   nand U13603 ( n13586,n13587,n13588 );
   not U13604 ( n13585,n13589 );
   nand U13605 ( n13583,n13590,n13587 );
   nor U13606 ( n13571,n13591,n13592 );
   nand U13607 ( n13592,n13593,n13594 );
   nand U13608 ( n13594,n13210,phyaddrpointer_reg_16_ );
   nand U13609 ( n13593,n13204,ebx_reg_16_ );
   nand U13610 ( n13591,n13595,n13596 );
   nand U13611 ( n13596,reip_reg_16_,n13597 );
   nand U13612 ( n13595,n13598,n9117 );
   nor U13613 ( n13598,n8782,n13599 );
   nor U13614 ( n13601,n13602,n13603 );
   nand U13615 ( n13603,n13604,n13605 );
   nand U13616 ( n13605,n8824,n13087 );
   xor U13617 ( n13087,n13606,n13579 );
   or U13618 ( n13604,n8826,n12052 );
   nand U13619 ( n13602,n13607,n13281 );
   nand U13620 ( n13607,n13340,n12051 );
   not U13621 ( n12051,n12888 );
   xor U13622 ( n12888,n13608,n13609 );
   nor U13623 ( n13600,n13610,n13611 );
   nand U13624 ( n13611,n13612,n13613 );
   nand U13625 ( n13613,n13210,phyaddrpointer_reg_17_ );
   nand U13626 ( n13612,n13204,ebx_reg_17_ );
   nand U13627 ( n13610,n13614,n13615 );
   nand U13628 ( n13615,reip_reg_17_,n13616 );
   nand U13629 ( n13616,n13617,n13618 );
   nand U13630 ( n13618,n8746,n9117 );
   not U13631 ( n13617,n13597 );
   nand U13632 ( n13597,n13167,n13619 );
   nand U13633 ( n13619,n8745,n13599 );
   nand U13634 ( n13614,n13620,n9112 );
   nor U13635 ( n13620,n13599,n13621 );
   nand U13636 ( n13621,n8747,reip_reg_16_ );
   not U13637 ( n13599,n13622 );
   nor U13638 ( n13624,n13625,n13626 );
   nand U13639 ( n13626,n13627,n13628 );
   nand U13640 ( n13628,n8824,n13629 );
   not U13641 ( n13629,n11355 );
   nand U13642 ( n11355,n13630,n13631 );
   nand U13643 ( n13630,n13632,n13633 );
   or U13644 ( n13627,n13165,n12066 );
   nand U13645 ( n13625,n13634,n13281 );
   nand U13646 ( n13634,n13340,n12065 );
   xor U13647 ( n12065,n13635,n13636 );
   nand U13648 ( n13636,n13637,n13609 );
   nand U13649 ( n13609,n13638,n13587 );
   nor U13650 ( n13623,n13639,n13640 );
   nand U13651 ( n13640,n13641,n13642 );
   nand U13652 ( n13642,n13210,phyaddrpointer_reg_18_ );
   nand U13653 ( n13641,n13204,ebx_reg_18_ );
   nand U13654 ( n13639,n13643,n13644 );
   nand U13655 ( n13644,reip_reg_18_,n13645 );
   nand U13656 ( n13643,n13646,n9107 );
   nor U13657 ( n13646,n8782,n13647 );
   nor U13658 ( n13649,n13650,n13651 );
   nand U13659 ( n13651,n13652,n13653 );
   nand U13660 ( n13653,n8824,n13096 );
   xor U13661 ( n13096,n13654,n13631 );
   or U13662 ( n13652,n8825,n12085 );
   nand U13663 ( n13650,n13655,n13281 );
   nand U13664 ( n13281,n8843,n8774 );
   nand U13665 ( n13655,n13340,n12084 );
   xor U13666 ( n12084,n13656,n13657 );
   and U13667 ( n13656,n13658,n13659 );
   nor U13668 ( n13648,n13660,n13661 );
   nand U13669 ( n13661,n13662,n13663 );
   nand U13670 ( n13663,n13210,phyaddrpointer_reg_19_ );
   nand U13671 ( n13662,n13204,ebx_reg_19_ );
   nand U13672 ( n13660,n13664,n13665 );
   nand U13673 ( n13665,reip_reg_19_,n13666 );
   nand U13674 ( n13666,n13667,n13668 );
   nand U13675 ( n13668,n8745,n9107 );
   not U13676 ( n9107,reip_reg_18_ );
   not U13677 ( n13667,n13645 );
   nand U13678 ( n13645,n13167,n13669 );
   nand U13679 ( n13669,n8745,n13647 );
   nand U13680 ( n13664,n13670,n9102 );
   not U13681 ( n9102,reip_reg_19_ );
   nor U13682 ( n13670,n13647,n13671 );
   nand U13683 ( n13671,n8746,reip_reg_18_ );
   nor U13684 ( n13673,n13674,n13675 );
   nand U13685 ( n13675,n13676,n13677 );
   nand U13686 ( n13677,n13340,n12102 );
   not U13687 ( n12102,n12909 );
   xor U13688 ( n12909,n13678,n13679 );
   nand U13689 ( n13676,n8824,n13680 );
   not U13690 ( n13680,n11403 );
   nand U13691 ( n11403,n13681,n13682 );
   nand U13692 ( n13681,n13683,n13684 );
   nor U13693 ( n13674,n12103,n8825 );
   nor U13694 ( n13672,n13685,n13686 );
   nand U13695 ( n13686,n13687,n13688 );
   nand U13696 ( n13688,n13210,phyaddrpointer_reg_20_ );
   nand U13697 ( n13687,n13204,ebx_reg_20_ );
   nand U13698 ( n13685,n13689,n13690 );
   nand U13699 ( n13690,reip_reg_20_,n13691 );
   nand U13700 ( n13689,n13692,n9097 );
   nor U13701 ( n13692,n13168,n13693 );
   nor U13702 ( n13695,n13696,n13697 );
   nand U13703 ( n13697,n13698,n13699 );
   nand U13704 ( n13699,n13340,n12119 );
   xor U13705 ( n12119,n13700,n13701 );
   nand U13706 ( n13698,n8824,n13105 );
   xor U13707 ( n13105,n13702,n13682 );
   nor U13708 ( n13696,n12120,n8826 );
   nor U13709 ( n13694,n13703,n13704 );
   nand U13710 ( n13704,n13705,n13706 );
   nand U13711 ( n13706,n13210,phyaddrpointer_reg_21_ );
   nand U13712 ( n13705,n13204,ebx_reg_21_ );
   nand U13713 ( n13703,n13707,n13708 );
   nand U13714 ( n13708,reip_reg_21_,n13709 );
   nand U13715 ( n13709,n13710,n13711 );
   nand U13716 ( n13711,n8746,n9097 );
   not U13717 ( n13710,n13691 );
   nand U13718 ( n13691,n13167,n13712 );
   nand U13719 ( n13712,n8747,n13693 );
   nand U13720 ( n13707,n13713,n9092 );
   nor U13721 ( n13713,n13693,n13714 );
   nand U13722 ( n13714,n8747,reip_reg_20_ );
   not U13723 ( n13693,n13715 );
   nor U13724 ( n13717,n13718,n13719 );
   nand U13725 ( n13719,n13720,n13721 );
   nand U13726 ( n13721,n13340,n12140 );
   not U13727 ( n12140,n12923 );
   xor U13728 ( n12923,n13722,n13723 );
   nor U13729 ( n13722,n13700,n13701 );
   nand U13730 ( n13701,n13724,n13679 );
   nand U13731 ( n13724,n13678,n13725 );
   nand U13732 ( n13725,n13726,n13727 );
   nand U13733 ( n13720,n8824,n13728 );
   not U13734 ( n13728,n11448 );
   nand U13735 ( n11448,n13729,n13730 );
   nand U13736 ( n13729,n13731,n13732 );
   nor U13737 ( n13718,n12141,n8825 );
   nor U13738 ( n13716,n13733,n13734 );
   nand U13739 ( n13734,n13735,n13736 );
   nand U13740 ( n13736,n13210,phyaddrpointer_reg_22_ );
   nand U13741 ( n13735,n13204,ebx_reg_22_ );
   nand U13742 ( n13733,n13737,n13738 );
   nand U13743 ( n13738,reip_reg_22_,n13739 );
   nand U13744 ( n13737,n13740,n9087 );
   nor U13745 ( n13740,n13168,n13741 );
   nor U13746 ( n13743,n13744,n13745 );
   nand U13747 ( n13745,n13746,n13747 );
   nand U13748 ( n13747,n13340,n12158 );
   not U13749 ( n12158,n12930 );
   xor U13750 ( n12930,n13748,n13749 );
   nand U13751 ( n13746,n8824,n13114 );
   xor U13752 ( n13114,n13750,n13730 );
   nor U13753 ( n13744,n12159,n13165 );
   nor U13754 ( n13742,n13751,n13752 );
   nand U13755 ( n13752,n13753,n13754 );
   nand U13756 ( n13754,n13210,phyaddrpointer_reg_23_ );
   nand U13757 ( n13753,n13204,ebx_reg_23_ );
   nand U13758 ( n13751,n13755,n13756 );
   nand U13759 ( n13756,reip_reg_23_,n13757 );
   nand U13760 ( n13757,n13758,n13759 );
   nand U13761 ( n13759,n8745,n9087 );
   not U13762 ( n9087,reip_reg_22_ );
   not U13763 ( n13758,n13739 );
   nand U13764 ( n13739,n13167,n13760 );
   nand U13765 ( n13760,n8745,n13741 );
   nand U13766 ( n13755,n13761,n9082 );
   not U13767 ( n9082,reip_reg_23_ );
   nor U13768 ( n13761,n13741,n13762 );
   nand U13769 ( n13762,n8747,reip_reg_22_ );
   nor U13770 ( n13764,n13765,n13766 );
   nand U13771 ( n13766,n13767,n13768 );
   nand U13772 ( n13768,n13340,n12175 );
   xor U13773 ( n12175,n13769,n13770 );
   nand U13774 ( n13770,n13771,n13749 );
   nand U13775 ( n13749,n13772,n13773 );
   nand U13776 ( n13773,n13774,n13775 );
   nor U13777 ( n13775,n13776,n13678 );
   nor U13778 ( n13774,n13700,n13723 );
   not U13779 ( n13700,n13777 );
   not U13780 ( n13771,n13748 );
   nand U13781 ( n13767,n8824,n13778 );
   not U13782 ( n13778,n11495 );
   nand U13783 ( n11495,n13779,n13780 );
   nand U13784 ( n13779,n13781,n13782 );
   nor U13785 ( n13765,n12176,n8825 );
   nor U13786 ( n13763,n13783,n13784 );
   nand U13787 ( n13784,n13785,n13786 );
   nand U13788 ( n13786,n13210,phyaddrpointer_reg_24_ );
   nand U13789 ( n13785,n13204,ebx_reg_24_ );
   nand U13790 ( n13783,n13787,n13788 );
   nand U13791 ( n13788,reip_reg_24_,n13789 );
   nand U13792 ( n13787,n13790,n9077 );
   nor U13793 ( n13790,n13168,n13791 );
   nor U13794 ( n13793,n13794,n13795 );
   nand U13795 ( n13795,n13796,n13797 );
   nand U13796 ( n13797,n13340,n12203 );
   xor U13797 ( n12203,n13798,n13799 );
   nand U13798 ( n13796,n8824,n13123 );
   xor U13799 ( n13123,n13800,n13780 );
   nor U13800 ( n13794,n12204,n8825 );
   nor U13801 ( n13792,n13801,n13802 );
   nand U13802 ( n13802,n13803,n13804 );
   nand U13803 ( n13804,n13210,phyaddrpointer_reg_25_ );
   nand U13804 ( n13803,n13204,ebx_reg_25_ );
   nand U13805 ( n13801,n13805,n13806 );
   nand U13806 ( n13806,reip_reg_25_,n13807 );
   nand U13807 ( n13807,n13808,n13809 );
   nand U13808 ( n13809,n8746,n9077 );
   not U13809 ( n13808,n13789 );
   nand U13810 ( n13789,n13167,n13810 );
   nand U13811 ( n13810,n8747,n13791 );
   nand U13812 ( n13805,n13811,n9072 );
   nor U13813 ( n13811,n13791,n13812 );
   nand U13814 ( n13812,n8747,reip_reg_24_ );
   not U13815 ( n13791,n13813 );
   nor U13816 ( n13815,n13816,n13817 );
   nand U13817 ( n13817,n13818,n13819 );
   nand U13818 ( n13819,n13340,n12222 );
   xor U13819 ( n12222,n13820,n13821 );
   nand U13820 ( n13818,n8824,n13822 );
   not U13821 ( n13822,n11541 );
   nand U13822 ( n11541,n13823,n13824 );
   nand U13823 ( n13823,n13825,n13826 );
   nor U13824 ( n13816,n12223,n8826 );
   nor U13825 ( n13814,n13827,n13828 );
   nand U13826 ( n13828,n13829,n13830 );
   nand U13827 ( n13830,n13210,phyaddrpointer_reg_26_ );
   nand U13828 ( n13829,n13204,ebx_reg_26_ );
   nand U13829 ( n13827,n13831,n13832 );
   nand U13830 ( n13832,reip_reg_26_,n13833 );
   nand U13831 ( n13831,n13834,n9067 );
   nor U13832 ( n13834,n8782,n13835 );
   nor U13833 ( n13837,n13838,n13839 );
   nand U13834 ( n13839,n13840,n13841 );
   nand U13835 ( n13841,n13340,n12238 );
   not U13836 ( n12238,n12958 );
   nand U13837 ( n12958,n13842,n13843 );
   nand U13838 ( n13843,n13844,n13845 );
   nand U13839 ( n13845,n13821,n13820 );
   not U13840 ( n13844,n13846 );
   nand U13841 ( n13842,n13847,n13820 );
   nand U13842 ( n13820,n13848,n13849 );
   nand U13843 ( n13840,n8824,n13132 );
   xor U13844 ( n13132,n13850,n13824 );
   nor U13845 ( n13838,n12239,n13165 );
   nor U13846 ( n13836,n13851,n13852 );
   nand U13847 ( n13852,n13853,n13854 );
   nand U13848 ( n13854,n13210,phyaddrpointer_reg_27_ );
   nand U13849 ( n13853,n13204,ebx_reg_27_ );
   nand U13850 ( n13851,n13855,n13856 );
   nand U13851 ( n13856,reip_reg_27_,n13857 );
   nand U13852 ( n13857,n13858,n13859 );
   nand U13853 ( n13859,n8745,n9067 );
   not U13854 ( n9067,reip_reg_26_ );
   not U13855 ( n13858,n13833 );
   nand U13856 ( n13833,n13167,n13860 );
   nand U13857 ( n13860,n8745,n13835 );
   nand U13858 ( n13855,n13861,n9062 );
   not U13859 ( n9062,reip_reg_27_ );
   nor U13860 ( n13861,n13835,n13862 );
   nand U13861 ( n13862,n8746,reip_reg_26_ );
   nor U13862 ( n13864,n13865,n13866 );
   nand U13863 ( n13866,n13867,n13868 );
   nand U13864 ( n13868,n13340,n12261 );
   not U13865 ( n12261,n12965 );
   xor U13866 ( n12965,n13869,n13870 );
   nand U13867 ( n13870,n13871,n13872 );
   nand U13868 ( n13872,n13873,n13847 );
   not U13869 ( n13847,n13874 );
   not U13870 ( n13871,n13875 );
   nand U13871 ( n13867,n8824,n13876 );
   not U13872 ( n13876,n11584 );
   nand U13873 ( n11584,n13877,n13878 );
   nand U13874 ( n13877,n13879,n13880 );
   nor U13875 ( n13865,n12262,n13165 );
   nor U13876 ( n13863,n13881,n13882 );
   nand U13877 ( n13882,n13883,n13884 );
   nand U13878 ( n13884,n13210,phyaddrpointer_reg_28_ );
   nand U13879 ( n13883,n13204,ebx_reg_28_ );
   nand U13880 ( n13881,n13885,n13886 );
   nand U13881 ( n13886,reip_reg_28_,n13887 );
   nand U13882 ( n13885,n13888,n9057 );
   nor U13883 ( n13888,n13168,n13889 );
   nor U13884 ( n13891,n13892,n13893 );
   nand U13885 ( n13893,n13894,n13895 );
   nand U13886 ( n13895,n13340,n12278 );
   xor U13887 ( n12278,n13896,n13897 );
   nor U13888 ( n13896,n13875,n13898 );
   nand U13889 ( n13898,n13899,n13900 );
   nand U13890 ( n13899,n13901,n13873 );
   not U13891 ( n13873,n13848 );
   nor U13892 ( n13901,n13869,n13874 );
   nand U13893 ( n13894,n8824,n13141 );
   xor U13894 ( n13141,n13902,n13878 );
   nor U13895 ( n13892,n12279,n8826 );
   nor U13896 ( n13890,n13903,n13904 );
   nand U13897 ( n13904,n13905,n13906 );
   nand U13898 ( n13906,n13210,phyaddrpointer_reg_29_ );
   nand U13899 ( n13905,n13204,ebx_reg_29_ );
   nand U13900 ( n13903,n13907,n13908 );
   or U13901 ( n13908,n13909,reip_reg_29_ );
   or U13902 ( n13907,n9052,n13910 );
   nor U13903 ( n13912,n13913,n13914 );
   nand U13904 ( n13914,n13915,n13916 );
   nand U13905 ( n13916,n13340,n12297 );
   not U13906 ( n12297,n12979 );
   xor U13907 ( n12979,n13917,n13918 );
   nor U13908 ( n13917,n13875,n13919 );
   nand U13909 ( n13919,n13900,n13920 );
   nand U13910 ( n13920,n13921,n13922 );
   nor U13911 ( n13921,n13874,n13848 );
   nand U13912 ( n13848,n13799,n13798 );
   nand U13913 ( n13798,n13923,n13924 );
   or U13914 ( n13924,n13925,n13678 );
   and U13915 ( n13678,n13926,n13927 );
   nand U13916 ( n13927,n13928,n13727 );
   nor U13917 ( n13926,n13929,n13930 );
   nor U13918 ( n13930,n13659,n13657 );
   and U13919 ( n13659,n13931,n13932 );
   nand U13920 ( n13932,n13933,n13934 );
   nand U13921 ( n13934,n13587,n13935 );
   nand U13922 ( n13935,n13727,n13936 );
   or U13923 ( n13587,n13937,n13938 );
   nand U13924 ( n13931,n13939,n13727 );
   nor U13925 ( n13923,n13940,n13941 );
   nor U13926 ( n13941,n13942,n13943 );
   nor U13927 ( n13942,n13944,n13945 );
   not U13928 ( n13940,n13772 );
   nand U13929 ( n13772,n13727,n13946 );
   nand U13930 ( n13946,n13947,n13948 );
   nor U13931 ( n13947,n13726,n13949 );
   nand U13932 ( n13900,n13727,n13950 );
   nand U13933 ( n13950,n13951,n13952 );
   nand U13934 ( n13875,n13849,n13953 );
   or U13935 ( n13953,n13954,n13943 );
   nand U13936 ( n13849,n13727,n13955 );
   nand U13937 ( n13915,n8824,n13147 );
   xor U13938 ( n13147,n13956,n13957 );
   nor U13939 ( n13913,n12298,n13165 );
   nand U13940 ( n13165,n13958,n12461 );
   nor U13941 ( n13958,n13959,n8948 );
   nor U13942 ( n13911,n13960,n13961 );
   nand U13943 ( n13961,n13962,n13963 );
   nand U13944 ( n13963,n8798,phyaddrpointer_reg_30_ );
   not U13945 ( n13210,n13164 );
   nand U13946 ( n13962,n8822,ebx_reg_30_ );
   not U13947 ( n13204,n13183 );
   nand U13948 ( n13960,n13964,n13965 );
   nand U13949 ( n13965,reip_reg_30_,n13966 );
   nand U13950 ( n13964,n13967,n9047 );
   nor U13951 ( n13967,n9052,n13909 );
   nor U13952 ( n13969,n13970,n13971 );
   nand U13953 ( n13971,n13972,n13973 );
   nand U13954 ( n13973,n8819,n12308 );
   xor U13955 ( n12308,n13974,n13975 );
   nand U13956 ( n13975,n13976,n13977 );
   nand U13957 ( n13977,eax_reg_31_,n13978 );
   nor U13958 ( n13976,n8829,n13979 );
   nor U13959 ( n13979,n8803,n12466 );
   xor U13960 ( n13974,n8830,n13980 );
   nor U13961 ( n13980,n13981,n13982 );
   nand U13962 ( n13982,n13983,n13929 );
   nor U13963 ( n13929,n13658,n13657 );
   nor U13964 ( n13657,n13928,n13727 );
   xor U13965 ( n13928,n8831,n13984 );
   nand U13966 ( n13984,n13985,n13986 );
   nor U13967 ( n13986,n13987,n13988 );
   nor U13968 ( n13988,n12085,n8764 );
   xor U13969 ( n12085,phyaddrpointer_reg_19_,n13989 );
   nor U13970 ( n13987,n13990,n13991 );
   nor U13971 ( n13990,n13992,n13993 );
   nand U13972 ( n13993,n13994,n13995 );
   nor U13973 ( n13995,n13996,n13997 );
   nand U13974 ( n13997,n13998,n13999 );
   nand U13975 ( n13999,n14000,instqueue_reg_7__3_ );
   nand U13976 ( n13998,n14001,instqueue_reg_6__3_ );
   nand U13977 ( n13996,n14002,n14003 );
   nand U13978 ( n14003,n14004,instqueue_reg_5__3_ );
   nand U13979 ( n14002,n14005,instqueue_reg_4__3_ );
   nor U13980 ( n13994,n14006,n14007 );
   nand U13981 ( n14007,n14008,n14009 );
   nand U13982 ( n14009,n14010,instqueue_reg_3__3_ );
   nand U13983 ( n14008,n14011,instqueue_reg_2__3_ );
   nand U13984 ( n14006,n14012,n14013 );
   nand U13985 ( n14013,n14014,instqueue_reg_1__3_ );
   nand U13986 ( n14012,n14015,instqueue_reg_0__3_ );
   nand U13987 ( n13992,n14016,n14017 );
   nor U13988 ( n14017,n14018,n14019 );
   nand U13989 ( n14019,n14020,n14021 );
   nand U13990 ( n14021,n14022,instqueue_reg_15__3_ );
   nand U13991 ( n14020,n14023,instqueue_reg_14__3_ );
   nand U13992 ( n14018,n14024,n14025 );
   nand U13993 ( n14025,n14026,instqueue_reg_13__3_ );
   nand U13994 ( n14024,n14027,instqueue_reg_12__3_ );
   nor U13995 ( n14016,n14028,n14029 );
   nand U13996 ( n14029,n14030,n14031 );
   nand U13997 ( n14031,n14032,instqueue_reg_11__3_ );
   nand U13998 ( n14030,n14033,instqueue_reg_10__3_ );
   nand U13999 ( n14028,n14034,n14035 );
   nand U14000 ( n14035,n14036,instqueue_reg_9__3_ );
   nand U14001 ( n14034,n14037,instqueue_reg_8__3_ );
   nor U14002 ( n13985,n14038,n14039 );
   nor U14003 ( n14039,n8801,n12731 );
   not U14004 ( n12731,eax_reg_19_ );
   nor U14005 ( n14038,n8804,n12088 );
   nand U14006 ( n13658,n13933,n13590 );
   not U14007 ( n13590,n13638 );
   nand U14008 ( n13638,n13588,n13589 );
   nand U14009 ( n13589,n14041,n14042 );
   nor U14010 ( n14042,n14043,n14044 );
   nor U14011 ( n14044,n14045,n14046 );
   nand U14012 ( n14046,n13552,n13534 );
   nor U14013 ( n14045,n14047,n13556 );
   nor U14014 ( n13556,n14048,n14049 );
   nor U14015 ( n14047,n14050,n14051 );
   nand U14016 ( n14051,n13488,n13487 );
   nand U14017 ( n13487,n14052,n14053 );
   nand U14018 ( n13488,n14054,n14055 );
   nand U14019 ( n14055,n14056,n14057 );
   nor U14020 ( n14057,n13412,n13438 );
   not U14021 ( n13438,n14058 );
   nor U14022 ( n14056,n14059,n13411 );
   nand U14023 ( n13411,n13392,n13393 );
   nand U14024 ( n13393,n14060,n14061 );
   nand U14025 ( n14061,n14062,n14063 );
   nor U14026 ( n14060,n14064,n14065 );
   nor U14027 ( n14065,n14066,n14067 );
   nand U14028 ( n14067,n14068,n14069 );
   not U14029 ( n14066,n14070 );
   nor U14030 ( n14064,n13367,n14071 );
   nand U14031 ( n14071,n13313,n13311 );
   nand U14032 ( n13311,n14072,n14073 );
   nand U14033 ( n14073,n14074,n12418 );
   not U14034 ( n12418,n14075 );
   xor U14035 ( n14072,n8831,n14076 );
   nand U14036 ( n13313,n14077,n13310 );
   nand U14037 ( n13310,n14078,n8784 );
   nor U14038 ( n14078,n14076,n14075 );
   xor U14039 ( n14075,n14079,n14080 );
   nor U14040 ( n14079,n14081,n14082 );
   and U14041 ( n14076,n14083,n14084 );
   nor U14042 ( n14084,n14085,n14086 );
   nor U14043 ( n14086,n11850,n8766 );
   xor U14044 ( n11850,phyaddrpointer_reg_5_,n14087 );
   nor U14045 ( n14085,n14088,n14089 );
   or U14046 ( n14089,n14090,n14091 );
   nor U14047 ( n14083,n14092,n14093 );
   nor U14048 ( n14093,n14040,n12664 );
   not U14049 ( n12664,eax_reg_5_ );
   nor U14050 ( n14092,n8805,n11853 );
   not U14051 ( n14077,n13309 );
   nand U14052 ( n13309,n13285,n14094 );
   nand U14053 ( n14094,n13284,n13283 );
   nand U14054 ( n13283,n13252,n14095 );
   nand U14055 ( n14095,n14096,n14097 );
   nand U14056 ( n14097,n14098,n14099 );
   nand U14057 ( n14099,n14100,n14101 );
   nand U14058 ( n14101,n8765,n13172 );
   nand U14059 ( n13172,n14102,n14103 );
   and U14060 ( n14100,n13171,n13194 );
   nand U14061 ( n13194,n14104,n14105 );
   or U14062 ( n13171,n14103,n14102 );
   and U14063 ( n14102,state2_reg_2_,n14106 );
   nand U14064 ( n14106,n10642,n11679 );
   not U14065 ( n10642,n8905 );
   nand U14066 ( n8905,n14107,n14108 );
   nand U14067 ( n14108,n12454,n14109 );
   nand U14068 ( n14107,n14110,n14111 );
   nand U14069 ( n14111,n14112,n14113 );
   nor U14070 ( n14113,n14114,n14115 );
   nor U14071 ( n14114,n10825,n11732 );
   nor U14072 ( n14112,n8863,n14116 );
   xor U14073 ( n14103,n8830,n14117 );
   nand U14074 ( n14117,n14118,n14119 );
   nor U14075 ( n14119,n14120,n14121 );
   nor U14076 ( n14121,n8801,n12637 );
   not U14077 ( n12637,eax_reg_0_ );
   nor U14078 ( n14120,n8910,n14090 );
   nor U14079 ( n14118,n14122,n14123 );
   nor U14080 ( n14123,n14124,n11758 );
   not U14081 ( n11758,phyaddrpointer_reg_0_ );
   nor U14082 ( n14124,n8831,n7819 );
   nor U14083 ( n14122,n8968,n14125 );
   and U14084 ( n14098,n13193,n13225 );
   nand U14085 ( n13225,n14126,n14127 );
   nand U14086 ( n14127,n14128,n8803 );
   nand U14087 ( n14128,n14074,n8930 );
   or U14088 ( n13193,n14105,n14104 );
   xor U14089 ( n14104,n14129,n8829 );
   nor U14090 ( n14129,n14130,n14131 );
   nand U14091 ( n14131,n14132,n14133 );
   nand U14092 ( n14133,n11710,instqueuerd_addr_reg_1_ );
   nor U14093 ( n14132,n14134,n14135 );
   nor U14094 ( n14135,n8803,n11779 );
   nor U14095 ( n14134,phyaddrpointer_reg_1_,n8765 );
   nand U14096 ( n14130,n14136,n14137 );
   nand U14097 ( n14137,n14074,n9603 );
   nand U14098 ( n14136,eax_reg_1_,n13978 );
   nand U14099 ( n14105,n14074,n8917 );
   xor U14100 ( n8917,n14110,n14138 );
   nand U14101 ( n14138,n14139,n14140 );
   nor U14102 ( n14096,n13251,n13227 );
   not U14103 ( n13227,n13224 );
   nand U14104 ( n13224,n14141,n14142 );
   xor U14105 ( n14142,n14126,n8763 );
   nand U14106 ( n14126,n14143,n14144 );
   nor U14107 ( n14144,n14145,n14146 );
   nand U14108 ( n14146,n14147,n14148 );
   nand U14109 ( n14148,n13217,n8829 );
   not U14110 ( n13217,n11793 );
   nand U14111 ( n11793,n14149,n14150 );
   nand U14112 ( n14150,n11779,n11796 );
   not U14113 ( n11779,phyaddrpointer_reg_1_ );
   nand U14114 ( n14147,n14074,n10123 );
   nor U14115 ( n14145,n8803,n11796 );
   not U14116 ( n11796,phyaddrpointer_reg_2_ );
   nor U14117 ( n14143,n14151,n14152 );
   nor U14118 ( n14152,n10864,n14125 );
   nor U14119 ( n14151,n8802,n12649 );
   not U14120 ( n12649,eax_reg_2_ );
   nor U14121 ( n14141,n7819,n14153 );
   nor U14122 ( n14153,n9782,n8811 );
   not U14123 ( n9782,n8930 );
   nand U14124 ( n8930,n14154,n14155 );
   nand U14125 ( n14155,n14156,n14157 );
   nand U14126 ( n14157,n14158,n14159 );
   nand U14127 ( n14154,n14160,n14158 );
   nor U14128 ( n13251,n14161,n14162 );
   xor U14129 ( n14161,n14163,n8830 );
   nand U14130 ( n13252,n14162,n14163 );
   nand U14131 ( n14163,n14164,n14165 );
   nor U14132 ( n14165,n14166,n14167 );
   nand U14133 ( n14167,n14168,n14169 );
   nand U14134 ( n14169,n8830,n11814 );
   xor U14135 ( n11814,n11817,n14149 );
   nand U14136 ( n14168,n14074,n10466 );
   nor U14137 ( n14166,n8805,n11817 );
   nor U14138 ( n14164,n14170,n14171 );
   nor U14139 ( n14171,n14172,n14125 );
   nor U14140 ( n14170,n14040,n12654 );
   not U14141 ( n12654,eax_reg_3_ );
   nor U14142 ( n14162,n14090,n9781 );
   not U14143 ( n9781,n8944 );
   xor U14144 ( n8944,n14173,n14174 );
   nand U14145 ( n14174,n14175,n14176 );
   nor U14146 ( n14173,n14177,n14178 );
   nor U14147 ( n14177,n14179,n14180 );
   nand U14148 ( n13284,n14181,n14182 );
   nand U14149 ( n14182,n14074,n12409 );
   not U14150 ( n12409,n14183 );
   xor U14151 ( n14181,n14184,n8831 );
   nand U14152 ( n13285,n14185,n8784 );
   nor U14153 ( n14185,n14184,n14183 );
   xor U14154 ( n14183,n14186,n14187 );
   nand U14155 ( n14187,n14188,n14189 );
   and U14156 ( n14184,n14190,n14191 );
   nor U14157 ( n14191,n14192,n14193 );
   nand U14158 ( n14193,n14194,n14195 );
   nand U14159 ( n14195,n13297,n8829 );
   not U14160 ( n13297,n11835 );
   nand U14161 ( n11835,n14196,n14087 );
   nand U14162 ( n14196,n11838,n14197 );
   or U14163 ( n14197,n14149,n11817 );
   nand U14164 ( n14194,n14074,n10919 );
   xor U14165 ( n10919,n14091,n14088 );
   nand U14166 ( n14088,n14198,n14199 );
   nand U14167 ( n14091,instqueuerd_addr_reg_4_,n14200 );
   nand U14168 ( n14200,n9350,n10889 );
   nor U14169 ( n14192,n8804,n11838 );
   not U14170 ( n11838,phyaddrpointer_reg_4_ );
   nor U14171 ( n14190,n14201,n14202 );
   and U14172 ( n14202,instqueuerd_addr_reg_4_,n11710 );
   nor U14173 ( n14201,n8801,n12659 );
   not U14174 ( n12659,eax_reg_4_ );
   nand U14175 ( n13367,n14069,n13343 );
   or U14176 ( n13343,n14068,n14070 );
   nor U14177 ( n14070,n14090,n12422 );
   xor U14178 ( n12422,n14203,n14204 );
   nor U14179 ( n14203,n14205,n14206 );
   not U14180 ( n14206,n14207 );
   nand U14181 ( n14068,n14208,n14209 );
   nand U14182 ( n14209,n8829,n11865 );
   nand U14183 ( n11865,n14210,n14211 );
   nand U14184 ( n14210,n11868,n14212 );
   or U14185 ( n14212,n14087,n11853 );
   nor U14186 ( n14208,n14213,n14214 );
   nor U14187 ( n14214,n14040,n12669 );
   not U14188 ( n12669,eax_reg_6_ );
   nor U14189 ( n14213,n8805,n11868 );
   not U14190 ( n11868,phyaddrpointer_reg_6_ );
   not U14191 ( n14069,n13364 );
   nor U14192 ( n13364,n14063,n14062 );
   and U14193 ( n14062,n14215,n12426 );
   nor U14194 ( n12426,n14216,n14217 );
   and U14195 ( n14217,n14218,n14219 );
   nor U14196 ( n14219,n14205,n14082 );
   nor U14197 ( n14218,n14080,n14220 );
   and U14198 ( n14216,n14205,n14220 );
   nor U14199 ( n14215,n12427,n14090 );
   and U14200 ( n12427,n14221,n14204 );
   and U14201 ( n14221,n14207,n14220 );
   nand U14202 ( n14220,n14222,n14223 );
   xor U14203 ( n14063,n14224,n8765 );
   nor U14204 ( n14224,n14225,n14226 );
   nand U14205 ( n14226,n14227,n14228 );
   nand U14206 ( n14228,n8831,n11881 );
   xor U14207 ( n11881,n11884,n14211 );
   nand U14208 ( n14227,phyaddrpointer_reg_7_,n7819 );
   nor U14209 ( n14225,n8802,n12674 );
   not U14210 ( n12674,eax_reg_7_ );
   nand U14211 ( n13392,n14229,n14230 );
   nand U14212 ( n14230,n14074,n12361 );
   xor U14213 ( n14229,n8766,n14231 );
   nor U14214 ( n14054,n14232,n14233 );
   nor U14215 ( n14233,n14090,n14234 );
   nand U14216 ( n14234,n14235,n13458 );
   not U14217 ( n13458,n14059 );
   nand U14218 ( n14235,n14236,n14237 );
   nand U14219 ( n14237,n14238,n12441 );
   nand U14220 ( n14236,n12349,n14239 );
   nor U14221 ( n14232,n14240,n14241 );
   or U14222 ( n14241,n13461,n14059 );
   nor U14223 ( n14059,n14238,n14242 );
   and U14224 ( n14242,n14074,n12441 );
   xor U14225 ( n12441,n14243,n14244 );
   xor U14226 ( n14238,n14245,n8766 );
   nor U14227 ( n14245,n14246,n14247 );
   nand U14228 ( n14247,n14248,n14249 );
   nand U14229 ( n14249,n8829,n11956 );
   xor U14230 ( n11956,n11959,n14250 );
   nand U14231 ( n14248,phyaddrpointer_reg_11_,n7819 );
   nor U14232 ( n14246,n14040,n12692 );
   not U14233 ( n12692,eax_reg_11_ );
   nand U14234 ( n13461,n14074,n14251 );
   nand U14235 ( n14251,n14252,n14253 );
   nand U14236 ( n14253,n12361,n14231 );
   nand U14237 ( n14231,n14254,n14255 );
   nand U14238 ( n14255,eax_reg_8_,n13978 );
   nor U14239 ( n14254,n14256,n14257 );
   nor U14240 ( n14257,n8803,n11908 );
   nor U14241 ( n14256,n8763,n11905 );
   nand U14242 ( n11905,n14258,n14259 );
   nand U14243 ( n14259,n14260,n11908 );
   not U14244 ( n11908,phyaddrpointer_reg_8_ );
   or U14245 ( n14260,n14211,n11884 );
   xor U14246 ( n12361,n14261,n14262 );
   nand U14247 ( n14252,n12436,n14263 );
   not U14248 ( n12436,n12438 );
   nand U14249 ( n14240,n14058,n13460 );
   not U14250 ( n13460,n13412 );
   nor U14251 ( n13412,n14263,n14264 );
   nor U14252 ( n14264,n14090,n12438 );
   xor U14253 ( n12438,n14265,n14266 );
   nand U14254 ( n14266,n14261,n14262 );
   nand U14255 ( n14263,n14267,n14268 );
   nand U14256 ( n14268,n11920,n8830 );
   xor U14257 ( n11920,phyaddrpointer_reg_9_,n14258 );
   nor U14258 ( n14267,n14269,n14270 );
   nor U14259 ( n14270,n8801,n12683 );
   not U14260 ( n12683,eax_reg_9_ );
   nor U14261 ( n14269,n8804,n11923 );
   nand U14262 ( n14058,n14271,n14272 );
   nand U14263 ( n14272,n14074,n12349 );
   xor U14264 ( n12349,n14273,n14274 );
   xor U14265 ( n14271,n8764,n14239 );
   nand U14266 ( n14239,n14275,n14276 );
   nand U14267 ( n14276,eax_reg_10_,n13978 );
   nor U14268 ( n14275,n14277,n14278 );
   nor U14269 ( n14278,n8805,n11941 );
   nor U14270 ( n14277,n8763,n11938 );
   nand U14271 ( n11938,n14250,n14279 );
   nand U14272 ( n14279,n14280,n11941 );
   not U14273 ( n11941,phyaddrpointer_reg_10_ );
   or U14274 ( n14280,n14258,n11923 );
   not U14275 ( n14050,n13506 );
   nor U14276 ( n14043,n14281,n14282 );
   or U14277 ( n14282,n14283,n8811 );
   nand U14278 ( n14281,n12444,n13552 );
   nor U14279 ( n14041,n14284,n14285 );
   nor U14280 ( n14285,n14286,n14287 );
   nand U14281 ( n14287,n13558,n13552 );
   nand U14282 ( n13552,n14288,n14289 );
   nand U14283 ( n14289,n14074,n12448 );
   xor U14284 ( n14288,n14290,n8764 );
   nor U14285 ( n13558,n14053,n14052 );
   xor U14286 ( n14052,n14291,n8830 );
   nor U14287 ( n14291,n14292,n14293 );
   nand U14288 ( n14293,n14294,n14295 );
   nand U14289 ( n14295,n13485,n8831 );
   not U14290 ( n13485,n11976 );
   nand U14291 ( n11976,n14296,n14297 );
   nand U14292 ( n14296,n11979,n14298 );
   or U14293 ( n14298,n14250,n11959 );
   not U14294 ( n11979,phyaddrpointer_reg_12_ );
   nand U14295 ( n14294,phyaddrpointer_reg_12_,n7819 );
   nor U14296 ( n14292,n8802,n12697 );
   not U14297 ( n12697,eax_reg_12_ );
   nand U14298 ( n14053,n14074,n12344 );
   and U14299 ( n12344,n14299,n14300 );
   nand U14300 ( n14299,n14301,n14302 );
   nand U14301 ( n14302,n14244,n14243 );
   nand U14302 ( n14286,n13534,n13506 );
   nand U14303 ( n13506,n14049,n14048 );
   nand U14304 ( n14048,n14074,n12342 );
   xor U14305 ( n12342,n14303,n14304 );
   xor U14306 ( n14049,n14305,n8829 );
   nor U14307 ( n14305,n14306,n14307 );
   nand U14308 ( n14307,n14308,n14309 );
   nand U14309 ( n14309,n8830,n11991 );
   xor U14310 ( n11991,n11994,n14297 );
   nand U14311 ( n14308,phyaddrpointer_reg_13_,n7819 );
   nor U14312 ( n14306,n8802,n12702 );
   not U14313 ( n12702,eax_reg_13_ );
   nand U14314 ( n13534,n14283,n14310 );
   nand U14315 ( n14310,n14074,n12444 );
   not U14316 ( n12444,n12446 );
   nand U14317 ( n12446,n14311,n14312 );
   nand U14318 ( n14311,n14313,n14314 );
   nand U14319 ( n14314,n14303,n14304 );
   xor U14320 ( n14283,n8765,n14315 );
   nand U14321 ( n14315,n14316,n14317 );
   nand U14322 ( n14317,eax_reg_14_,n13978 );
   nor U14323 ( n14316,n14318,n14319 );
   nor U14324 ( n14319,n8803,n12009 );
   nor U14325 ( n14318,n8764,n12006 );
   nand U14326 ( n12006,n14320,n14321 );
   nand U14327 ( n14321,n14322,n12009 );
   not U14328 ( n12009,phyaddrpointer_reg_14_ );
   or U14329 ( n14322,n14297,n11994 );
   nor U14330 ( n14284,n14090,n14323 );
   nand U14331 ( n14323,n12448,n14290 );
   nand U14332 ( n14290,n14324,n14325 );
   nand U14333 ( n14325,eax_reg_15_,n13978 );
   not U14334 ( n13978,n8802 );
   nor U14335 ( n14324,n14326,n14327 );
   nor U14336 ( n14327,n8805,n12024 );
   nor U14337 ( n14326,n8765,n12021 );
   nand U14338 ( n12021,n14328,n14329 );
   nand U14339 ( n14329,n14320,n12024 );
   xor U14340 ( n12448,n14330,n14312 );
   nand U14341 ( n13588,n13938,n13937 );
   xor U14342 ( n13937,n8763,n14331 );
   nand U14343 ( n14331,n14332,n14333 );
   nor U14344 ( n14333,n14334,n14335 );
   nor U14345 ( n14335,n8764,n12036 );
   nand U14346 ( n12036,n14336,n14337 );
   nand U14347 ( n14336,n12039,n14328 );
   nor U14348 ( n14334,n14338,n13991 );
   nor U14349 ( n14338,n14339,n14340 );
   nand U14350 ( n14340,n14341,n14342 );
   nor U14351 ( n14342,n14343,n14344 );
   nand U14352 ( n14344,n14345,n14346 );
   nand U14353 ( n14346,n14000,instqueue_reg_7__0_ );
   nand U14354 ( n14345,n14001,instqueue_reg_6__0_ );
   nand U14355 ( n14343,n14347,n14348 );
   nand U14356 ( n14348,n14004,instqueue_reg_5__0_ );
   nand U14357 ( n14347,n14005,instqueue_reg_4__0_ );
   nor U14358 ( n14341,n14349,n14350 );
   nand U14359 ( n14350,n14351,n14352 );
   nand U14360 ( n14352,n14010,instqueue_reg_3__0_ );
   nand U14361 ( n14351,n14011,instqueue_reg_2__0_ );
   nand U14362 ( n14349,n14353,n14354 );
   nand U14363 ( n14354,n14014,instqueue_reg_1__0_ );
   nand U14364 ( n14353,n14015,instqueue_reg_0__0_ );
   nand U14365 ( n14339,n14355,n14356 );
   nor U14366 ( n14356,n14357,n14358 );
   nand U14367 ( n14358,n14359,n14360 );
   nand U14368 ( n14360,n14022,instqueue_reg_15__0_ );
   nand U14369 ( n14359,n14023,instqueue_reg_14__0_ );
   nand U14370 ( n14357,n14361,n14362 );
   nand U14371 ( n14362,n14026,instqueue_reg_13__0_ );
   nand U14372 ( n14361,n14027,instqueue_reg_12__0_ );
   nor U14373 ( n14355,n14363,n14364 );
   nand U14374 ( n14364,n14365,n14366 );
   nand U14375 ( n14366,n14032,instqueue_reg_11__0_ );
   nand U14376 ( n14365,n14033,instqueue_reg_10__0_ );
   nand U14377 ( n14363,n14367,n14368 );
   nand U14378 ( n14368,n14036,instqueue_reg_9__0_ );
   nand U14379 ( n14367,n14037,instqueue_reg_8__0_ );
   nor U14380 ( n14332,n14369,n14370 );
   nor U14381 ( n14370,n8801,n12715 );
   not U14382 ( n12715,eax_reg_16_ );
   nor U14383 ( n14369,n8805,n12039 );
   and U14384 ( n13938,n13943,n14371 );
   nand U14385 ( n14371,n14372,n8784 );
   and U14386 ( n14372,n8796,n12453 );
   nor U14387 ( n13933,n13608,n13635 );
   nor U14388 ( n13635,n13939,n13727 );
   xor U14389 ( n13939,n8829,n14374 );
   nand U14390 ( n14374,n14375,n14376 );
   nor U14391 ( n14376,n14377,n14378 );
   nor U14392 ( n14378,n8766,n12066 );
   nand U14393 ( n12066,n14379,n13989 );
   nand U14394 ( n14379,n12069,n14380 );
   nor U14395 ( n14377,n14381,n13991 );
   nor U14396 ( n14381,n14382,n14383 );
   nand U14397 ( n14383,n14384,n14385 );
   nor U14398 ( n14385,n14386,n14387 );
   nand U14399 ( n14387,n14388,n14389 );
   nand U14400 ( n14389,n14000,instqueue_reg_7__2_ );
   nand U14401 ( n14388,n14001,instqueue_reg_6__2_ );
   nand U14402 ( n14386,n14390,n14391 );
   nand U14403 ( n14391,n14004,instqueue_reg_5__2_ );
   nand U14404 ( n14390,n14005,instqueue_reg_4__2_ );
   nor U14405 ( n14384,n14392,n14393 );
   nand U14406 ( n14393,n14394,n14395 );
   nand U14407 ( n14395,n14010,instqueue_reg_3__2_ );
   nand U14408 ( n14394,n14011,instqueue_reg_2__2_ );
   nand U14409 ( n14392,n14396,n14397 );
   nand U14410 ( n14397,n14014,instqueue_reg_1__2_ );
   nand U14411 ( n14396,n14015,instqueue_reg_0__2_ );
   nand U14412 ( n14382,n14398,n14399 );
   nor U14413 ( n14399,n14400,n14401 );
   nand U14414 ( n14401,n14402,n14403 );
   nand U14415 ( n14403,n14022,instqueue_reg_15__2_ );
   nand U14416 ( n14402,n14023,instqueue_reg_14__2_ );
   nand U14417 ( n14400,n14404,n14405 );
   nand U14418 ( n14405,n14026,instqueue_reg_13__2_ );
   nand U14419 ( n14404,n14027,instqueue_reg_12__2_ );
   nor U14420 ( n14398,n14406,n14407 );
   nand U14421 ( n14407,n14408,n14409 );
   nand U14422 ( n14409,n14032,instqueue_reg_11__2_ );
   nand U14423 ( n14408,n14033,instqueue_reg_10__2_ );
   nand U14424 ( n14406,n14410,n14411 );
   nand U14425 ( n14411,n14036,instqueue_reg_9__2_ );
   nand U14426 ( n14410,n14037,instqueue_reg_8__2_ );
   nor U14427 ( n14375,n14412,n14413 );
   nor U14428 ( n14413,n8802,n12726 );
   not U14429 ( n12726,eax_reg_18_ );
   nor U14430 ( n14412,n8803,n12069 );
   not U14431 ( n13608,n13637 );
   nand U14432 ( n13637,n14414,n13943 );
   xor U14433 ( n14414,n13936,n8766 );
   nand U14434 ( n13936,n14415,n14416 );
   nor U14435 ( n14416,n14417,n14418 );
   nor U14436 ( n14418,n14419,n13991 );
   nor U14437 ( n14419,n14420,n14421 );
   nand U14438 ( n14421,n14422,n14423 );
   nor U14439 ( n14423,n14424,n14425 );
   nand U14440 ( n14425,n14426,n14427 );
   nand U14441 ( n14427,n14022,instqueue_reg_15__1_ );
   nand U14442 ( n14426,n14032,instqueue_reg_11__1_ );
   nand U14443 ( n14424,n14428,n14429 );
   nand U14444 ( n14429,n14000,instqueue_reg_7__1_ );
   nand U14445 ( n14428,n14010,instqueue_reg_3__1_ );
   nor U14446 ( n14422,n14430,n14431 );
   nand U14447 ( n14431,n14432,n14433 );
   nand U14448 ( n14433,n14036,instqueue_reg_9__1_ );
   nand U14449 ( n14432,n14037,instqueue_reg_8__1_ );
   nand U14450 ( n14430,n14434,n14435 );
   nand U14451 ( n14435,n14027,instqueue_reg_12__1_ );
   nand U14452 ( n14434,n14033,instqueue_reg_10__1_ );
   nand U14453 ( n14420,n14436,n14437 );
   nor U14454 ( n14437,n14438,n14439 );
   nand U14455 ( n14439,n14440,n14441 );
   nand U14456 ( n14441,n14026,instqueue_reg_13__1_ );
   nand U14457 ( n14440,n14023,instqueue_reg_14__1_ );
   nand U14458 ( n14438,n14442,n14443 );
   nand U14459 ( n14443,n14014,instqueue_reg_1__1_ );
   nand U14460 ( n14442,n14015,instqueue_reg_0__1_ );
   nor U14461 ( n14436,n14444,n14445 );
   nand U14462 ( n14445,n14446,n14447 );
   nand U14463 ( n14447,n14005,instqueue_reg_4__1_ );
   nand U14464 ( n14446,n14011,instqueue_reg_2__1_ );
   nand U14465 ( n14444,n14448,n14449 );
   nand U14466 ( n14449,n14004,instqueue_reg_5__1_ );
   nand U14467 ( n14448,n14001,instqueue_reg_6__1_ );
   nor U14468 ( n14417,n8763,n12052 );
   nand U14469 ( n12052,n14380,n14450 );
   nand U14470 ( n14450,n14337,n12055 );
   nor U14471 ( n14415,n14451,n14452 );
   nor U14472 ( n14452,n14040,n12721 );
   not U14473 ( n12721,eax_reg_17_ );
   nor U14474 ( n14451,n8804,n12055 );
   nor U14475 ( n13983,n13925,n13874 );
   nand U14476 ( n13874,n13821,n13846 );
   nand U14477 ( n13846,n14453,n13943 );
   xor U14478 ( n14453,n13951,n8831 );
   and U14479 ( n13951,n14454,n14455 );
   nor U14480 ( n14455,n14456,n14457 );
   nor U14481 ( n14457,n8801,n12771 );
   not U14482 ( n12771,eax_reg_27_ );
   nor U14483 ( n14456,n8764,n12239 );
   nand U14484 ( n12239,n14458,n14459 );
   nand U14485 ( n14459,n14460,n12242 );
   nor U14486 ( n14454,n14461,n14462 );
   xor U14487 ( n14462,n14463,n14464 );
   nor U14488 ( n14461,n8804,n12242 );
   nand U14489 ( n13821,n13954,n13943 );
   xor U14490 ( n13954,n8765,n14465 );
   nand U14491 ( n14465,n14466,n14467 );
   nor U14492 ( n14467,n14468,n14469 );
   nor U14493 ( n14469,n8766,n12223 );
   nand U14494 ( n12223,n14470,n14460 );
   nand U14495 ( n14470,n12226,n14471 );
   nor U14496 ( n14468,n14472,n14473 );
   nor U14497 ( n14473,n14474,n14475 );
   not U14498 ( n14472,n14464 );
   nor U14499 ( n14466,n14476,n14477 );
   nor U14500 ( n14477,n8801,n12766 );
   not U14501 ( n12766,eax_reg_26_ );
   nor U14502 ( n14476,n8805,n12226 );
   nand U14503 ( n13925,n14478,n14479 );
   nor U14504 ( n14479,n13723,n14480 );
   nand U14505 ( n14480,n13777,n13679 );
   not U14506 ( n13679,n13776 );
   nor U14507 ( n13776,n13726,n13727 );
   xor U14508 ( n13726,n8829,n14481 );
   nand U14509 ( n14481,n14482,n14483 );
   nor U14510 ( n14483,n14484,n14485 );
   nor U14511 ( n14485,n8763,n12103 );
   nand U14512 ( n12103,n14486,n14487 );
   nand U14513 ( n14486,n12106,n14488 );
   nand U14514 ( n14488,n14489,phyaddrpointer_reg_19_ );
   nor U14515 ( n14484,n14490,n13991 );
   nor U14516 ( n14490,n14491,n14492 );
   nand U14517 ( n14492,n14493,n14494 );
   nor U14518 ( n14494,n14495,n14496 );
   nand U14519 ( n14496,n14497,n14498 );
   nand U14520 ( n14498,n14000,instqueue_reg_7__4_ );
   nand U14521 ( n14497,n14001,instqueue_reg_6__4_ );
   nand U14522 ( n14495,n14499,n14500 );
   nand U14523 ( n14500,n14004,instqueue_reg_5__4_ );
   nand U14524 ( n14499,n14005,instqueue_reg_4__4_ );
   nor U14525 ( n14493,n14501,n14502 );
   nand U14526 ( n14502,n14503,n14504 );
   nand U14527 ( n14504,n14010,instqueue_reg_3__4_ );
   nand U14528 ( n14503,n14011,instqueue_reg_2__4_ );
   nand U14529 ( n14501,n14505,n14506 );
   nand U14530 ( n14506,n14014,instqueue_reg_1__4_ );
   nand U14531 ( n14505,n14015,instqueue_reg_0__4_ );
   nand U14532 ( n14491,n14507,n14508 );
   nor U14533 ( n14508,n14509,n14510 );
   nand U14534 ( n14510,n14511,n14512 );
   nand U14535 ( n14512,n14022,instqueue_reg_15__4_ );
   nand U14536 ( n14511,n14023,instqueue_reg_14__4_ );
   nand U14537 ( n14509,n14513,n14514 );
   nand U14538 ( n14514,n14026,instqueue_reg_13__4_ );
   nand U14539 ( n14513,n14027,instqueue_reg_12__4_ );
   nor U14540 ( n14507,n14515,n14516 );
   nand U14541 ( n14516,n14517,n14518 );
   nand U14542 ( n14518,n14032,instqueue_reg_11__4_ );
   nand U14543 ( n14517,n14033,instqueue_reg_10__4_ );
   nand U14544 ( n14515,n14519,n14520 );
   nand U14545 ( n14520,n14036,instqueue_reg_9__4_ );
   nand U14546 ( n14519,n14037,instqueue_reg_8__4_ );
   nor U14547 ( n14482,n14521,n14522 );
   nor U14548 ( n14522,n14040,n12736 );
   not U14549 ( n12736,eax_reg_20_ );
   nor U14550 ( n14521,n8805,n12106 );
   not U14551 ( n12106,phyaddrpointer_reg_20_ );
   nand U14552 ( n13777,n14523,n13943 );
   xor U14553 ( n14523,n13949,n8763 );
   nand U14554 ( n13949,n14524,n14525 );
   nor U14555 ( n14525,n14526,n14527 );
   nor U14556 ( n14527,n8802,n12741 );
   not U14557 ( n12741,eax_reg_21_ );
   nor U14558 ( n14526,n12120,n8763 );
   xor U14559 ( n12120,phyaddrpointer_reg_21_,n14487 );
   nor U14560 ( n14524,n14528,n14529 );
   nor U14561 ( n14529,n8805,n12123 );
   nor U14562 ( n14528,n14530,n13991 );
   nor U14563 ( n14530,n14531,n14532 );
   nand U14564 ( n14532,n14533,n14534 );
   nor U14565 ( n14534,n14535,n14536 );
   nand U14566 ( n14536,n14537,n14538 );
   nand U14567 ( n14538,n14022,instqueue_reg_15__5_ );
   nand U14568 ( n14537,n14032,instqueue_reg_11__5_ );
   nand U14569 ( n14535,n14539,n14540 );
   nand U14570 ( n14540,n14000,instqueue_reg_7__5_ );
   nand U14571 ( n14539,n14010,instqueue_reg_3__5_ );
   nor U14572 ( n14533,n14541,n14542 );
   nand U14573 ( n14542,n14543,n14544 );
   nand U14574 ( n14544,n14036,instqueue_reg_9__5_ );
   nand U14575 ( n14543,n14037,instqueue_reg_8__5_ );
   nand U14576 ( n14541,n14545,n14546 );
   nand U14577 ( n14546,n14027,instqueue_reg_12__5_ );
   nand U14578 ( n14545,n14033,instqueue_reg_10__5_ );
   nand U14579 ( n14531,n14547,n14548 );
   nor U14580 ( n14548,n14549,n14550 );
   nand U14581 ( n14550,n14551,n14552 );
   nand U14582 ( n14552,n14026,instqueue_reg_13__5_ );
   nand U14583 ( n14551,n14023,instqueue_reg_14__5_ );
   nand U14584 ( n14549,n14553,n14554 );
   nand U14585 ( n14554,n14014,instqueue_reg_1__5_ );
   nand U14586 ( n14553,n14015,instqueue_reg_0__5_ );
   nor U14587 ( n14547,n14555,n14556 );
   nand U14588 ( n14556,n14557,n14558 );
   nand U14589 ( n14558,n14005,instqueue_reg_4__5_ );
   nand U14590 ( n14557,n14011,instqueue_reg_2__5_ );
   nand U14591 ( n14555,n14559,n14560 );
   nand U14592 ( n14560,n14004,instqueue_reg_5__5_ );
   nand U14593 ( n14559,n14001,instqueue_reg_6__5_ );
   and U14594 ( n13723,n14561,n13943 );
   xor U14595 ( n14561,n13948,n8830 );
   and U14596 ( n13948,n14562,n14563 );
   nor U14597 ( n14563,n14564,n14565 );
   nor U14598 ( n14565,n8802,n12746 );
   not U14599 ( n12746,eax_reg_22_ );
   nor U14600 ( n14564,n8764,n12141 );
   nand U14601 ( n12141,n14566,n14567 );
   nand U14602 ( n14567,n14568,n12144 );
   or U14603 ( n14568,n14487,n12123 );
   nor U14604 ( n14562,n14569,n14570 );
   nor U14605 ( n14570,n8804,n12144 );
   not U14606 ( n12144,phyaddrpointer_reg_22_ );
   nor U14607 ( n14569,n14571,n13991 );
   nand U14608 ( n13991,n14074,n14572 );
   nor U14609 ( n14571,n14573,n14574 );
   nand U14610 ( n14574,n14575,n14576 );
   nor U14611 ( n14576,n14577,n14578 );
   nand U14612 ( n14578,n14579,n14580 );
   nand U14613 ( n14580,n14022,instqueue_reg_15__6_ );
   not U14614 ( n14022,n14581 );
   nand U14615 ( n14579,n14032,instqueue_reg_11__6_ );
   not U14616 ( n14032,n14582 );
   nand U14617 ( n14577,n14583,n14584 );
   nand U14618 ( n14584,n14000,instqueue_reg_7__6_ );
   not U14619 ( n14000,n14585 );
   nand U14620 ( n14583,n14010,instqueue_reg_3__6_ );
   not U14621 ( n14010,n14586 );
   nor U14622 ( n14575,n14587,n14588 );
   nand U14623 ( n14588,n14589,n14590 );
   nand U14624 ( n14590,n14036,instqueue_reg_9__6_ );
   not U14625 ( n14036,n14591 );
   nand U14626 ( n14589,n14037,instqueue_reg_8__6_ );
   not U14627 ( n14037,n14592 );
   nand U14628 ( n14587,n14593,n14594 );
   nand U14629 ( n14594,n14027,instqueue_reg_12__6_ );
   not U14630 ( n14027,n14595 );
   nand U14631 ( n14593,n14033,instqueue_reg_10__6_ );
   not U14632 ( n14033,n14596 );
   nand U14633 ( n14573,n14597,n14598 );
   nor U14634 ( n14598,n14599,n14600 );
   nand U14635 ( n14600,n14601,n14602 );
   nand U14636 ( n14602,n14026,instqueue_reg_13__6_ );
   not U14637 ( n14026,n14603 );
   nand U14638 ( n14601,n14023,instqueue_reg_14__6_ );
   not U14639 ( n14023,n14604 );
   nand U14640 ( n14599,n14605,n14606 );
   nand U14641 ( n14606,n14014,instqueue_reg_1__6_ );
   not U14642 ( n14014,n14607 );
   nand U14643 ( n14605,n14015,instqueue_reg_0__6_ );
   not U14644 ( n14015,n14608 );
   nor U14645 ( n14597,n14609,n14610 );
   nand U14646 ( n14610,n14611,n14612 );
   nand U14647 ( n14612,n14005,instqueue_reg_4__6_ );
   not U14648 ( n14005,n14613 );
   nand U14649 ( n14611,n14011,instqueue_reg_2__6_ );
   not U14650 ( n14011,n14614 );
   nand U14651 ( n14609,n14615,n14616 );
   nand U14652 ( n14616,n14004,instqueue_reg_5__6_ );
   not U14653 ( n14004,n14617 );
   nand U14654 ( n14615,n14001,instqueue_reg_6__6_ );
   not U14655 ( n14001,n14618 );
   nor U14656 ( n14478,n13748,n13769 );
   nor U14657 ( n13769,n13945,n13727 );
   xor U14658 ( n13945,n8830,n14619 );
   nand U14659 ( n14619,n14620,n14621 );
   nor U14660 ( n14621,n14622,n14623 );
   nor U14661 ( n14623,n8766,n12176 );
   nand U14662 ( n12176,n14624,n14625 );
   nand U14663 ( n14624,n12179,n14626 );
   nor U14664 ( n14622,n14090,n14627 );
   nand U14665 ( n14627,n14628,n14629 );
   nand U14666 ( n14628,n14630,n14631 );
   nand U14667 ( n14631,n14632,n14572 );
   or U14668 ( n14630,n14633,n14634 );
   nor U14669 ( n14620,n14635,n14636 );
   nor U14670 ( n14636,n8801,n12756 );
   not U14671 ( n12756,eax_reg_24_ );
   nor U14672 ( n14635,n8803,n12179 );
   nor U14673 ( n13748,n13944,n13727 );
   not U14674 ( n13727,n13943 );
   xor U14675 ( n13944,n8829,n14637 );
   nand U14676 ( n14637,n14638,n14639 );
   nor U14677 ( n14639,n14640,n14641 );
   nor U14678 ( n14641,n8765,n12159 );
   nand U14679 ( n12159,n14626,n14642 );
   nand U14680 ( n14642,n14566,n12162 );
   nor U14681 ( n14640,n14643,n8811 );
   xor U14682 ( n14643,n14634,n14644 );
   nor U14683 ( n14638,n14645,n14646 );
   nor U14684 ( n14646,n14040,n12751 );
   not U14685 ( n12751,eax_reg_23_ );
   nor U14686 ( n14645,n8804,n12162 );
   nand U14687 ( n13981,n13922,n14647 );
   and U14688 ( n14647,n13918,n13799 );
   nand U14689 ( n13799,n14648,n13943 );
   xor U14690 ( n14648,n13955,n8765 );
   nand U14691 ( n13955,n14649,n14650 );
   nor U14692 ( n14650,n14651,n14652 );
   nor U14693 ( n14652,n8766,n12204 );
   nand U14694 ( n12204,n14471,n14653 );
   nand U14695 ( n14653,n14625,n12207 );
   and U14696 ( n14651,n14654,n8784 );
   xor U14697 ( n14654,n14655,n14629 );
   nor U14698 ( n14649,n14656,n14657 );
   nor U14699 ( n14657,n8802,n12761 );
   not U14700 ( n12761,eax_reg_25_ );
   nor U14701 ( n14656,n8804,n12207 );
   nand U14702 ( n13918,n14658,n13943 );
   xor U14703 ( n14658,n14659,n8763 );
   nand U14704 ( n14659,n14660,n14661 );
   nor U14705 ( n14661,n14662,n14663 );
   nand U14706 ( n14663,n14664,n14665 );
   nand U14707 ( n14665,n14666,n14667 );
   nor U14708 ( n14666,n14668,n14669 );
   nand U14709 ( n14664,n14670,n14671 );
   or U14710 ( n14671,n14669,n14668 );
   not U14711 ( n14670,n14667 );
   nand U14712 ( n14667,n14572,n14672 );
   nand U14713 ( n14672,n14673,n14674 );
   nor U14714 ( n14674,n14675,n14676 );
   nand U14715 ( n14676,n14677,n14678 );
   nor U14716 ( n14678,n14679,n14680 );
   nor U14717 ( n14680,n14681,n14682 );
   nor U14718 ( n14679,n14683,n14684 );
   nor U14719 ( n14677,n14685,n14686 );
   nor U14720 ( n14686,n14687,n14688 );
   nor U14721 ( n14685,n10750,n14689 );
   nand U14722 ( n14675,n14690,n14691 );
   nor U14723 ( n14691,n14692,n14693 );
   nor U14724 ( n14693,n14694,n14695 );
   nor U14725 ( n14692,n14696,n14697 );
   nor U14726 ( n14690,n14698,n14699 );
   nor U14727 ( n14699,n14700,n14701 );
   nor U14728 ( n14698,n14702,n14703 );
   nor U14729 ( n14673,n14704,n14705 );
   nand U14730 ( n14705,n14706,n14707 );
   nor U14731 ( n14707,n14708,n14709 );
   nor U14732 ( n14709,n14710,n14711 );
   nor U14733 ( n14708,n14712,n14713 );
   nor U14734 ( n14706,n14714,n14715 );
   nor U14735 ( n14715,n14716,n14717 );
   nor U14736 ( n14714,n14718,n14719 );
   nand U14737 ( n14704,n14720,n14721 );
   nor U14738 ( n14721,n14722,n14723 );
   nor U14739 ( n14723,n14724,n14725 );
   nor U14740 ( n14722,n14726,n14727 );
   nor U14741 ( n14720,n14728,n14729 );
   nor U14742 ( n14729,n14730,n14731 );
   nor U14743 ( n14728,n14732,n14733 );
   nor U14744 ( n14662,n8765,n12298 );
   nand U14745 ( n12298,n14734,n14735 );
   or U14746 ( n14735,n14736,phyaddrpointer_reg_30_ );
   nor U14747 ( n14660,n14737,n14738 );
   nor U14748 ( n14738,n8801,n12786 );
   not U14749 ( n12786,eax_reg_30_ );
   nor U14750 ( n14737,n8803,n12301 );
   not U14751 ( n12301,phyaddrpointer_reg_30_ );
   nor U14752 ( n13922,n13869,n13897 );
   and U14753 ( n13897,n14739,n13943 );
   xor U14754 ( n14739,n14740,n8764 );
   nand U14755 ( n14740,n14741,n14742 );
   nor U14756 ( n14742,n14743,n14744 );
   nor U14757 ( n14744,n8803,n12282 );
   nor U14758 ( n14743,n12279,n8764 );
   xor U14759 ( n12279,phyaddrpointer_reg_29_,n14745 );
   nor U14760 ( n14741,n14746,n14747 );
   xor U14761 ( n14747,n14669,n14668 );
   nand U14762 ( n14669,n14572,n14748 );
   nand U14763 ( n14748,n14749,n14750 );
   nor U14764 ( n14750,n14751,n14752 );
   nand U14765 ( n14752,n14753,n14754 );
   nor U14766 ( n14754,n14755,n14756 );
   nor U14767 ( n14756,n14757,n14682 );
   nor U14768 ( n14755,n14758,n14684 );
   nor U14769 ( n14753,n14759,n14760 );
   nor U14770 ( n14760,n14761,n14688 );
   nor U14771 ( n14759,n10761,n14689 );
   nand U14772 ( n14751,n14762,n14763 );
   nor U14773 ( n14763,n14764,n14765 );
   nor U14774 ( n14765,n14766,n14695 );
   nor U14775 ( n14764,n14767,n14697 );
   nor U14776 ( n14762,n14768,n14769 );
   nor U14777 ( n14769,n14770,n14701 );
   nor U14778 ( n14768,n14771,n14703 );
   nor U14779 ( n14749,n14772,n14773 );
   nand U14780 ( n14773,n14774,n14775 );
   nor U14781 ( n14775,n14776,n14777 );
   nor U14782 ( n14777,n14778,n14711 );
   nor U14783 ( n14776,n14779,n14713 );
   nor U14784 ( n14774,n14780,n14781 );
   nor U14785 ( n14781,n14782,n14717 );
   nor U14786 ( n14780,n14783,n14719 );
   nand U14787 ( n14772,n14784,n14785 );
   nor U14788 ( n14785,n14786,n14787 );
   nor U14789 ( n14787,n14788,n14725 );
   nor U14790 ( n14786,n14789,n14727 );
   nor U14791 ( n14784,n14790,n14791 );
   nor U14792 ( n14791,n14792,n14731 );
   nor U14793 ( n14790,n14793,n14733 );
   nor U14794 ( n14746,n14040,n12781 );
   not U14795 ( n12781,eax_reg_29_ );
   and U14796 ( n13869,n13952,n13943 );
   nand U14797 ( n13943,n14794,n8784 );
   not U14798 ( n14074,n14090 );
   nand U14799 ( n14090,state2_reg_2_,n14795 );
   nand U14800 ( n14795,n10906,n10758 );
   nor U14801 ( n14794,n12453,n8796 );
   nor U14802 ( n12453,n14312,n14330 );
   and U14803 ( n14330,n14796,n14797 );
   nor U14804 ( n14796,n14798,n14799 );
   nor U14805 ( n14799,n8796,n14800 );
   nor U14806 ( n14798,n14801,n14802 );
   not U14807 ( n14801,n14800 );
   nand U14808 ( n14800,n14803,n14804 );
   nor U14809 ( n14804,n14805,n14806 );
   nand U14810 ( n14806,n14807,n14808 );
   nor U14811 ( n14808,n14809,n14810 );
   nor U14812 ( n14810,n14716,n14811 );
   nor U14813 ( n14809,n14718,n14812 );
   nor U14814 ( n14807,n14813,n14814 );
   nor U14815 ( n14814,n14710,n14815 );
   nor U14816 ( n14813,n14712,n14816 );
   nand U14817 ( n14805,n14817,n14818 );
   nor U14818 ( n14818,n14819,n14820 );
   nor U14819 ( n14820,n14730,n14821 );
   nor U14820 ( n14819,n14732,n14822 );
   nor U14821 ( n14817,n14823,n14824 );
   nor U14822 ( n14824,n14724,n14825 );
   nor U14823 ( n14823,n14726,n14826 );
   nor U14824 ( n14803,n14827,n14828 );
   nand U14825 ( n14828,n14829,n14830 );
   nor U14826 ( n14830,n14831,n14832 );
   nor U14827 ( n14832,n14683,n14833 );
   nor U14828 ( n14831,n14687,n14834 );
   nor U14829 ( n14829,n14835,n14836 );
   nor U14830 ( n14836,n14702,n14837 );
   nor U14831 ( n14835,n14681,n14838 );
   nand U14832 ( n14827,n14839,n14840 );
   nor U14833 ( n14840,n14841,n14842 );
   nor U14834 ( n14842,n14696,n14843 );
   nor U14835 ( n14841,n14700,n14844 );
   nor U14836 ( n14839,n14845,n14846 );
   nor U14837 ( n14846,n10750,n14847 );
   nor U14838 ( n14845,n14694,n14848 );
   nand U14839 ( n14312,n14849,n14303 );
   not U14840 ( n14303,n14300 );
   nand U14841 ( n14300,n14850,n14244 );
   and U14842 ( n14244,n14273,n14274 );
   nand U14843 ( n14274,n14851,n14797 );
   nor U14844 ( n14851,n14852,n14853 );
   nor U14845 ( n14853,n8796,n14854 );
   nor U14846 ( n14852,n14855,n14802 );
   not U14847 ( n14855,n14854 );
   nand U14848 ( n14854,n14856,n14857 );
   nor U14849 ( n14857,n14858,n14859 );
   nand U14850 ( n14859,n14860,n14861 );
   nor U14851 ( n14861,n14862,n14863 );
   nor U14852 ( n14863,n14864,n14811 );
   nor U14853 ( n14862,n14865,n14812 );
   nor U14854 ( n14860,n14866,n14867 );
   nor U14855 ( n14867,n14868,n14815 );
   nor U14856 ( n14866,n14869,n14816 );
   nand U14857 ( n14858,n14870,n14871 );
   nor U14858 ( n14871,n14872,n14873 );
   nor U14859 ( n14873,n14874,n14821 );
   nor U14860 ( n14872,n14875,n14822 );
   nor U14861 ( n14870,n14876,n14877 );
   nor U14862 ( n14877,n14878,n14825 );
   nor U14863 ( n14876,n14879,n14826 );
   nor U14864 ( n14856,n14880,n14881 );
   nand U14865 ( n14881,n14882,n14883 );
   nor U14866 ( n14883,n14884,n14885 );
   nor U14867 ( n14885,n14886,n14833 );
   nor U14868 ( n14884,n14887,n14834 );
   nor U14869 ( n14882,n14888,n14889 );
   nor U14870 ( n14889,n14890,n14837 );
   nor U14871 ( n14888,n14891,n14838 );
   nand U14872 ( n14880,n14892,n14893 );
   nor U14873 ( n14893,n14894,n14895 );
   nor U14874 ( n14895,n14896,n14843 );
   nor U14875 ( n14894,n14897,n14844 );
   nor U14876 ( n14892,n14898,n14899 );
   nor U14877 ( n14899,n10801,n14847 );
   nor U14878 ( n14898,n14900,n14848 );
   and U14879 ( n14273,n14901,n14265 );
   nand U14880 ( n14265,n14902,n14797 );
   nor U14881 ( n14902,n14903,n14904 );
   nor U14882 ( n14904,n8796,n14905 );
   nor U14883 ( n14903,n14906,n14802 );
   not U14884 ( n14906,n14905 );
   nand U14885 ( n14905,n14907,n14908 );
   nor U14886 ( n14908,n14909,n14910 );
   nand U14887 ( n14910,n14911,n14912 );
   nor U14888 ( n14912,n14913,n14914 );
   nor U14889 ( n14914,n14915,n14811 );
   nor U14890 ( n14913,n14916,n14812 );
   nor U14891 ( n14911,n14917,n14918 );
   nor U14892 ( n14918,n14919,n14815 );
   nor U14893 ( n14917,n14920,n14816 );
   nand U14894 ( n14909,n14921,n14922 );
   nor U14895 ( n14922,n14923,n14924 );
   nor U14896 ( n14924,n14925,n14821 );
   nor U14897 ( n14923,n14926,n14822 );
   nor U14898 ( n14921,n14927,n14928 );
   nor U14899 ( n14928,n14929,n14825 );
   nor U14900 ( n14927,n14930,n14826 );
   nor U14901 ( n14907,n14931,n14932 );
   nand U14902 ( n14932,n14933,n14934 );
   nor U14903 ( n14934,n14935,n14936 );
   nor U14904 ( n14936,n14937,n14833 );
   nor U14905 ( n14935,n14938,n14834 );
   nor U14906 ( n14933,n14939,n14940 );
   nor U14907 ( n14940,n14941,n14837 );
   nor U14908 ( n14939,n14942,n14838 );
   nand U14909 ( n14931,n14943,n14944 );
   nor U14910 ( n14944,n14945,n14946 );
   nor U14911 ( n14946,n14947,n14843 );
   nor U14912 ( n14945,n14948,n14844 );
   nor U14913 ( n14943,n14949,n14950 );
   nor U14914 ( n14950,n10811,n14847 );
   nor U14915 ( n14949,n14951,n14848 );
   and U14916 ( n14901,n14261,n14262 );
   nand U14917 ( n14262,n14223,n14952 );
   nand U14918 ( n14952,n14953,n14222 );
   or U14919 ( n14222,n14954,n12454 );
   nand U14920 ( n14953,n14207,n14955 );
   or U14921 ( n14955,n14204,n14205 );
   nor U14922 ( n14205,n14956,n14957 );
   nor U14923 ( n14204,n14081,n14958 );
   nor U14924 ( n14958,n14080,n14082 );
   and U14925 ( n14082,n14959,n14960 );
   and U14926 ( n14080,n14189,n14961 );
   nand U14927 ( n14961,n14186,n14188 );
   or U14928 ( n14188,n14962,n14963 );
   nand U14929 ( n14186,n14175,n14964 );
   nand U14930 ( n14964,n14965,n14176 );
   nand U14931 ( n14176,n14966,n14967 );
   nor U14932 ( n14965,n14179,n14160 );
   nor U14933 ( n14160,n14156,n14178 );
   not U14934 ( n14178,n14159 );
   nand U14935 ( n14159,n14968,n14969 );
   or U14936 ( n14969,n14970,n12454 );
   nor U14937 ( n14968,n14971,n12397 );
   not U14938 ( n14156,n14180 );
   nand U14939 ( n14180,n14140,n14972 );
   nand U14940 ( n14972,n14110,n14139 );
   or U14941 ( n14139,n14973,n14974 );
   nor U14942 ( n14110,n14109,n12454 );
   and U14943 ( n14109,n14975,n14976 );
   or U14944 ( n14976,n14116,n8821 );
   nand U14945 ( n14116,n14977,n14978 );
   nand U14946 ( n14978,n14979,n12382 );
   nand U14947 ( n14977,n11708,n12430 );
   xor U14948 ( n14975,n14115,n12454 );
   nand U14949 ( n14115,n14980,n14981 );
   nand U14950 ( n14981,n9348,n8821 );
   not U14951 ( n9348,n8910 );
   nand U14952 ( n8910,n14982,n14983 );
   nand U14953 ( n14983,n14984,n14985 );
   nor U14954 ( n14980,n14986,n14987 );
   nor U14955 ( n14987,n12382,n8796 );
   and U14956 ( n14986,n12382,n14988 );
   nand U14957 ( n12382,n14989,n14990 );
   nor U14958 ( n14990,n14991,n14992 );
   nand U14959 ( n14992,n14993,n14994 );
   nor U14960 ( n14994,n14995,n14996 );
   nor U14961 ( n14996,n14997,n14998 );
   nor U14962 ( n14995,n14999,n15000 );
   nor U14963 ( n14993,n15001,n15002 );
   nor U14964 ( n15002,n15003,n15004 );
   nor U14965 ( n15001,n15005,n15006 );
   nand U14966 ( n14991,n15007,n15008 );
   nor U14967 ( n15008,n15009,n15010 );
   nor U14968 ( n15010,n15011,n15012 );
   nor U14969 ( n15009,n15013,n15014 );
   nor U14970 ( n15007,n15015,n15016 );
   nor U14971 ( n15016,n15017,n15018 );
   nor U14972 ( n15015,n15019,n15020 );
   nor U14973 ( n14989,n15021,n15022 );
   nand U14974 ( n15022,n15023,n15024 );
   nor U14975 ( n15024,n15025,n15026 );
   nor U14976 ( n15026,n15027,n15028 );
   nor U14977 ( n15025,n15029,n15030 );
   nor U14978 ( n15023,n15031,n15032 );
   nor U14979 ( n15032,n15033,n15034 );
   nor U14980 ( n15031,n15035,n15036 );
   nand U14981 ( n15021,n15037,n15038 );
   nor U14982 ( n15038,n15039,n15040 );
   nor U14983 ( n15040,n10825,n15041 );
   nor U14984 ( n15039,n15042,n15043 );
   nor U14985 ( n15037,n15044,n15045 );
   nor U14986 ( n15045,n15046,n15047 );
   nor U14987 ( n15044,n15048,n15049 );
   nand U14988 ( n14140,n14974,n14973 );
   xor U14989 ( n14973,n14373,n15050 );
   nand U14990 ( n15050,n15051,n15052 );
   nand U14991 ( n15052,n9603,n8821 );
   not U14992 ( n9603,n8920 );
   xor U14993 ( n8920,n15053,n15054 );
   xor U14994 ( n15053,n15055,n14982 );
   nor U14995 ( n15051,n15056,n15057 );
   nor U14996 ( n15057,n8796,n12433 );
   nor U14997 ( n15056,n12389,n15058 );
   and U14998 ( n14974,n15059,n15060 );
   nand U14999 ( n15060,n15061,instqueue_reg_0__1_ );
   nor U15000 ( n15059,n14988,n15062 );
   nor U15001 ( n15062,n12389,n15063 );
   not U15002 ( n12389,n12433 );
   nand U15003 ( n12433,n15064,n15065 );
   nor U15004 ( n15065,n15066,n15067 );
   nand U15005 ( n15067,n15068,n15069 );
   nor U15006 ( n15069,n15070,n15071 );
   nor U15007 ( n15071,n14951,n14998 );
   nor U15008 ( n15070,n14947,n15000 );
   nor U15009 ( n15068,n15072,n15073 );
   nor U15010 ( n15073,n14948,n15004 );
   nor U15011 ( n15072,n14942,n15006 );
   nand U15012 ( n15066,n15074,n15075 );
   nor U15013 ( n15075,n15076,n15077 );
   nor U15014 ( n15077,n14937,n15012 );
   nor U15015 ( n15076,n14938,n15014 );
   nor U15016 ( n15074,n15078,n15079 );
   nor U15017 ( n15079,n14930,n15018 );
   nor U15018 ( n15078,n14925,n15020 );
   nor U15019 ( n15064,n15080,n15081 );
   nand U15020 ( n15081,n15082,n15083 );
   nor U15021 ( n15083,n15084,n15085 );
   nor U15022 ( n15085,n14926,n15028 );
   nor U15023 ( n15084,n14920,n15030 );
   nor U15024 ( n15082,n15086,n15087 );
   nor U15025 ( n15087,n14915,n15034 );
   nor U15026 ( n15086,n14916,n15036 );
   nand U15027 ( n15080,n15088,n15089 );
   nor U15028 ( n15089,n15090,n15091 );
   nor U15029 ( n15091,n10811,n15041 );
   nor U15030 ( n15090,n14941,n15043 );
   nor U15031 ( n15088,n15092,n15093 );
   nor U15032 ( n15093,n14929,n15047 );
   nor U15033 ( n15092,n14919,n15049 );
   not U15034 ( n14988,n15058 );
   not U15035 ( n14179,n14158 );
   nand U15036 ( n14158,n15094,n15095 );
   xor U15037 ( n15095,n14970,n14373 );
   nand U15038 ( n14970,n15096,n15097 );
   nand U15039 ( n15097,n10123,n8821 );
   not U15040 ( n10123,n8933 );
   xor U15041 ( n8933,n15098,n15099 );
   nor U15042 ( n15098,n15100,n15101 );
   nor U15043 ( n15096,n15102,n15103 );
   nor U15044 ( n15103,n8796,n15104 );
   nor U15045 ( n15102,n12397,n15058 );
   nor U15046 ( n15094,n15105,n15106 );
   nor U15047 ( n15106,n11732,n10801 );
   nor U15048 ( n15105,n12397,n15063 );
   not U15049 ( n12397,n15104 );
   nand U15050 ( n15104,n15107,n15108 );
   nor U15051 ( n15108,n15109,n15110 );
   nand U15052 ( n15110,n15111,n15112 );
   nor U15053 ( n15112,n15113,n15114 );
   nor U15054 ( n15114,n14900,n14998 );
   nor U15055 ( n15113,n14896,n15000 );
   nor U15056 ( n15111,n15115,n15116 );
   nor U15057 ( n15116,n14897,n15004 );
   nor U15058 ( n15115,n14891,n15006 );
   nand U15059 ( n15109,n15117,n15118 );
   nor U15060 ( n15118,n15119,n15120 );
   nor U15061 ( n15120,n14886,n15012 );
   nor U15062 ( n15119,n14887,n15014 );
   nor U15063 ( n15117,n15121,n15122 );
   nor U15064 ( n15122,n14879,n15018 );
   nor U15065 ( n15121,n14874,n15020 );
   nor U15066 ( n15107,n15123,n15124 );
   nand U15067 ( n15124,n15125,n15126 );
   nor U15068 ( n15126,n15127,n15128 );
   nor U15069 ( n15128,n14875,n15028 );
   nor U15070 ( n15127,n14869,n15030 );
   nor U15071 ( n15125,n15129,n15130 );
   nor U15072 ( n15130,n14864,n15034 );
   nor U15073 ( n15129,n14865,n15036 );
   nand U15074 ( n15123,n15131,n15132 );
   nor U15075 ( n15132,n15133,n15134 );
   nor U15076 ( n15134,n10801,n15041 );
   nor U15077 ( n15133,n14890,n15043 );
   nor U15078 ( n15131,n15135,n15136 );
   nor U15079 ( n15136,n14878,n15047 );
   nor U15080 ( n15135,n14868,n15049 );
   or U15081 ( n14175,n14967,n14966 );
   and U15082 ( n14966,n15137,n15138 );
   nand U15083 ( n15138,n14979,n12403 );
   nand U15084 ( n15137,instqueue_reg_0__3_,n15061 );
   xor U15085 ( n14967,n14373,n15139 );
   nand U15086 ( n15139,n15140,n15141 );
   nand U15087 ( n15141,n10466,n8821 );
   xor U15088 ( n10466,n14199,n14198 );
   nor U15089 ( n14198,n15142,n15099 );
   nand U15090 ( n15099,n15143,n15144 );
   nand U15091 ( n15144,n15145,n14982 );
   or U15092 ( n14982,n14985,n14984 );
   and U15093 ( n14984,n15146,n15147 );
   nor U15094 ( n15147,n15148,n15149 );
   nand U15095 ( n15149,n15150,n11669 );
   nand U15096 ( n11669,n15151,n9391 );
   nor U15097 ( n15151,n15152,n15153 );
   nor U15098 ( n15153,n10778,n12383 );
   nor U15099 ( n15152,n15154,n15155 );
   nand U15100 ( n15155,n15156,n10906 );
   nor U15101 ( n15156,n15157,n15158 );
   nor U15102 ( n15158,n11627,n15159 );
   nor U15103 ( n15159,n10778,n15160 );
   nand U15104 ( n15160,n15161,n13156 );
   nor U15105 ( n15157,n10798,n15162 );
   nand U15106 ( n15162,n15163,n13156 );
   nand U15107 ( n15163,n11679,n10778 );
   nand U15108 ( n15154,n10745,n15164 );
   nand U15109 ( n15150,n15165,n10808 );
   nand U15110 ( n15165,n15166,n15167 );
   nor U15111 ( n15167,n15168,n9391 );
   nor U15112 ( n15166,n11672,n11728 );
   nor U15113 ( n11672,n12874,n11708 );
   nor U15114 ( n15148,n15169,n15170 );
   nor U15115 ( n15170,n8874,n15171 );
   nor U15116 ( n15171,n15161,n11663 );
   nor U15117 ( n15169,n15172,n15173 );
   nand U15118 ( n15173,n11721,n11708 );
   nand U15119 ( n15172,n10788,n11722 );
   nor U15120 ( n15146,n15174,n9288 );
   nand U15121 ( n9288,n8960,state2_reg_0_ );
   nor U15122 ( n15174,n9391,n11627 );
   nand U15123 ( n14985,n15175,n15176 );
   nand U15124 ( n15176,n15177,n15178 );
   nand U15125 ( n15178,instqueuerd_addr_reg_0_,n15179 );
   nor U15126 ( n15177,instqueuewr_addr_reg_0_,n8858 );
   nand U15127 ( n15175,n9275,n15180 );
   nand U15128 ( n15180,n15181,n15182 );
   nand U15129 ( n15182,n15183,instqueuewr_addr_reg_0_ );
   nand U15130 ( n15181,n12469,n8968 );
   nand U15131 ( n15145,n15055,n15054 );
   or U15132 ( n15143,n15055,n15054 );
   nand U15133 ( n15054,n15184,n15185 );
   nand U15134 ( n15185,instqueuerd_addr_reg_1_,n15179 );
   nor U15135 ( n15184,n15186,n15187 );
   nor U15136 ( n15187,n9275,n9356 );
   nor U15137 ( n15186,n10126,n12469 );
   nor U15138 ( n10126,n9698,n9611 );
   nor U15139 ( n9611,n9356,instqueuewr_addr_reg_0_ );
   nor U15140 ( n9698,n15188,instqueuewr_addr_reg_1_ );
   nand U15141 ( n15055,n15189,n15190 );
   nand U15142 ( n15190,n15191,n15192 );
   nor U15143 ( n15192,n10768,n15193 );
   nand U15144 ( n15193,n10906,state2_reg_0_ );
   nor U15145 ( n15191,n11748,n11663 );
   nand U15146 ( n11663,n15168,n9391 );
   not U15147 ( n15168,n13155 );
   nand U15148 ( n13155,n11627,n11631 );
   nor U15149 ( n15189,n15194,n15195 );
   not U15150 ( n15195,n15196 );
   or U15151 ( n15142,n15101,n15100 );
   and U15152 ( n15100,n15197,n10864 );
   and U15153 ( n15101,n15197,n15183 );
   and U15154 ( n15197,n15198,n15199 );
   nand U15155 ( n15199,n8858,n9958 );
   not U15156 ( n9958,n9605 );
   xor U15157 ( n9605,instqueuewr_addr_reg_2_,n9334 );
   not U15158 ( n8858,n12469 );
   nand U15159 ( n15198,instqueuewr_addr_reg_2_,n12996 );
   nand U15160 ( n14199,n15200,n15201 );
   nand U15161 ( n15201,instqueuewr_addr_reg_3_,n12996 );
   nor U15162 ( n15200,n15202,n15203 );
   nor U15163 ( n15203,n15183,n14172 );
   not U15164 ( n15183,n15179 );
   nand U15165 ( n15179,n15204,n15205 );
   nor U15166 ( n15205,n15206,n15207 );
   nand U15167 ( n15207,n15196,n15208 );
   nand U15168 ( n15208,n15061,n11722 );
   nand U15169 ( n15196,n15209,n10914 );
   nor U15170 ( n15209,n15210,n8863 );
   nor U15171 ( n15210,n15211,n15212 );
   nor U15172 ( n15212,n15213,n12359 );
   nand U15173 ( n15206,n15214,n15215 );
   nand U15174 ( n15214,n15216,n8757 );
   nor U15175 ( n15216,n11680,n8821 );
   not U15176 ( n11680,n11728 );
   nand U15177 ( n11728,n11721,n15217 );
   nand U15178 ( n15217,n12874,n11708 );
   nor U15179 ( n15204,n15218,n15219 );
   nand U15180 ( n15219,n15220,n15221 );
   nand U15181 ( n15221,n15222,state2_reg_0_ );
   not U15182 ( n15222,n11671 );
   nand U15183 ( n15220,n12994,n15223 );
   nand U15184 ( n15223,n10788,n15164 );
   nand U15185 ( n15164,n10788,n10881 );
   nor U15186 ( n15218,n15224,n8863 );
   nor U15187 ( n15224,n15225,n15226 );
   nand U15188 ( n15226,n11627,n15227 );
   nand U15189 ( n15227,n8874,n15228 );
   nand U15190 ( n15228,n11721,n15229 );
   nand U15191 ( n15229,n11679,n15230 );
   and U15192 ( n11721,n10745,n13156 );
   nand U15193 ( n13156,n12386,n10758 );
   not U15194 ( n15225,n10894 );
   nand U15195 ( n10894,n8757,n9390 );
   nor U15196 ( n15202,n10639,n12469 );
   not U15197 ( n10639,n9959 );
   nand U15198 ( n9959,n15231,n15232 );
   nand U15199 ( n15232,instqueuewr_addr_reg_3_,n9334 );
   nor U15200 ( n15231,n9876,n10214 );
   not U15201 ( n10214,n10140 );
   nand U15202 ( n10140,n10302,n9521 );
   not U15203 ( n9521,n9334 );
   nand U15204 ( n9334,instqueuewr_addr_reg_0_,instqueuewr_addr_reg_1_ );
   nor U15205 ( n10302,n9354,instqueuewr_addr_reg_3_ );
   nor U15206 ( n9876,n9788,instqueuewr_addr_reg_2_ );
   nor U15207 ( n15140,n15233,n15234 );
   nor U15208 ( n15234,n14373,n12403 );
   nor U15209 ( n15233,n12432,n15058 );
   not U15210 ( n12432,n12403 );
   nand U15211 ( n12403,n15235,n15236 );
   nor U15212 ( n15236,n15237,n15238 );
   nand U15213 ( n15238,n15239,n15240 );
   nor U15214 ( n15240,n15241,n15242 );
   nor U15215 ( n15242,n15243,n14998 );
   nor U15216 ( n15241,n15244,n15000 );
   nor U15217 ( n15239,n15245,n15246 );
   nor U15218 ( n15246,n15247,n15004 );
   nor U15219 ( n15245,n15248,n15006 );
   nand U15220 ( n15237,n15249,n15250 );
   nor U15221 ( n15250,n15251,n15252 );
   nor U15222 ( n15252,n15253,n15012 );
   nor U15223 ( n15251,n15254,n15014 );
   nor U15224 ( n15249,n15255,n15256 );
   nor U15225 ( n15256,n15257,n15018 );
   nor U15226 ( n15255,n15258,n15020 );
   nor U15227 ( n15235,n15259,n15260 );
   nand U15228 ( n15260,n15261,n15262 );
   nor U15229 ( n15262,n15263,n15264 );
   nor U15230 ( n15264,n15265,n15028 );
   nor U15231 ( n15263,n15266,n15030 );
   nor U15232 ( n15261,n15267,n15268 );
   nor U15233 ( n15268,n15269,n15034 );
   nor U15234 ( n15267,n15270,n15036 );
   nand U15235 ( n15259,n15271,n15272 );
   nor U15236 ( n15272,n15273,n15274 );
   nor U15237 ( n15274,n10791,n15041 );
   nor U15238 ( n15273,n15275,n15043 );
   nor U15239 ( n15271,n15276,n15277 );
   nor U15240 ( n15277,n15278,n15047 );
   nor U15241 ( n15276,n15279,n15049 );
   nand U15242 ( n14189,n14963,n14962 );
   nand U15243 ( n14962,n15280,n15281 );
   nand U15244 ( n15281,n14979,n12407 );
   nand U15245 ( n15280,n15061,instqueue_reg_0__4_ );
   and U15246 ( n14963,n15282,n12407 );
   nand U15247 ( n12407,n15283,n15284 );
   nor U15248 ( n15284,n15285,n15286 );
   nand U15249 ( n15286,n15287,n15288 );
   nor U15250 ( n15288,n15289,n15290 );
   nor U15251 ( n15290,n15291,n14998 );
   nor U15252 ( n15289,n15292,n15000 );
   nor U15253 ( n15287,n15293,n15294 );
   nor U15254 ( n15294,n15295,n15004 );
   nor U15255 ( n15293,n15296,n15006 );
   nand U15256 ( n15285,n15297,n15298 );
   nor U15257 ( n15298,n15299,n15300 );
   nor U15258 ( n15300,n15301,n15012 );
   nor U15259 ( n15299,n15302,n15014 );
   nor U15260 ( n15297,n15303,n15304 );
   nor U15261 ( n15304,n15305,n15018 );
   nor U15262 ( n15303,n15306,n15020 );
   nor U15263 ( n15283,n15307,n15308 );
   nand U15264 ( n15308,n15309,n15310 );
   nor U15265 ( n15310,n15311,n15312 );
   nor U15266 ( n15312,n15313,n15028 );
   nor U15267 ( n15311,n15314,n15030 );
   nor U15268 ( n15309,n15315,n15316 );
   nor U15269 ( n15316,n15317,n15034 );
   nor U15270 ( n15315,n15318,n15036 );
   nand U15271 ( n15307,n15319,n15320 );
   nor U15272 ( n15320,n15321,n15322 );
   nor U15273 ( n15322,n10781,n15041 );
   nor U15274 ( n15321,n15323,n15043 );
   nor U15275 ( n15319,n15324,n15325 );
   nor U15276 ( n15325,n15326,n15047 );
   nor U15277 ( n15324,n15327,n15049 );
   nor U15278 ( n14081,n14960,n14959 );
   and U15279 ( n14959,n15328,n15329 );
   nand U15280 ( n15329,n14979,n12417 );
   nand U15281 ( n15328,n15061,instqueue_reg_0__5_ );
   nand U15282 ( n14960,n15282,n12417 );
   nand U15283 ( n12417,n15330,n15331 );
   nor U15284 ( n15331,n15332,n15333 );
   nand U15285 ( n15333,n15334,n15335 );
   nor U15286 ( n15335,n15336,n15337 );
   nor U15287 ( n15337,n15338,n14998 );
   nor U15288 ( n15336,n15339,n15000 );
   nor U15289 ( n15334,n15340,n15341 );
   nor U15290 ( n15341,n15342,n15004 );
   nor U15291 ( n15340,n15343,n15006 );
   nand U15292 ( n15332,n15344,n15345 );
   nor U15293 ( n15345,n15346,n15347 );
   nor U15294 ( n15347,n15348,n15012 );
   nor U15295 ( n15346,n15349,n15014 );
   nor U15296 ( n15344,n15350,n15351 );
   nor U15297 ( n15351,n15352,n15018 );
   nor U15298 ( n15350,n15353,n15020 );
   nor U15299 ( n15330,n15354,n15355 );
   nand U15300 ( n15355,n15356,n15357 );
   nor U15301 ( n15357,n15358,n15359 );
   nor U15302 ( n15359,n15360,n15028 );
   nor U15303 ( n15358,n15361,n15030 );
   nor U15304 ( n15356,n15362,n15363 );
   nor U15305 ( n15363,n15364,n15034 );
   nor U15306 ( n15362,n15365,n15036 );
   nand U15307 ( n15354,n15366,n15367 );
   nor U15308 ( n15367,n15368,n15369 );
   nor U15309 ( n15369,n10771,n15041 );
   nor U15310 ( n15368,n15370,n15043 );
   nor U15311 ( n15366,n15371,n15372 );
   nor U15312 ( n15372,n15373,n15047 );
   nor U15313 ( n15371,n15374,n15049 );
   nand U15314 ( n14207,n14957,n14956 );
   nand U15315 ( n14956,n15375,n15376 );
   nand U15316 ( n15376,n14979,n12434 );
   nand U15317 ( n15375,instqueue_reg_0__6_,n15061 );
   and U15318 ( n14957,n15282,n12434 );
   nand U15319 ( n12434,n15377,n15378 );
   nor U15320 ( n15378,n15379,n15380 );
   nand U15321 ( n15380,n15381,n15382 );
   nor U15322 ( n15382,n15383,n15384 );
   nor U15323 ( n15384,n14766,n14998 );
   nor U15324 ( n15383,n14767,n15000 );
   nor U15325 ( n15381,n15385,n15386 );
   nor U15326 ( n15386,n14770,n15004 );
   nor U15327 ( n15385,n14757,n15006 );
   nand U15328 ( n15379,n15387,n15388 );
   nor U15329 ( n15388,n15389,n15390 );
   nor U15330 ( n15390,n14758,n15012 );
   nor U15331 ( n15389,n14761,n15014 );
   nor U15332 ( n15387,n15391,n15392 );
   nor U15333 ( n15392,n14789,n15018 );
   nor U15334 ( n15391,n14792,n15020 );
   nor U15335 ( n15377,n15393,n15394 );
   nand U15336 ( n15394,n15395,n15396 );
   nor U15337 ( n15396,n15397,n15398 );
   nor U15338 ( n15398,n14793,n15028 );
   nor U15339 ( n15397,n14779,n15030 );
   nor U15340 ( n15395,n15399,n15400 );
   nor U15341 ( n15400,n14782,n15034 );
   nor U15342 ( n15399,n14783,n15036 );
   nand U15343 ( n15393,n15401,n15402 );
   nor U15344 ( n15402,n15403,n15404 );
   nor U15345 ( n15404,n10761,n15041 );
   nor U15346 ( n15403,n14771,n15043 );
   nor U15347 ( n15401,n15405,n15406 );
   nor U15348 ( n15406,n14788,n15047 );
   nor U15349 ( n15405,n14778,n15049 );
   nand U15350 ( n15282,n8796,n15058 );
   nand U15351 ( n15058,n12357,n15407 );
   not U15352 ( n12357,n12430 );
   nand U15353 ( n14223,n12454,n14954 );
   nand U15354 ( n14954,n15408,n15409 );
   nand U15355 ( n15409,n14979,n12430 );
   nand U15356 ( n15408,instqueue_reg_0__7_,n15061 );
   nand U15357 ( n14261,n15410,n14797 );
   nor U15358 ( n15410,n15411,n15412 );
   nor U15359 ( n15412,n14373,n15413 );
   nor U15360 ( n15411,n15414,n14802 );
   not U15361 ( n15414,n15413 );
   nand U15362 ( n15413,n15415,n15416 );
   nor U15363 ( n15416,n15417,n15418 );
   nand U15364 ( n15418,n15419,n15420 );
   nor U15365 ( n15420,n15421,n15422 );
   nor U15366 ( n15422,n15033,n14811 );
   nor U15367 ( n15421,n15035,n14812 );
   nor U15368 ( n15419,n15423,n15424 );
   nor U15369 ( n15424,n15048,n14815 );
   nor U15370 ( n15423,n15029,n14816 );
   nand U15371 ( n15417,n15425,n15426 );
   nor U15372 ( n15426,n15427,n15428 );
   nor U15373 ( n15428,n15019,n14821 );
   nor U15374 ( n15427,n15027,n14822 );
   nor U15375 ( n15425,n15429,n15430 );
   nor U15376 ( n15430,n15046,n14825 );
   nor U15377 ( n15429,n15017,n14826 );
   nor U15378 ( n15415,n15431,n15432 );
   nand U15379 ( n15432,n15433,n15434 );
   nor U15380 ( n15434,n15435,n15436 );
   nor U15381 ( n15436,n15011,n14833 );
   nor U15382 ( n15435,n15013,n14834 );
   nor U15383 ( n15433,n15437,n15438 );
   nor U15384 ( n15438,n15042,n14837 );
   nor U15385 ( n15437,n15005,n14838 );
   nand U15386 ( n15431,n15439,n15440 );
   nor U15387 ( n15440,n15441,n15442 );
   nor U15388 ( n15442,n14999,n14843 );
   nor U15389 ( n15441,n15003,n14844 );
   nor U15390 ( n15439,n15443,n15444 );
   nor U15391 ( n15444,n10825,n14847 );
   nor U15392 ( n15443,n14997,n14848 );
   nor U15393 ( n14850,n15445,n14301 );
   xor U15394 ( n14301,n15446,n14373 );
   nor U15395 ( n15446,n15447,n14971 );
   nor U15396 ( n15447,n15448,n15449 );
   nand U15397 ( n15449,n15450,n15451 );
   nor U15398 ( n15451,n15452,n15453 );
   nand U15399 ( n15453,n15454,n15455 );
   nand U15400 ( n15455,n15456,instqueue_reg_1__4_ );
   nand U15401 ( n15454,n15457,instqueue_reg_0__4_ );
   nand U15402 ( n15452,n15458,n15459 );
   nand U15403 ( n15459,n15460,instqueue_reg_3__4_ );
   nand U15404 ( n15458,n15461,instqueue_reg_2__4_ );
   nor U15405 ( n15450,n15462,n15463 );
   nand U15406 ( n15463,n15464,n15465 );
   nand U15407 ( n15465,n15466,instqueue_reg_5__4_ );
   nand U15408 ( n15464,n15467,instqueue_reg_4__4_ );
   nand U15409 ( n15462,n15468,n15469 );
   nand U15410 ( n15469,n15470,instqueue_reg_7__4_ );
   nand U15411 ( n15468,n15471,instqueue_reg_6__4_ );
   nand U15412 ( n15448,n15472,n15473 );
   nor U15413 ( n15473,n15474,n15475 );
   nand U15414 ( n15475,n15476,n15477 );
   nand U15415 ( n15477,n15478,instqueue_reg_9__4_ );
   nand U15416 ( n15476,n15479,instqueue_reg_8__4_ );
   nand U15417 ( n15474,n15480,n15481 );
   nand U15418 ( n15481,n15482,instqueue_reg_11__4_ );
   nand U15419 ( n15480,n15483,instqueue_reg_10__4_ );
   nor U15420 ( n15472,n15484,n15485 );
   nand U15421 ( n15485,n15486,n15487 );
   nand U15422 ( n15487,n15488,instqueue_reg_13__4_ );
   nand U15423 ( n15486,n15489,instqueue_reg_12__4_ );
   nand U15424 ( n15484,n15490,n15491 );
   nand U15425 ( n15491,n15492,instqueue_reg_15__4_ );
   nand U15426 ( n15490,n15493,instqueue_reg_14__4_ );
   not U15427 ( n15445,n14243 );
   nand U15428 ( n14243,n15494,n14797 );
   nor U15429 ( n15494,n15495,n15496 );
   nor U15430 ( n15496,n8796,n15497 );
   nor U15431 ( n15495,n15498,n14802 );
   not U15432 ( n15498,n15497 );
   nand U15433 ( n15497,n15499,n15500 );
   nor U15434 ( n15500,n15501,n15502 );
   nand U15435 ( n15502,n15503,n15504 );
   nor U15436 ( n15504,n15505,n15506 );
   nor U15437 ( n15506,n15269,n14811 );
   nor U15438 ( n15505,n15270,n14812 );
   nor U15439 ( n15503,n15507,n15508 );
   nor U15440 ( n15508,n15279,n14815 );
   nor U15441 ( n15507,n15266,n14816 );
   nand U15442 ( n15501,n15509,n15510 );
   nor U15443 ( n15510,n15511,n15512 );
   nor U15444 ( n15512,n15258,n14821 );
   nor U15445 ( n15511,n15265,n14822 );
   nor U15446 ( n15509,n15513,n15514 );
   nor U15447 ( n15514,n15278,n14825 );
   nor U15448 ( n15513,n15257,n14826 );
   nor U15449 ( n15499,n15515,n15516 );
   nand U15450 ( n15516,n15517,n15518 );
   nor U15451 ( n15518,n15519,n15520 );
   nor U15452 ( n15520,n15253,n14833 );
   nor U15453 ( n15519,n15254,n14834 );
   nor U15454 ( n15517,n15521,n15522 );
   nor U15455 ( n15522,n15275,n14837 );
   nor U15456 ( n15521,n15248,n14838 );
   nand U15457 ( n15515,n15523,n15524 );
   nor U15458 ( n15524,n15525,n15526 );
   nor U15459 ( n15526,n15244,n14843 );
   nor U15460 ( n15525,n15247,n14844 );
   nor U15461 ( n15523,n15527,n15528 );
   nor U15462 ( n15528,n10791,n14847 );
   nor U15463 ( n15527,n15243,n14848 );
   nor U15464 ( n14849,n15529,n14313 );
   xor U15465 ( n14313,n15530,n14373 );
   nor U15466 ( n15530,n15531,n14971 );
   nor U15467 ( n15531,n15532,n15533 );
   nand U15468 ( n15533,n15534,n15535 );
   nor U15469 ( n15535,n15536,n15537 );
   nand U15470 ( n15537,n15538,n15539 );
   nand U15471 ( n15539,n15456,instqueue_reg_1__6_ );
   not U15472 ( n15456,n14848 );
   nand U15473 ( n15538,n15457,instqueue_reg_0__6_ );
   not U15474 ( n15457,n14847 );
   nand U15475 ( n15536,n15540,n15541 );
   nand U15476 ( n15541,n15460,instqueue_reg_3__6_ );
   not U15477 ( n15460,n14844 );
   nand U15478 ( n15540,n15461,instqueue_reg_2__6_ );
   not U15479 ( n15461,n14843 );
   nor U15480 ( n15534,n15542,n15543 );
   nand U15481 ( n15543,n15544,n15545 );
   nand U15482 ( n15545,n15466,instqueue_reg_5__6_ );
   not U15483 ( n15466,n14838 );
   nand U15484 ( n15544,n15467,instqueue_reg_4__6_ );
   not U15485 ( n15467,n14837 );
   nand U15486 ( n15542,n15546,n15547 );
   nand U15487 ( n15547,n15470,instqueue_reg_7__6_ );
   not U15488 ( n15470,n14834 );
   nand U15489 ( n15546,n15471,instqueue_reg_6__6_ );
   not U15490 ( n15471,n14833 );
   nand U15491 ( n15532,n15548,n15549 );
   nor U15492 ( n15549,n15550,n15551 );
   nand U15493 ( n15551,n15552,n15553 );
   nand U15494 ( n15553,n15478,instqueue_reg_9__6_ );
   not U15495 ( n15478,n14826 );
   nand U15496 ( n15552,n15479,instqueue_reg_8__6_ );
   not U15497 ( n15479,n14825 );
   nand U15498 ( n15550,n15554,n15555 );
   nand U15499 ( n15555,n15482,instqueue_reg_11__6_ );
   not U15500 ( n15482,n14822 );
   nand U15501 ( n15554,n15483,instqueue_reg_10__6_ );
   not U15502 ( n15483,n14821 );
   nor U15503 ( n15548,n15556,n15557 );
   nand U15504 ( n15557,n15558,n15559 );
   nand U15505 ( n15559,n15488,instqueue_reg_13__6_ );
   not U15506 ( n15488,n14816 );
   nand U15507 ( n15558,n15489,instqueue_reg_12__6_ );
   not U15508 ( n15489,n14815 );
   nand U15509 ( n15556,n15560,n15561 );
   nand U15510 ( n15561,n15492,instqueue_reg_15__6_ );
   not U15511 ( n15492,n14812 );
   nand U15512 ( n15560,n15493,instqueue_reg_14__6_ );
   not U15513 ( n15493,n14811 );
   not U15514 ( n15529,n14304 );
   nand U15515 ( n14304,n15562,n14797 );
   nand U15516 ( n14797,n14971,n12454 );
   nor U15517 ( n15562,n15563,n15564 );
   nor U15518 ( n15564,n8796,n15565 );
   nor U15519 ( n15563,n15566,n14802 );
   or U15520 ( n14802,n12454,n14971 );
   nor U15521 ( n14971,n15061,n14979 );
   not U15522 ( n12454,n14373 );
   nand U15523 ( n14373,n15407,n12430 );
   nand U15524 ( n12430,n15567,n15568 );
   nor U15525 ( n15568,n15569,n15570 );
   nand U15526 ( n15570,n15571,n15572 );
   nor U15527 ( n15572,n15573,n15574 );
   nor U15528 ( n15574,n14694,n14998 );
   nand U15529 ( n14998,n15575,n15576 );
   nor U15530 ( n15573,n14696,n15000 );
   nand U15531 ( n15000,n15575,n15577 );
   nor U15532 ( n15571,n15578,n15579 );
   nor U15533 ( n15579,n14700,n15004 );
   nand U15534 ( n15004,n15575,n15580 );
   nor U15535 ( n15578,n14681,n15006 );
   nand U15536 ( n15006,n15576,n15581 );
   nand U15537 ( n15569,n15582,n15583 );
   nor U15538 ( n15583,n15584,n15585 );
   nor U15539 ( n15585,n14683,n15012 );
   nand U15540 ( n15012,n15577,n15581 );
   nor U15541 ( n15584,n14687,n15014 );
   nand U15542 ( n15014,n15580,n15581 );
   nor U15543 ( n15582,n15586,n15587 );
   nor U15544 ( n15587,n14726,n15018 );
   nand U15545 ( n15018,n15576,n15588 );
   nor U15546 ( n15586,n14730,n15020 );
   nand U15547 ( n15020,n15588,n15577 );
   nor U15548 ( n15567,n15589,n15590 );
   nand U15549 ( n15590,n15591,n15592 );
   nor U15550 ( n15592,n15593,n15594 );
   nor U15551 ( n15594,n14732,n15028 );
   nand U15552 ( n15028,n15588,n15580 );
   nor U15553 ( n15593,n14712,n15030 );
   nand U15554 ( n15030,n15595,n15576 );
   nor U15555 ( n15591,n15596,n15597 );
   nor U15556 ( n15597,n14716,n15034 );
   nand U15557 ( n15034,n15595,n15577 );
   nor U15558 ( n15596,n14718,n15036 );
   nand U15559 ( n15036,n15595,n15580 );
   nand U15560 ( n15589,n15598,n15599 );
   nor U15561 ( n15599,n15600,n15601 );
   nor U15562 ( n15601,n10750,n15041 );
   nand U15563 ( n15041,n15602,n15575 );
   nor U15564 ( n15575,n9005,n8989 );
   nor U15565 ( n15600,n14702,n15043 );
   nand U15566 ( n15043,n15602,n15581 );
   nor U15567 ( n15581,n9005,n10878 );
   nor U15568 ( n15598,n15603,n15604 );
   nor U15569 ( n15604,n14724,n15047 );
   nand U15570 ( n15047,n15602,n15588 );
   nor U15571 ( n15588,n8989,n10854 );
   not U15572 ( n8989,n10878 );
   nor U15573 ( n15603,n14710,n15049 );
   nand U15574 ( n15049,n15595,n15602 );
   nor U15575 ( n15595,n10878,n10854 );
   not U15576 ( n10854,n9005 );
   nand U15577 ( n9005,n15605,n15606 );
   or U15578 ( n15606,n14172,n15607 );
   nor U15579 ( n10878,n15608,n15609 );
   nor U15580 ( n15608,n10864,n10861 );
   not U15581 ( n15566,n15565 );
   nand U15582 ( n15565,n15610,n15611 );
   nor U15583 ( n15611,n15612,n15613 );
   nand U15584 ( n15613,n15614,n15615 );
   nor U15585 ( n15615,n15616,n15617 );
   nor U15586 ( n15617,n15364,n14811 );
   nand U15587 ( n14811,n15618,n15619 );
   nor U15588 ( n15616,n15365,n14812 );
   nand U15589 ( n14812,n15618,n15620 );
   nor U15590 ( n15614,n15621,n15622 );
   nor U15591 ( n15622,n15374,n14815 );
   nand U15592 ( n14815,n15618,n15623 );
   nor U15593 ( n15621,n15361,n14816 );
   nand U15594 ( n14816,n15618,n10861 );
   nor U15595 ( n15618,n10867,n10884 );
   nand U15596 ( n15612,n15624,n15625 );
   nor U15597 ( n15625,n15626,n15627 );
   nor U15598 ( n15627,n15353,n14821 );
   nand U15599 ( n14821,n15628,n15619 );
   nor U15600 ( n15626,n15360,n14822 );
   nand U15601 ( n14822,n15628,n15620 );
   nor U15602 ( n15624,n15629,n15630 );
   nor U15603 ( n15630,n15373,n14825 );
   nand U15604 ( n14825,n15628,n15623 );
   nor U15605 ( n15629,n15352,n14826 );
   nand U15606 ( n14826,n15628,n10861 );
   nor U15607 ( n15628,n15631,n10867 );
   nor U15608 ( n15610,n15632,n15633 );
   nand U15609 ( n15633,n15634,n15635 );
   nor U15610 ( n15635,n15636,n15637 );
   nor U15611 ( n15637,n15348,n14833 );
   nand U15612 ( n14833,n15638,n15619 );
   nor U15613 ( n15636,n15349,n14834 );
   nand U15614 ( n14834,n15638,n15620 );
   nor U15615 ( n15634,n15639,n15640 );
   nor U15616 ( n15640,n15370,n14837 );
   nand U15617 ( n14837,n15638,n15623 );
   nor U15618 ( n15639,n15343,n14838 );
   nand U15619 ( n14838,n15638,n10861 );
   nor U15620 ( n15638,n10884,n15641 );
   nand U15621 ( n15632,n15642,n15643 );
   nor U15622 ( n15643,n15644,n15645 );
   nor U15623 ( n15645,n15339,n14843 );
   nand U15624 ( n14843,n15646,n15619 );
   nor U15625 ( n15644,n15342,n14844 );
   nand U15626 ( n14844,n15646,n15620 );
   nor U15627 ( n15642,n15647,n15648 );
   nor U15628 ( n15648,n10771,n14847 );
   nand U15629 ( n14847,n15646,n15623 );
   nor U15630 ( n15647,n15338,n14848 );
   nand U15631 ( n14848,n15646,n10861 );
   nor U15632 ( n15646,n15631,n15641 );
   not U15633 ( n15641,n10867 );
   nand U15634 ( n10867,n15649,n15650 );
   nand U15635 ( n15650,n15651,instqueuerd_addr_reg_2_ );
   nor U15636 ( n15651,n15652,n9339 );
   nand U15637 ( n15649,n15653,n14172 );
   nand U15638 ( n15653,n15652,instqueuerd_addr_reg_1_ );
   not U15639 ( n15631,n10884 );
   xor U15640 ( n10884,instqueuerd_addr_reg_2_,n9339 );
   xor U15641 ( n13952,n8764,n15654 );
   nand U15642 ( n15654,n15655,n15656 );
   nor U15643 ( n15656,n15657,n15658 );
   nor U15644 ( n15658,n8765,n12262 );
   nand U15645 ( n12262,n15659,n14745 );
   nand U15646 ( n15659,n12265,n14458 );
   nor U15647 ( n15657,n15660,n15661 );
   nor U15648 ( n15661,n15662,n15663 );
   not U15649 ( n15660,n14668 );
   nand U15650 ( n14668,n15662,n15663 );
   and U15651 ( n15663,n15664,n14572 );
   nand U15652 ( n15664,n15665,n15666 );
   nor U15653 ( n15666,n15667,n15668 );
   nand U15654 ( n15668,n15669,n15670 );
   nor U15655 ( n15670,n15671,n15672 );
   nor U15656 ( n15672,n15373,n14725 );
   nor U15657 ( n15671,n15352,n14727 );
   nor U15658 ( n15669,n15673,n15674 );
   nor U15659 ( n15674,n15353,n14731 );
   nor U15660 ( n15673,n15360,n14733 );
   nand U15661 ( n15667,n15675,n15676 );
   nor U15662 ( n15676,n15677,n15678 );
   nor U15663 ( n15678,n15374,n14711 );
   nor U15664 ( n15677,n15361,n14713 );
   nor U15665 ( n15675,n15679,n15680 );
   nor U15666 ( n15680,n15364,n14717 );
   nor U15667 ( n15679,n15365,n14719 );
   nor U15668 ( n15665,n15681,n15682 );
   nand U15669 ( n15682,n15683,n15684 );
   nor U15670 ( n15684,n15685,n15686 );
   nor U15671 ( n15686,n15338,n14695 );
   nor U15672 ( n15685,n15339,n14697 );
   nor U15673 ( n15683,n15687,n15688 );
   nor U15674 ( n15688,n15342,n14701 );
   nor U15675 ( n15687,n15370,n14703 );
   nand U15676 ( n15681,n15689,n15690 );
   nor U15677 ( n15690,n15691,n15692 );
   nor U15678 ( n15692,n15343,n14682 );
   nor U15679 ( n15691,n15348,n14684 );
   nor U15680 ( n15689,n15693,n15694 );
   nor U15681 ( n15694,n15349,n14688 );
   nor U15682 ( n15693,n10771,n14689 );
   nor U15683 ( n15662,n14464,n14463 );
   nand U15684 ( n14463,n14572,n15695 );
   nand U15685 ( n15695,n15696,n15697 );
   nor U15686 ( n15697,n15698,n15699 );
   nand U15687 ( n15699,n15700,n15701 );
   nor U15688 ( n15701,n15702,n15703 );
   nor U15689 ( n15703,n15296,n14682 );
   nor U15690 ( n15702,n15301,n14684 );
   nor U15691 ( n15700,n15704,n15705 );
   nor U15692 ( n15705,n15302,n14688 );
   nor U15693 ( n15704,n10781,n14689 );
   nand U15694 ( n15698,n15706,n15707 );
   nor U15695 ( n15707,n15708,n15709 );
   nor U15696 ( n15709,n15291,n14695 );
   nor U15697 ( n15708,n15292,n14697 );
   nor U15698 ( n15706,n15710,n15711 );
   nor U15699 ( n15711,n15295,n14701 );
   nor U15700 ( n15710,n15323,n14703 );
   nor U15701 ( n15696,n15712,n15713 );
   nand U15702 ( n15713,n15714,n15715 );
   nor U15703 ( n15715,n15716,n15717 );
   nor U15704 ( n15717,n15327,n14711 );
   nor U15705 ( n15716,n15314,n14713 );
   nor U15706 ( n15714,n15718,n15719 );
   nor U15707 ( n15719,n15317,n14717 );
   nor U15708 ( n15718,n15318,n14719 );
   nand U15709 ( n15712,n15720,n15721 );
   nor U15710 ( n15721,n15722,n15723 );
   nor U15711 ( n15723,n15326,n14725 );
   nor U15712 ( n15722,n15305,n14727 );
   nor U15713 ( n15720,n15724,n15725 );
   nor U15714 ( n15725,n15306,n14731 );
   nor U15715 ( n15724,n15313,n14733 );
   nand U15716 ( n14464,n14474,n14475 );
   and U15717 ( n14475,n14572,n15726 );
   nand U15718 ( n15726,n15727,n15728 );
   nor U15719 ( n15728,n15729,n15730 );
   nand U15720 ( n15730,n15731,n15732 );
   nor U15721 ( n15732,n15733,n15734 );
   nor U15722 ( n15734,n15248,n14682 );
   nor U15723 ( n15733,n15253,n14684 );
   nor U15724 ( n15731,n15735,n15736 );
   nor U15725 ( n15736,n15254,n14688 );
   nor U15726 ( n15735,n10791,n14689 );
   nand U15727 ( n15729,n15737,n15738 );
   nor U15728 ( n15738,n15739,n15740 );
   nor U15729 ( n15740,n15243,n14695 );
   nor U15730 ( n15739,n15244,n14697 );
   nor U15731 ( n15737,n15741,n15742 );
   nor U15732 ( n15742,n15247,n14701 );
   nor U15733 ( n15741,n15275,n14703 );
   nor U15734 ( n15727,n15743,n15744 );
   nand U15735 ( n15744,n15745,n15746 );
   nor U15736 ( n15746,n15747,n15748 );
   nor U15737 ( n15748,n15279,n14711 );
   nor U15738 ( n15747,n15266,n14713 );
   nor U15739 ( n15745,n15749,n15750 );
   nor U15740 ( n15750,n15269,n14717 );
   nor U15741 ( n15749,n15270,n14719 );
   nand U15742 ( n15743,n15751,n15752 );
   nor U15743 ( n15752,n15753,n15754 );
   nor U15744 ( n15754,n15278,n14725 );
   nor U15745 ( n15753,n15257,n14727 );
   nor U15746 ( n15751,n15755,n15756 );
   nor U15747 ( n15756,n15258,n14731 );
   nor U15748 ( n15755,n15265,n14733 );
   nor U15749 ( n14474,n14655,n14629 );
   nand U15750 ( n14629,n15757,n14644 );
   not U15751 ( n14644,n14633 );
   nand U15752 ( n14633,n14572,n15758 );
   nand U15753 ( n15758,n15759,n15760 );
   nor U15754 ( n15760,n15761,n15762 );
   nand U15755 ( n15762,n15763,n15764 );
   nor U15756 ( n15764,n15765,n15766 );
   nor U15757 ( n15766,n15005,n14682 );
   nor U15758 ( n15765,n15011,n14684 );
   nor U15759 ( n15763,n15767,n15768 );
   nor U15760 ( n15768,n15013,n14688 );
   nor U15761 ( n15767,n10825,n14689 );
   nand U15762 ( n15761,n15769,n15770 );
   nor U15763 ( n15770,n15771,n15772 );
   nor U15764 ( n15772,n14997,n14695 );
   nor U15765 ( n15771,n14999,n14697 );
   nor U15766 ( n15769,n15773,n15774 );
   nor U15767 ( n15774,n15003,n14701 );
   nor U15768 ( n15773,n15042,n14703 );
   nor U15769 ( n15759,n15775,n15776 );
   nand U15770 ( n15776,n15777,n15778 );
   nor U15771 ( n15778,n15779,n15780 );
   nor U15772 ( n15780,n15048,n14711 );
   nor U15773 ( n15779,n15029,n14713 );
   nor U15774 ( n15777,n15781,n15782 );
   nor U15775 ( n15782,n15033,n14717 );
   nor U15776 ( n15781,n15035,n14719 );
   nand U15777 ( n15775,n15783,n15784 );
   nor U15778 ( n15784,n15785,n15786 );
   nor U15779 ( n15786,n15046,n14725 );
   nor U15780 ( n15785,n15017,n14727 );
   nor U15781 ( n15783,n15787,n15788 );
   nor U15782 ( n15788,n15019,n14731 );
   nor U15783 ( n15787,n15027,n14733 );
   nor U15784 ( n15757,n15789,n14634 );
   nand U15785 ( n14634,n14572,n15790 );
   nand U15786 ( n15790,n15791,n15792 );
   nor U15787 ( n15792,n15793,n15794 );
   nand U15788 ( n15794,n15795,n15796 );
   nor U15789 ( n15796,n15797,n15798 );
   nor U15790 ( n15798,n14702,n14613 );
   nand U15791 ( n14613,n15799,n15577 );
   nor U15792 ( n15797,n14681,n14617 );
   nand U15793 ( n14617,n15799,n15580 );
   nor U15794 ( n15795,n15800,n15801 );
   nor U15795 ( n15801,n14683,n14618 );
   nand U15796 ( n14618,n15799,n15602 );
   nor U15797 ( n15800,n14687,n14585 );
   nand U15798 ( n14585,n15799,n15576 );
   nor U15799 ( n15799,n15802,n15803 );
   nand U15800 ( n15793,n15804,n15805 );
   nor U15801 ( n15805,n15806,n15807 );
   nor U15802 ( n15807,n10750,n14608 );
   nand U15803 ( n14608,n15808,n15577 );
   nor U15804 ( n15806,n14694,n14607 );
   nand U15805 ( n14607,n15808,n15580 );
   nor U15806 ( n15804,n15809,n15810 );
   nor U15807 ( n15810,n14696,n14614 );
   nand U15808 ( n14614,n15808,n15602 );
   nor U15809 ( n15809,n14700,n14586 );
   nand U15810 ( n14586,n15808,n15576 );
   nor U15811 ( n15808,n15802,n15811 );
   nor U15812 ( n15791,n15812,n15813 );
   nand U15813 ( n15813,n15814,n15815 );
   nor U15814 ( n15815,n15816,n15817 );
   nor U15815 ( n15817,n14710,n14595 );
   nand U15816 ( n14595,n15818,n15577 );
   nor U15817 ( n15816,n14712,n14603 );
   nand U15818 ( n14603,n15818,n15580 );
   nor U15819 ( n15814,n15819,n15820 );
   nor U15820 ( n15820,n14716,n14604 );
   nand U15821 ( n14604,n15818,n15602 );
   nor U15822 ( n15819,n14718,n14581 );
   nand U15823 ( n14581,n15818,n15576 );
   nor U15824 ( n15818,n15803,n15821 );
   not U15825 ( n15803,n15811 );
   nand U15826 ( n15812,n15822,n15823 );
   nor U15827 ( n15823,n15824,n15825 );
   nor U15828 ( n15825,n14724,n14592 );
   nand U15829 ( n14592,n15826,n15577 );
   nor U15830 ( n15577,n15827,n8968 );
   nor U15831 ( n15824,n14726,n14591 );
   nand U15832 ( n14591,n15826,n15580 );
   nor U15833 ( n15580,n15827,instqueuerd_addr_reg_0_ );
   nor U15834 ( n15822,n15828,n15829 );
   nor U15835 ( n15829,n14730,n14596 );
   nand U15836 ( n14596,n15826,n15602 );
   nor U15837 ( n15602,n8968,n8977 );
   nor U15838 ( n15828,n14732,n14582 );
   nand U15839 ( n14582,n15826,n15576 );
   nor U15840 ( n15576,n8977,instqueuerd_addr_reg_0_ );
   not U15841 ( n8977,n15827 );
   nand U15842 ( n15827,n15830,n10868 );
   nor U15843 ( n15826,n15821,n15811 );
   nor U15844 ( n15811,n15831,n15832 );
   not U15845 ( n15821,n15802 );
   nand U15846 ( n15802,n15833,n15834 );
   or U15847 ( n15834,n14172,n15831 );
   nor U15848 ( n15831,n10864,n15619 );
   nand U15849 ( n15833,n15652,n10868 );
   not U15850 ( n15789,n14632 );
   nand U15851 ( n14632,n15835,n15836 );
   nor U15852 ( n15836,n15837,n15838 );
   nand U15853 ( n15838,n15839,n15840 );
   nor U15854 ( n15840,n15841,n15842 );
   nor U15855 ( n15842,n14929,n14725 );
   nor U15856 ( n15841,n14930,n14727 );
   nor U15857 ( n15839,n15843,n15844 );
   nor U15858 ( n15844,n14925,n14731 );
   nor U15859 ( n15843,n14926,n14733 );
   nand U15860 ( n15837,n15845,n15846 );
   nor U15861 ( n15846,n15847,n15848 );
   nor U15862 ( n15848,n14919,n14711 );
   nor U15863 ( n15847,n14920,n14713 );
   nor U15864 ( n15845,n15849,n15850 );
   nor U15865 ( n15850,n14915,n14717 );
   nor U15866 ( n15849,n14916,n14719 );
   nor U15867 ( n15835,n15851,n15852 );
   nand U15868 ( n15852,n15853,n15854 );
   nor U15869 ( n15854,n15855,n15856 );
   nor U15870 ( n15856,n14951,n14695 );
   nor U15871 ( n15855,n14947,n14697 );
   nor U15872 ( n15853,n15857,n15858 );
   nor U15873 ( n15858,n14948,n14701 );
   nor U15874 ( n15857,n14941,n14703 );
   nand U15875 ( n15851,n15859,n15860 );
   nor U15876 ( n15860,n15861,n15862 );
   nor U15877 ( n15862,n14942,n14682 );
   nor U15878 ( n15861,n14937,n14684 );
   nor U15879 ( n15859,n15863,n15864 );
   nor U15880 ( n15864,n14938,n14688 );
   nor U15881 ( n15863,n10811,n14689 );
   nand U15882 ( n14655,n14572,n15865 );
   nand U15883 ( n15865,n15866,n15867 );
   nor U15884 ( n15867,n15868,n15869 );
   nand U15885 ( n15869,n15870,n15871 );
   nor U15886 ( n15871,n15872,n15873 );
   nor U15887 ( n15873,n14891,n14682 );
   nand U15888 ( n14682,n15874,n15875 );
   nor U15889 ( n15874,instqueuerd_addr_reg_2_,n15876 );
   nor U15890 ( n15872,n14886,n14684 );
   nand U15891 ( n14684,n15877,n15875 );
   nor U15892 ( n15877,instqueuerd_addr_reg_2_,n15878 );
   nor U15893 ( n15870,n15879,n15880 );
   nor U15894 ( n15880,n14887,n14688 );
   nand U15895 ( n14688,n15875,n15609 );
   nor U15896 ( n15879,n10801,n14689 );
   nand U15897 ( n14689,n15875,n15881 );
   nand U15898 ( n15868,n15882,n15883 );
   nor U15899 ( n15883,n15884,n15885 );
   nor U15900 ( n15885,n14900,n14695 );
   nand U15901 ( n14695,n15875,n15886 );
   nor U15902 ( n15884,n14896,n14697 );
   nand U15903 ( n14697,n15875,n15887 );
   nor U15904 ( n15882,n15888,n15889 );
   nor U15905 ( n15889,n14897,n14701 );
   nand U15906 ( n14701,n15875,n15607 );
   nor U15907 ( n15888,n14890,n14703 );
   nand U15908 ( n14703,n15875,n15832 );
   nor U15909 ( n15866,n15890,n15891 );
   nand U15910 ( n15891,n15892,n15893 );
   nor U15911 ( n15893,n15894,n15895 );
   nor U15912 ( n15895,n14868,n14711 );
   nand U15913 ( n14711,n15832,n15896 );
   nor U15914 ( n15894,n14869,n14713 );
   nand U15915 ( n14713,n15897,n15620 );
   nor U15916 ( n15892,n15898,n15899 );
   nor U15917 ( n15899,n14864,n14717 );
   nand U15918 ( n14717,n15897,n15623 );
   nor U15919 ( n15897,instqueuerd_addr_reg_2_,n15875 );
   nor U15920 ( n15898,n14865,n14719 );
   nand U15921 ( n14719,n15609,n15896 );
   nand U15922 ( n15890,n15900,n15901 );
   nor U15923 ( n15901,n15902,n15903 );
   nor U15924 ( n15903,n14878,n14725 );
   nand U15925 ( n14725,n15881,n15896 );
   nor U15926 ( n15902,n14879,n14727 );
   nand U15927 ( n14727,n15886,n15896 );
   nor U15928 ( n15900,n15904,n15905 );
   nor U15929 ( n15905,n14874,n14731 );
   nand U15930 ( n14731,n15887,n15896 );
   nor U15931 ( n15904,n14875,n14733 );
   nand U15932 ( n14733,n15607,n15896 );
   not U15933 ( n15896,n15875 );
   nor U15934 ( n15875,n15906,n15652 );
   nand U15935 ( n14572,n15907,n15908 );
   nand U15936 ( n15908,n10877,state2_reg_0_ );
   not U15937 ( n10877,n9365 );
   nand U15938 ( n9365,n15909,n8757 );
   and U15939 ( n15909,n10818,n9367 );
   nand U15940 ( n15907,n12994,n9367 );
   nor U15941 ( n9367,n10881,n10798 );
   nand U15942 ( n10881,n15910,n12874 );
   not U15943 ( n12874,n11722 );
   nand U15944 ( n11722,n11679,n10768 );
   nor U15945 ( n15910,n11708,n11661 );
   nor U15946 ( n15655,n15911,n15912 );
   nor U15947 ( n15912,n14040,n12776 );
   not U15948 ( n12776,eax_reg_28_ );
   nand U15949 ( n14040,n11661,state2_reg_2_ );
   not U15950 ( n11661,n10745 );
   nor U15951 ( n15911,n8804,n12265 );
   not U15952 ( n13340,n13314 );
   nand U15953 ( n13314,n15913,state2_reg_1_ );
   nor U15954 ( n15913,n13959,n12461 );
   xor U15955 ( n12461,phyaddrpointer_reg_31_,n14734 );
   nand U15956 ( n14734,phyaddrpointer_reg_30_,n14736 );
   nor U15957 ( n14736,n14745,n12282 );
   not U15958 ( n12282,phyaddrpointer_reg_29_ );
   or U15959 ( n14745,n12265,n14458 );
   or U15960 ( n14458,n12242,n14460 );
   or U15961 ( n14460,n12226,n14471 );
   or U15962 ( n14471,n12207,n14625 );
   or U15963 ( n14625,n12179,n14626 );
   or U15964 ( n14626,n12162,n14566 );
   nand U15965 ( n14566,n15914,phyaddrpointer_reg_22_ );
   nor U15966 ( n15914,n12123,n14487 );
   nand U15967 ( n14487,n15915,phyaddrpointer_reg_20_ );
   nor U15968 ( n15915,n12088,n13989 );
   not U15969 ( n13989,n14489 );
   nor U15970 ( n14489,n12069,n14380 );
   or U15971 ( n14380,n12055,n14337 );
   or U15972 ( n14337,n12039,n14328 );
   or U15973 ( n14328,n12024,n14320 );
   nand U15974 ( n14320,n15916,phyaddrpointer_reg_14_ );
   nor U15975 ( n15916,n11994,n14297 );
   nand U15976 ( n14297,n15917,phyaddrpointer_reg_12_ );
   nor U15977 ( n15917,n11959,n14250 );
   nand U15978 ( n14250,n15918,phyaddrpointer_reg_10_ );
   nor U15979 ( n15918,n11923,n14258 );
   nand U15980 ( n14258,n15919,phyaddrpointer_reg_8_ );
   nor U15981 ( n15919,n11884,n14211 );
   nand U15982 ( n14211,n15920,phyaddrpointer_reg_6_ );
   nor U15983 ( n15920,n11853,n14087 );
   nand U15984 ( n14087,n15921,phyaddrpointer_reg_4_ );
   nor U15985 ( n15921,n11817,n14149 );
   nand U15986 ( n14149,phyaddrpointer_reg_2_,phyaddrpointer_reg_1_ );
   not U15987 ( n11817,phyaddrpointer_reg_3_ );
   not U15988 ( n11853,phyaddrpointer_reg_5_ );
   not U15989 ( n11884,phyaddrpointer_reg_7_ );
   not U15990 ( n11923,phyaddrpointer_reg_9_ );
   not U15991 ( n11959,phyaddrpointer_reg_11_ );
   not U15992 ( n11994,phyaddrpointer_reg_13_ );
   not U15993 ( n12024,phyaddrpointer_reg_15_ );
   not U15994 ( n12039,phyaddrpointer_reg_16_ );
   not U15995 ( n12055,phyaddrpointer_reg_17_ );
   not U15996 ( n12069,phyaddrpointer_reg_18_ );
   not U15997 ( n12088,phyaddrpointer_reg_19_ );
   not U15998 ( n12123,phyaddrpointer_reg_21_ );
   not U15999 ( n12162,phyaddrpointer_reg_23_ );
   not U16000 ( n12179,phyaddrpointer_reg_24_ );
   not U16001 ( n12207,phyaddrpointer_reg_25_ );
   not U16002 ( n12226,phyaddrpointer_reg_26_ );
   not U16003 ( n12242,phyaddrpointer_reg_27_ );
   not U16004 ( n12265,phyaddrpointer_reg_28_ );
   nand U16005 ( n13972,n8824,n13150 );
   not U16006 ( n13150,n11705 );
   xor U16007 ( n11705,n15922,n15923 );
   nand U16008 ( n15923,n13956,n13957 );
   xor U16009 ( n13957,n8757,n15924 );
   nand U16010 ( n15924,n15925,n15926 );
   nand U16011 ( n15926,ebx_reg_30_,n8725 );
   nand U16012 ( n15925,instaddrpointer_reg_30_,n8818 );
   nor U16013 ( n13956,n13878,n13902 );
   xor U16014 ( n13902,n8759,n15928 );
   nand U16015 ( n15928,n15929,n15930 );
   nand U16016 ( n15930,ebx_reg_29_,n8725 );
   nand U16017 ( n15929,instaddrpointer_reg_29_,n13197 );
   or U16018 ( n13878,n13880,n13879 );
   xor U16019 ( n13879,n8761,n15931 );
   nand U16020 ( n15931,n15932,n15933 );
   nand U16021 ( n15933,ebx_reg_28_,n15927 );
   nand U16022 ( n15932,instaddrpointer_reg_28_,n8818 );
   or U16023 ( n13880,n13824,n13850 );
   xor U16024 ( n13850,n15934,n8759 );
   nand U16025 ( n15934,n15935,n15936 );
   nand U16026 ( n15936,ebx_reg_27_,n8725 );
   nand U16027 ( n15935,instaddrpointer_reg_27_,n8818 );
   or U16028 ( n13824,n13826,n13825 );
   xor U16029 ( n13825,n8760,n15937 );
   nand U16030 ( n15937,n15938,n15939 );
   nand U16031 ( n15939,ebx_reg_26_,n15927 );
   nand U16032 ( n15938,instaddrpointer_reg_26_,n13197 );
   or U16033 ( n13826,n13780,n13800 );
   xor U16034 ( n13800,n8761,n15940 );
   nand U16035 ( n15940,n15941,n15942 );
   nand U16036 ( n15942,ebx_reg_25_,n15927 );
   nand U16037 ( n15941,instaddrpointer_reg_25_,n8818 );
   or U16038 ( n13780,n13782,n13781 );
   xor U16039 ( n13781,n8759,n15943 );
   nand U16040 ( n15943,n15944,n15945 );
   nand U16041 ( n15945,ebx_reg_24_,n15927 );
   nand U16042 ( n15944,instaddrpointer_reg_24_,n8818 );
   or U16043 ( n13782,n13730,n13750 );
   xor U16044 ( n13750,n8758,n15946 );
   nand U16045 ( n15946,n15947,n15948 );
   nand U16046 ( n15948,ebx_reg_23_,n15927 );
   nand U16047 ( n15947,instaddrpointer_reg_23_,n8818 );
   or U16048 ( n13730,n13732,n13731 );
   xor U16049 ( n13731,n8761,n15949 );
   nand U16050 ( n15949,n15950,n15951 );
   nand U16051 ( n15951,ebx_reg_22_,n15927 );
   nand U16052 ( n15950,instaddrpointer_reg_22_,n13197 );
   or U16053 ( n13732,n13682,n13702 );
   xor U16054 ( n13702,n8758,n15952 );
   nand U16055 ( n15952,n15953,n15954 );
   nand U16056 ( n15954,ebx_reg_21_,n15927 );
   nand U16057 ( n15953,instaddrpointer_reg_21_,n13197 );
   or U16058 ( n13682,n13684,n13683 );
   xor U16059 ( n13683,n8758,n15955 );
   nand U16060 ( n15955,n15956,n15957 );
   nand U16061 ( n15957,ebx_reg_20_,n15927 );
   nand U16062 ( n15956,instaddrpointer_reg_20_,n13197 );
   or U16063 ( n13684,n13631,n13654 );
   xor U16064 ( n13654,n8760,n15958 );
   nand U16065 ( n15958,n15959,n15960 );
   nand U16066 ( n15960,ebx_reg_19_,n15927 );
   nand U16067 ( n15959,instaddrpointer_reg_19_,n13197 );
   or U16068 ( n13631,n13633,n13632 );
   xor U16069 ( n13632,n8760,n15961 );
   nand U16070 ( n15961,n15962,n15963 );
   nand U16071 ( n15963,ebx_reg_18_,n15927 );
   nand U16072 ( n15962,instaddrpointer_reg_18_,n13197 );
   or U16073 ( n13633,n13579,n13606 );
   xor U16074 ( n13606,n8761,n15964 );
   nand U16075 ( n15964,n15965,n15966 );
   nand U16076 ( n15966,ebx_reg_17_,n15927 );
   nand U16077 ( n15965,instaddrpointer_reg_17_,n13197 );
   or U16078 ( n13579,n13581,n13580 );
   xor U16079 ( n13580,n8760,n15967 );
   nand U16080 ( n15967,n15968,n15969 );
   nand U16081 ( n15969,ebx_reg_16_,n15927 );
   nand U16082 ( n15968,instaddrpointer_reg_16_,n8818 );
   or U16083 ( n13581,n13529,n13550 );
   xor U16084 ( n13550,n8759,n15970 );
   nand U16085 ( n15970,n15971,n15972 );
   nand U16086 ( n15972,ebx_reg_15_,n15927 );
   nand U16087 ( n15971,instaddrpointer_reg_15_,n13197 );
   or U16088 ( n13529,n13531,n13530 );
   xor U16089 ( n13530,n8758,n15973 );
   nand U16090 ( n15973,n15974,n15975 );
   nand U16091 ( n15975,ebx_reg_14_,n15927 );
   nand U16092 ( n15974,instaddrpointer_reg_14_,n13197 );
   or U16093 ( n13531,n13482,n13504 );
   xor U16094 ( n13504,n8759,n15976 );
   nand U16095 ( n15976,n15977,n15978 );
   nand U16096 ( n15978,ebx_reg_13_,n15927 );
   nand U16097 ( n15977,instaddrpointer_reg_13_,n13197 );
   or U16098 ( n13482,n13484,n13483 );
   xor U16099 ( n13483,n8760,n15979 );
   nand U16100 ( n15979,n15980,n15981 );
   nand U16101 ( n15981,ebx_reg_12_,n15927 );
   nand U16102 ( n15980,instaddrpointer_reg_12_,n13197 );
   or U16103 ( n13484,n13434,n13455 );
   xor U16104 ( n13455,n8759,n15982 );
   nand U16105 ( n15982,n15983,n15984 );
   nand U16106 ( n15984,ebx_reg_11_,n15927 );
   nand U16107 ( n15983,instaddrpointer_reg_11_,n8818 );
   or U16108 ( n13434,n13436,n13435 );
   xor U16109 ( n13435,n8758,n15985 );
   nand U16110 ( n15985,n15986,n15987 );
   nand U16111 ( n15987,ebx_reg_10_,n15927 );
   nand U16112 ( n15986,instaddrpointer_reg_10_,n13197 );
   or U16113 ( n13436,n13388,n13409 );
   xor U16114 ( n13409,n8760,n15988 );
   nand U16115 ( n15988,n15989,n15990 );
   nand U16116 ( n15990,ebx_reg_9_,n8725 );
   nand U16117 ( n15989,instaddrpointer_reg_9_,n13197 );
   or U16118 ( n13388,n13390,n13389 );
   xor U16119 ( n13389,n8760,n15991 );
   nand U16120 ( n15991,n15992,n15993 );
   nand U16121 ( n15993,ebx_reg_8_,n8725 );
   nand U16122 ( n15992,instaddrpointer_reg_8_,n13197 );
   or U16123 ( n13390,n13336,n13360 );
   xor U16124 ( n13360,n8761,n15994 );
   nand U16125 ( n15994,n15995,n15996 );
   nand U16126 ( n15996,ebx_reg_7_,n8725 );
   nand U16127 ( n15995,instaddrpointer_reg_7_,n13197 );
   or U16128 ( n13336,n13338,n13337 );
   xor U16129 ( n13337,n8758,n15997 );
   nand U16130 ( n15997,n15998,n15999 );
   nand U16131 ( n15999,ebx_reg_6_,n8725 );
   nand U16132 ( n15998,instaddrpointer_reg_6_,n13197 );
   or U16133 ( n13338,n13275,n13304 );
   xor U16134 ( n13304,n8758,n16000 );
   nand U16135 ( n16000,n16001,n16002 );
   nand U16136 ( n16002,ebx_reg_5_,n8725 );
   nand U16137 ( n16001,instaddrpointer_reg_5_,n13197 );
   or U16138 ( n13275,n13277,n13276 );
   xor U16139 ( n13276,n8761,n16003 );
   nand U16140 ( n16003,n16004,n16005 );
   nand U16141 ( n16005,ebx_reg_4_,n8725 );
   nand U16142 ( n16004,instaddrpointer_reg_4_,n13197 );
   or U16143 ( n13277,n13253,n13254 );
   xor U16144 ( n13254,n8761,n16006 );
   nand U16145 ( n16006,n16007,n16008 );
   nand U16146 ( n16008,ebx_reg_3_,n8725 );
   nand U16147 ( n16007,instaddrpointer_reg_3_,n13197 );
   or U16148 ( n13253,n13229,n13228 );
   xor U16149 ( n13228,n8759,n16009 );
   nand U16150 ( n16009,n16010,n16011 );
   nand U16151 ( n16011,ebx_reg_2_,n8725 );
   nand U16152 ( n16010,instaddrpointer_reg_2_,n8818 );
   not U16153 ( n13197,n16012 );
   nand U16154 ( n13229,n16013,n16014 );
   nand U16155 ( n16014,n16015,n16012 );
   or U16156 ( n16015,n13195,n13198 );
   nand U16157 ( n16013,n13195,n13198 );
   nand U16158 ( n13198,n13180,n8725 );
   xor U16159 ( n13180,n16016,n8759 );
   nor U16160 ( n16016,n16017,n16018 );
   nor U16161 ( n16018,n8965,n16012 );
   not U16162 ( n8965,instaddrpointer_reg_0_ );
   nor U16163 ( n16017,n13179,n13182 );
   not U16164 ( n13182,ebx_reg_0_ );
   xor U16165 ( n13195,n16019,n8757 );
   nor U16166 ( n16019,n16020,n16021 );
   nor U16167 ( n16021,n8996,n16012 );
   not U16168 ( n8996,instaddrpointer_reg_1_ );
   and U16169 ( n16020,n15927,ebx_reg_1_ );
   nor U16170 ( n15922,n8757,n16022 );
   nor U16171 ( n16022,n16023,n16024 );
   nor U16172 ( n16024,n8997,n16012 );
   nand U16173 ( n16012,n12992,n16025 );
   nand U16174 ( n16025,n15213,n10818 );
   not U16175 ( n8997,instaddrpointer_reg_31_ );
   nor U16176 ( n16023,n13179,n16026 );
   not U16177 ( n13179,n15927 );
   nand U16178 ( n15927,n8761,n11671 );
   nand U16179 ( n11671,n11631,n10818 );
   and U16180 ( n13177,n16027,n16028 );
   nor U16181 ( n16028,n16029,n12992 );
   and U16182 ( n16027,ebx_reg_31_,n13279 );
   nor U16183 ( n13970,n12466,n13164 );
   nand U16184 ( n13164,state2_reg_3_,n8774 );
   not U16185 ( n12466,phyaddrpointer_reg_31_ );
   nor U16186 ( n13968,n16030,n16031 );
   nand U16187 ( n16031,n16032,n16033 );
   nand U16188 ( n16033,reip_reg_31_,n16034 );
   nand U16189 ( n16034,n16035,n16036 );
   nand U16190 ( n16036,n8746,n9047 );
   not U16191 ( n9047,reip_reg_30_ );
   not U16192 ( n16035,n13966 );
   nand U16193 ( n13966,n13910,n16037 );
   nand U16194 ( n16037,n8746,n9052 );
   not U16195 ( n9052,reip_reg_29_ );
   nor U16196 ( n13910,n13887,n16038 );
   nor U16197 ( n16038,n13168,reip_reg_28_ );
   nand U16198 ( n13887,n13167,n16039 );
   nand U16199 ( n16039,n8747,n13889 );
   not U16200 ( n13889,n16040 );
   nand U16201 ( n16032,n16041,n9045 );
   not U16202 ( n9045,reip_reg_31_ );
   nor U16203 ( n16041,n13909,n16042 );
   nand U16204 ( n16042,reip_reg_29_,reip_reg_30_ );
   nand U16205 ( n13909,n16043,n16040 );
   nor U16206 ( n16040,n16044,n13835 );
   nand U16207 ( n13835,n16045,n13813 );
   nor U16208 ( n13813,n16046,n13741 );
   nand U16209 ( n13741,n16047,n13715 );
   nor U16210 ( n13715,n16048,n13647 );
   nand U16211 ( n13647,n16049,n13622 );
   nor U16212 ( n13622,n16050,n13543 );
   nand U16213 ( n13543,n16051,n13520 );
   nor U16214 ( n13520,n16052,n13448 );
   nand U16215 ( n13448,n16053,n13425 );
   nor U16216 ( n13425,n16054,n13353 );
   nand U16217 ( n13353,n16055,n13293 );
   not U16218 ( n13293,n13325 );
   nand U16219 ( n13325,n16056,reip_reg_2_ );
   nor U16220 ( n16056,n9192,n9182 );
   not U16221 ( n9182,reip_reg_3_ );
   nor U16222 ( n16055,n9172,n9177 );
   not U16223 ( n9177,reip_reg_4_ );
   not U16224 ( n9172,reip_reg_5_ );
   nand U16225 ( n16054,reip_reg_7_,reip_reg_6_ );
   nor U16226 ( n16053,n9152,n9157 );
   not U16227 ( n9157,reip_reg_8_ );
   not U16228 ( n9152,reip_reg_9_ );
   nand U16229 ( n16052,reip_reg_11_,reip_reg_10_ );
   nor U16230 ( n16051,n9132,n9137 );
   not U16231 ( n9137,reip_reg_12_ );
   not U16232 ( n9132,reip_reg_13_ );
   nand U16233 ( n16050,reip_reg_15_,reip_reg_14_ );
   nor U16234 ( n16049,n9112,n9117 );
   not U16235 ( n9117,reip_reg_16_ );
   not U16236 ( n9112,reip_reg_17_ );
   nand U16237 ( n16048,reip_reg_19_,reip_reg_18_ );
   nor U16238 ( n16047,n9092,n9097 );
   not U16239 ( n9097,reip_reg_20_ );
   not U16240 ( n9092,reip_reg_21_ );
   nand U16241 ( n16046,reip_reg_23_,reip_reg_22_ );
   nor U16242 ( n16045,n9072,n9077 );
   not U16243 ( n9077,reip_reg_24_ );
   not U16244 ( n9072,reip_reg_25_ );
   nand U16245 ( n16044,reip_reg_27_,reip_reg_26_ );
   nor U16246 ( n16043,n9057,n8782 );
   nand U16247 ( n13168,n16057,n13279 );
   nor U16248 ( n16057,n16058,n16059 );
   nor U16249 ( n16058,n16060,n15211 );
   nor U16250 ( n16060,n8867,n12359 );
   not U16251 ( n9057,reip_reg_28_ );
   nor U16252 ( n16030,n16026,n13183 );
   nand U16253 ( n13183,n13279,n16061 );
   nand U16254 ( n16061,n16062,n16063 );
   nand U16255 ( n16063,n16064,n15211 );
   nor U16256 ( n16064,ebx_reg_31_,n16029 );
   nand U16257 ( n16062,n8874,n9310 );
   nand U16258 ( n9310,n16029,n8876 );
   not U16259 ( n16029,n16059 );
   nand U16260 ( n16059,n10838,n8862 );
   nor U16261 ( n13279,n8789,n13959 );
   not U16262 ( n13959,n13167 );
   nand U16263 ( n13167,n16065,n16066 );
   nor U16264 ( n16066,n16067,n9283 );
   and U16265 ( n9283,n16068,n8830 );
   nor U16266 ( n16068,state2_reg_0_,n8948 );
   not U16267 ( n16067,n9293 );
   nand U16268 ( n9293,n16069,n8868 );
   nor U16269 ( n8868,state2_reg_1_,state2_reg_2_ );
   nor U16270 ( n16069,n8863,n9018 );
   nor U16271 ( n16065,n8842,n11734 );
   nor U16272 ( n11734,state2_reg_2_,n12469 );
   nand U16273 ( n12469,n8960,n8821 );
   not U16274 ( n8960,n8981 );
   nand U16275 ( n8981,n8948,n9018 );
   not U16276 ( n9018,state2_reg_3_ );
   and U16277 ( n8842,n9275,n16070 );
   nand U16278 ( n16070,n16071,n16072 );
   nand U16279 ( n16072,n15194,n11741 );
   nor U16280 ( n15194,n10889,n8863 );
   nand U16281 ( n10889,n8845,n16073 );
   nor U16282 ( n16071,n16074,n16075 );
   nor U16283 ( n16075,n9350,n16076 );
   nand U16284 ( n16076,state2_reg_0_,n9384 );
   nand U16285 ( n9350,n13278,n16073 );
   nor U16286 ( n13278,n10906,n10818 );
   not U16287 ( n16026,ebx_reg_31_ );
   nor U16288 ( n16077,n16079,n16080 );
   nor U16289 ( n16080,n8888,n16081 );
   or U16290 ( n16081,datawidth_reg_1_,reip_reg_1_ );
   and U16291 ( n16079,n8888,byteenable_reg_3_ );
   nand U16292 ( n16083,byteenable_reg_1_,n8888 );
   and U16293 ( n16082,n16078,n8885 );
   not U16294 ( n8885,n8892 );
   nor U16295 ( n8892,n9192,n8888 );
   not U16296 ( n9192,reip_reg_1_ );
   nand U16297 ( n16078,n16084,n16085 );
   nor U16298 ( n16085,reip_reg_0_,datawidth_reg_1_ );
   nor U16299 ( n16084,datawidth_reg_0_,n8888 );
   nand U16300 ( n8888,n16086,n16087 );
   nor U16301 ( n16087,n16088,n16089 );
   nand U16302 ( n16089,n16090,n16091 );
   nor U16303 ( n16091,n16092,n16093 );
   nand U16304 ( n16093,n9264,n9265 );
   not U16305 ( n9265,datawidth_reg_29_ );
   not U16306 ( n9264,datawidth_reg_28_ );
   nand U16307 ( n16092,n9238,n9266 );
   not U16308 ( n9266,datawidth_reg_30_ );
   not U16309 ( n9238,datawidth_reg_2_ );
   nor U16310 ( n16090,n16094,n16095 );
   nand U16311 ( n16095,n9260,n9261 );
   not U16312 ( n9261,datawidth_reg_25_ );
   not U16313 ( n9260,datawidth_reg_24_ );
   nand U16314 ( n16094,n9262,n9263 );
   not U16315 ( n9263,datawidth_reg_27_ );
   not U16316 ( n9262,datawidth_reg_26_ );
   nand U16317 ( n16088,n16096,n16097 );
   nor U16318 ( n16097,n16098,n16099 );
   nand U16319 ( n16099,n9242,n9243 );
   not U16320 ( n9243,datawidth_reg_7_ );
   not U16321 ( n9242,datawidth_reg_6_ );
   nand U16322 ( n16098,n9244,n9245 );
   not U16323 ( n9245,datawidth_reg_9_ );
   not U16324 ( n9244,datawidth_reg_8_ );
   nor U16325 ( n16096,n16100,n16101 );
   nand U16326 ( n16101,n9267,n9239 );
   not U16327 ( n9239,datawidth_reg_3_ );
   not U16328 ( n9267,datawidth_reg_31_ );
   nand U16329 ( n16100,n9240,n9241 );
   not U16330 ( n9241,datawidth_reg_5_ );
   not U16331 ( n9240,datawidth_reg_4_ );
   nor U16332 ( n16086,n16102,n16103 );
   nand U16333 ( n16103,n16104,n16105 );
   nor U16334 ( n16105,n16106,n16107 );
   nand U16335 ( n16107,n9248,n9249 );
   not U16336 ( n9249,datawidth_reg_13_ );
   not U16337 ( n9248,datawidth_reg_12_ );
   nand U16338 ( n16106,n9250,n9251 );
   not U16339 ( n9251,datawidth_reg_15_ );
   not U16340 ( n9250,datawidth_reg_14_ );
   nor U16341 ( n16104,n16108,n16109 );
   nand U16342 ( n16109,n9246,n9247 );
   not U16343 ( n9247,datawidth_reg_11_ );
   not U16344 ( n9246,datawidth_reg_10_ );
   and U16345 ( n16108,datawidth_reg_0_,datawidth_reg_1_ );
   nand U16346 ( n16102,n16110,n16111 );
   nor U16347 ( n16111,n16112,n16113 );
   nand U16348 ( n16113,n9256,n9257 );
   not U16349 ( n9257,datawidth_reg_21_ );
   not U16350 ( n9256,datawidth_reg_20_ );
   nand U16351 ( n16112,n9258,n9259 );
   not U16352 ( n9259,datawidth_reg_23_ );
   not U16353 ( n9258,datawidth_reg_22_ );
   nor U16354 ( n16110,n16114,n16115 );
   nand U16355 ( n16115,n9252,n9253 );
   not U16356 ( n9253,datawidth_reg_17_ );
   not U16357 ( n9252,datawidth_reg_16_ );
   nand U16358 ( n16114,n9254,n9255 );
   not U16359 ( n9255,datawidth_reg_19_ );
   not U16360 ( n9254,datawidth_reg_18_ );
   nand U16361 ( n16116,flush_reg,n8881 );
   not U16362 ( n8881,n8879 );
   nor U16363 ( n8879,n9015,n9369 );
   and U16364 ( n9369,n16117,n16118 );
   nand U16365 ( n16118,n8862,n16119 );
   nand U16366 ( n16119,n16120,n8867 );
   not U16367 ( n8867,n8876 );
   nor U16368 ( n8876,n15213,state_reg_0_ );
   nand U16369 ( n15213,n9027,n16121 );
   nand U16370 ( n16121,state_reg_2_,state_reg_1_ );
   nor U16371 ( n16120,n15211,n8845 );
   not U16372 ( n8845,n11632 );
   not U16373 ( n15211,n12992 );
   not U16374 ( n8862,ready_n );
   nand U16375 ( n12470,n16122,n16123 );
   nor U16376 ( n16123,n9392,n16124 );
   nand U16377 ( n16124,n9384,n8948 );
   nor U16378 ( n16122,n14125,n16125 );
   not U16379 ( n14125,n11710 );
   nor U16380 ( n11710,n11748,n8871 );
   not U16381 ( n8871,state2_reg_2_ );
   nor U16382 ( n16126,n16128,n16129 );
   nor U16383 ( n16129,n10838,n8755 );
   not U16384 ( n9025,n9023 );
   not U16385 ( n10838,statebs16_reg );
   nor U16386 ( n16128,n9023,n9026 );
   not U16387 ( n9026,bs16_n );
   nand U16388 ( n16127,n9031,n9202 );
   not U16389 ( n9031,n9027 );
   nand U16390 ( n9027,n9203,n9208 );
   not U16391 ( n9208,state_reg_2_ );
   nor U16392 ( n16130,n16131,n16132 );
   and U16393 ( n16132,d_c_n_reg,n8742 );
   nor U16394 ( n16131,codefetch_reg,n8741 );
   nand U16395 ( n8848,state_reg_1_,n9202 );
   not U16396 ( n9202,state_reg_0_ );
   nand U16397 ( n16134,codefetch_reg,n16135 );
   nand U16398 ( n16135,n16117,n9287 );
   and U16399 ( n16117,n16136,n16137 );
   nand U16400 ( n16137,n16138,n16139 );
   or U16401 ( n16139,n9388,n9393 );
   not U16402 ( n9393,n9384 );
   nand U16403 ( n16138,n16073,n9391 );
   nor U16404 ( n16136,n11731,n16140 );
   nor U16405 ( n16140,n11741,n11632 );
   nand U16406 ( n11632,n10906,n9391 );
   not U16407 ( n11741,n9380 );
   nor U16408 ( n11731,n9384,n10906 );
   nand U16409 ( n16133,n8843,state2_reg_0_ );
   nand U16410 ( n16141,ads_n_reg,state_reg_0_ );
   nor U16411 ( n9023,n16142,n9228 );
   nor U16412 ( n9228,state_reg_0_,state_reg_1_ );
   and U16413 ( n16142,n16143,state_reg_0_ );
   nor U16414 ( n16143,state_reg_2_,n9203 );
   not U16415 ( n9203,state_reg_1_ );
   nand U16416 ( n16145,memoryfetch_reg,n16146 );
   nand U16417 ( n16146,n16147,n16148 );
   nor U16418 ( n16148,n9380,n12996 );
   nand U16419 ( n9380,n16149,n16150 );
   nand U16420 ( n16150,n16151,n16152 );
   nor U16421 ( n16152,n16153,n16154 );
   nor U16422 ( n16151,n16155,n16156 );
   not U16423 ( n16156,n16157 );
   nor U16424 ( n16147,n15063,n13002 );
   not U16425 ( n13002,n16073 );
   nor U16426 ( n16073,n11726,n11627 );
   nand U16427 ( n11726,n9390,n11631 );
   not U16428 ( n11631,n10788 );
   nor U16429 ( n9390,n16158,n11748 );
   nand U16430 ( n11748,n10745,n10758 );
   nand U16431 ( n16158,n10768,n11708 );
   nor U16432 ( n16144,n16074,n8843 );
   and U16433 ( n8843,n8857,n8948 );
   nor U16434 ( n8857,state2_reg_2_,state2_reg_3_ );
   nor U16435 ( n16074,n11745,n9388 );
   nand U16436 ( n9388,n10914,n10818 );
   not U16437 ( n10914,n10890 );
   nand U16438 ( n10890,n16159,n16160 );
   nor U16439 ( n16160,n15161,n10778 );
   nand U16440 ( n15161,n11679,n10745 );
   nand U16441 ( n10745,n16161,n16162 );
   nor U16442 ( n16162,n16163,n16164 );
   nand U16443 ( n16164,n16165,n16166 );
   nor U16444 ( n16166,n16167,n16168 );
   nor U16445 ( n16168,n16169,n14730 );
   not U16446 ( n14730,instqueue_reg_10__7_ );
   nor U16447 ( n16167,n16170,n14724 );
   not U16448 ( n14724,instqueue_reg_8__7_ );
   nor U16449 ( n16165,n16171,n16172 );
   nor U16450 ( n16172,n16173,n14718 );
   not U16451 ( n14718,instqueue_reg_15__7_ );
   nor U16452 ( n16171,n16174,n14716 );
   not U16453 ( n14716,instqueue_reg_14__7_ );
   nand U16454 ( n16163,n16175,n16176 );
   nor U16455 ( n16176,n16177,n16178 );
   nor U16456 ( n16178,n16179,n10750 );
   not U16457 ( n10750,instqueue_reg_0__7_ );
   nor U16458 ( n16177,n16180,n14700 );
   not U16459 ( n14700,instqueue_reg_3__7_ );
   nor U16460 ( n16175,n16181,n16182 );
   nor U16461 ( n16182,n16183,n14710 );
   not U16462 ( n14710,instqueue_reg_12__7_ );
   nor U16463 ( n16181,n16184,n14732 );
   not U16464 ( n14732,instqueue_reg_11__7_ );
   nor U16465 ( n16161,n16185,n16186 );
   nand U16466 ( n16186,n16187,n16188 );
   nor U16467 ( n16188,n16189,n16190 );
   nor U16468 ( n16190,n16191,n14683 );
   not U16469 ( n14683,instqueue_reg_6__7_ );
   nor U16470 ( n16189,n16192,n14681 );
   not U16471 ( n14681,instqueue_reg_5__7_ );
   nor U16472 ( n16187,n16193,n16194 );
   nor U16473 ( n16194,n16195,n14702 );
   not U16474 ( n14702,instqueue_reg_4__7_ );
   nor U16475 ( n16193,n16196,n14696 );
   not U16476 ( n14696,instqueue_reg_2__7_ );
   nand U16477 ( n16185,n16197,n16198 );
   nor U16478 ( n16198,n16199,n16200 );
   nor U16479 ( n16200,n16201,n14726 );
   not U16480 ( n14726,instqueue_reg_9__7_ );
   nor U16481 ( n16199,n16202,n14712 );
   not U16482 ( n14712,instqueue_reg_13__7_ );
   nor U16483 ( n16197,n16203,n16204 );
   nor U16484 ( n16204,n16205,n14694 );
   not U16485 ( n14694,instqueue_reg_1__7_ );
   nor U16486 ( n16203,n15605,n14687 );
   not U16487 ( n14687,instqueue_reg_7__7_ );
   not U16488 ( n11679,n10758 );
   nand U16489 ( n10758,n16206,n16207 );
   nor U16490 ( n16207,n16208,n16209 );
   nand U16491 ( n16209,n16210,n16211 );
   nor U16492 ( n16211,n16212,n16213 );
   nor U16493 ( n16213,n16169,n14792 );
   not U16494 ( n14792,instqueue_reg_10__6_ );
   nor U16495 ( n16212,n16170,n14788 );
   not U16496 ( n14788,instqueue_reg_8__6_ );
   nor U16497 ( n16210,n16214,n16215 );
   nor U16498 ( n16215,n16173,n14783 );
   not U16499 ( n14783,instqueue_reg_15__6_ );
   nor U16500 ( n16214,n16174,n14782 );
   not U16501 ( n14782,instqueue_reg_14__6_ );
   nand U16502 ( n16208,n16216,n16217 );
   nor U16503 ( n16217,n16218,n16219 );
   nor U16504 ( n16219,n16179,n10761 );
   not U16505 ( n10761,instqueue_reg_0__6_ );
   nor U16506 ( n16218,n16220,n14770 );
   not U16507 ( n14770,instqueue_reg_3__6_ );
   nor U16508 ( n16216,n16221,n16222 );
   nor U16509 ( n16222,n16183,n14778 );
   not U16510 ( n14778,instqueue_reg_12__6_ );
   nor U16511 ( n16221,n16184,n14793 );
   not U16512 ( n14793,instqueue_reg_11__6_ );
   nor U16513 ( n16206,n16223,n16224 );
   nand U16514 ( n16224,n16225,n16226 );
   nor U16515 ( n16226,n16227,n16228 );
   nor U16516 ( n16228,n16191,n14758 );
   not U16517 ( n14758,instqueue_reg_6__6_ );
   nor U16518 ( n16227,n16192,n14757 );
   not U16519 ( n14757,instqueue_reg_5__6_ );
   nor U16520 ( n16225,n16229,n16230 );
   nor U16521 ( n16230,n16195,n14771 );
   not U16522 ( n14771,instqueue_reg_4__6_ );
   nor U16523 ( n16229,n16196,n14767 );
   not U16524 ( n14767,instqueue_reg_2__6_ );
   nand U16525 ( n16223,n16231,n16232 );
   nor U16526 ( n16232,n16233,n16234 );
   nor U16527 ( n16234,n16201,n14789 );
   not U16528 ( n14789,instqueue_reg_9__6_ );
   nor U16529 ( n16233,n16202,n14779 );
   not U16530 ( n14779,instqueue_reg_13__6_ );
   nor U16531 ( n16231,n16235,n16236 );
   nor U16532 ( n16236,n16205,n14766 );
   not U16533 ( n14766,instqueue_reg_1__6_ );
   nor U16534 ( n16235,n15605,n14761 );
   not U16535 ( n14761,instqueue_reg_7__6_ );
   nor U16536 ( n16159,n10768,n9392 );
   nand U16537 ( n9392,n11627,n10788 );
   nand U16538 ( n10788,n16237,n16238 );
   nor U16539 ( n16238,n16239,n16240 );
   nand U16540 ( n16240,n16241,n16242 );
   nor U16541 ( n16242,n16243,n16244 );
   nor U16542 ( n16244,n16169,n15258 );
   not U16543 ( n15258,instqueue_reg_10__3_ );
   nor U16544 ( n16243,n16170,n15278 );
   not U16545 ( n15278,instqueue_reg_8__3_ );
   nor U16546 ( n16241,n16245,n16246 );
   nor U16547 ( n16246,n16173,n15270 );
   not U16548 ( n15270,instqueue_reg_15__3_ );
   nor U16549 ( n16245,n16174,n15269 );
   not U16550 ( n15269,instqueue_reg_14__3_ );
   nand U16551 ( n16239,n16247,n16248 );
   nor U16552 ( n16248,n16249,n16250 );
   nor U16553 ( n16250,n16179,n10791 );
   not U16554 ( n10791,instqueue_reg_0__3_ );
   nor U16555 ( n16249,n16180,n15247 );
   not U16556 ( n15247,instqueue_reg_3__3_ );
   nor U16557 ( n16247,n16251,n16252 );
   nor U16558 ( n16252,n16183,n15279 );
   not U16559 ( n15279,instqueue_reg_12__3_ );
   nor U16560 ( n16251,n16184,n15265 );
   not U16561 ( n15265,instqueue_reg_11__3_ );
   nor U16562 ( n16237,n16253,n16254 );
   nand U16563 ( n16254,n16255,n16256 );
   nor U16564 ( n16256,n16257,n16258 );
   nor U16565 ( n16258,n16191,n15253 );
   not U16566 ( n15253,instqueue_reg_6__3_ );
   nor U16567 ( n16257,n16192,n15248 );
   not U16568 ( n15248,instqueue_reg_5__3_ );
   nor U16569 ( n16255,n16259,n16260 );
   nor U16570 ( n16260,n16195,n15275 );
   not U16571 ( n15275,instqueue_reg_4__3_ );
   nor U16572 ( n16259,n16196,n15244 );
   not U16573 ( n15244,instqueue_reg_2__3_ );
   nand U16574 ( n16253,n16261,n16262 );
   nor U16575 ( n16262,n16263,n16264 );
   nor U16576 ( n16264,n16201,n15257 );
   not U16577 ( n15257,instqueue_reg_9__3_ );
   nor U16578 ( n16263,n16202,n15266 );
   not U16579 ( n15266,instqueue_reg_13__3_ );
   nor U16580 ( n16261,n16265,n16266 );
   nor U16581 ( n16266,n16205,n15243 );
   not U16582 ( n15243,instqueue_reg_1__3_ );
   nor U16583 ( n16265,n15605,n15254 );
   not U16584 ( n15254,instqueue_reg_7__3_ );
   not U16585 ( n11627,n10798 );
   nand U16586 ( n10798,n16267,n16268 );
   nor U16587 ( n16268,n16269,n16270 );
   nand U16588 ( n16270,n16271,n16272 );
   nor U16589 ( n16272,n16273,n16274 );
   nor U16590 ( n16274,n16169,n14874 );
   not U16591 ( n14874,instqueue_reg_10__2_ );
   nor U16592 ( n16273,n16170,n14878 );
   not U16593 ( n14878,instqueue_reg_8__2_ );
   nor U16594 ( n16271,n16275,n16276 );
   nor U16595 ( n16276,n16173,n14865 );
   not U16596 ( n14865,instqueue_reg_15__2_ );
   nor U16597 ( n16275,n16174,n14864 );
   not U16598 ( n14864,instqueue_reg_14__2_ );
   nand U16599 ( n16269,n16277,n16278 );
   nor U16600 ( n16278,n16279,n16280 );
   nor U16601 ( n16280,n16179,n10801 );
   not U16602 ( n10801,instqueue_reg_0__2_ );
   nor U16603 ( n16279,n16180,n14897 );
   not U16604 ( n14897,instqueue_reg_3__2_ );
   nor U16605 ( n16277,n16281,n16282 );
   nor U16606 ( n16282,n16183,n14868 );
   not U16607 ( n14868,instqueue_reg_12__2_ );
   nor U16608 ( n16281,n16184,n14875 );
   not U16609 ( n14875,instqueue_reg_11__2_ );
   nor U16610 ( n16267,n16283,n16284 );
   nand U16611 ( n16284,n16285,n16286 );
   nor U16612 ( n16286,n16287,n16288 );
   nor U16613 ( n16288,n16191,n14886 );
   not U16614 ( n14886,instqueue_reg_6__2_ );
   nor U16615 ( n16287,n16192,n14891 );
   not U16616 ( n14891,instqueue_reg_5__2_ );
   nor U16617 ( n16285,n16289,n16290 );
   nor U16618 ( n16290,n16195,n14890 );
   not U16619 ( n14890,instqueue_reg_4__2_ );
   nor U16620 ( n16289,n16196,n14896 );
   not U16621 ( n14896,instqueue_reg_2__2_ );
   nand U16622 ( n16283,n16291,n16292 );
   nor U16623 ( n16292,n16293,n16294 );
   nor U16624 ( n16294,n16201,n14879 );
   not U16625 ( n14879,instqueue_reg_9__2_ );
   nor U16626 ( n16293,n16202,n14869 );
   not U16627 ( n14869,instqueue_reg_13__2_ );
   nor U16628 ( n16291,n16295,n16296 );
   nor U16629 ( n16296,n16205,n14900 );
   not U16630 ( n14900,instqueue_reg_1__2_ );
   nor U16631 ( n16295,n15605,n14887 );
   not U16632 ( n14887,instqueue_reg_7__2_ );
   nand U16633 ( n11745,n9287,n9384 );
   nand U16634 ( n9384,n16297,n16298 );
   nand U16635 ( n16298,n16299,n16300 );
   nand U16636 ( n16300,n16301,n16302 );
   nand U16637 ( n16302,n16303,n16304 );
   nand U16638 ( n16303,n16305,n16306 );
   nand U16639 ( n16306,n16154,n11732 );
   nand U16640 ( n16305,n16307,n16153 );
   nand U16641 ( n16301,n16308,n16309 );
   nand U16642 ( n16309,n16310,n16311 );
   nor U16643 ( n16308,n16312,n16313 );
   nor U16644 ( n16313,n16314,n16315 );
   nor U16645 ( n16315,n16316,n16317 );
   and U16646 ( n16317,n16318,n16319 );
   nor U16647 ( n16316,n16320,n16321 );
   nor U16648 ( n16321,n16319,n16318 );
   nand U16649 ( n16318,n16322,n16323 );
   nand U16650 ( n16323,n16324,n12341 );
   not U16651 ( n12341,n12383 );
   nand U16652 ( n12383,n10808,n10768 );
   nor U16653 ( n16324,n16325,n11732 );
   nand U16654 ( n16322,n16326,n16327 );
   nor U16655 ( n16326,n16325,n16328 );
   nor U16656 ( n16328,n16329,n16330 );
   and U16657 ( n16325,n16331,n16125 );
   nand U16658 ( n16125,n16332,n15407 );
   not U16659 ( n15407,n16333 );
   nor U16660 ( n16332,n12386,n9391 );
   and U16661 ( n16331,n16330,n16334 );
   and U16662 ( n16330,n16335,n16336 );
   nand U16663 ( n16336,instqueuewr_addr_reg_0_,n8968 );
   nand U16664 ( n16319,n16337,n16338 );
   nor U16665 ( n16338,n12386,n8866 );
   nor U16666 ( n16337,n16339,n16340 );
   nor U16667 ( n16340,n10906,n16333 );
   nor U16668 ( n16339,n16157,n11732 );
   nor U16669 ( n16320,n16329,n16157 );
   xor U16670 ( n16157,n16341,n16335 );
   xor U16671 ( n16341,instqueuewr_addr_reg_1_,instqueuerd_addr_reg_1_ );
   nor U16672 ( n16314,n16310,n16311 );
   nand U16673 ( n16311,n16334,n16342 );
   nand U16674 ( n16342,n16155,n15061 );
   nand U16675 ( n16334,n10906,n16343 );
   or U16676 ( n16343,n10768,n12994 );
   not U16677 ( n10768,n12386 );
   and U16678 ( n16310,n16327,n16344 );
   nand U16679 ( n16344,n16155,n16304 );
   xor U16680 ( n16155,n16345,n16346 );
   xor U16681 ( n16345,instqueuewr_addr_reg_2_,instqueuerd_addr_reg_2_ );
   nand U16682 ( n16327,n15063,n16333 );
   nor U16683 ( n16312,n11732,n16347 );
   nand U16684 ( n16347,n16154,n16329 );
   xor U16685 ( n16154,n16348,n16349 );
   xor U16686 ( n16348,instqueuewr_addr_reg_3_,instqueuerd_addr_reg_3_ );
   nor U16687 ( n16299,n16350,n16351 );
   nor U16688 ( n16351,n16329,n16352 );
   nand U16689 ( n16352,n16353,n11732 );
   not U16690 ( n16329,n16304 );
   nor U16691 ( n16350,n16307,n16304 );
   and U16692 ( n16307,n16354,n16355 );
   nand U16693 ( n16355,n15061,n16153 );
   xor U16694 ( n16153,n16356,n16357 );
   xor U16695 ( n16356,instqueuewr_addr_reg_4_,instqueuerd_addr_reg_4_ );
   not U16696 ( n15061,n11732 );
   nand U16697 ( n16354,instqueuerd_addr_reg_4_,n8821 );
   nand U16698 ( n16297,n16358,n16353 );
   not U16699 ( n16353,n16149 );
   nand U16700 ( n16149,n16359,n16360 );
   nand U16701 ( n16360,instqueuewr_addr_reg_4_,n16361 );
   nand U16702 ( n16361,instqueuerd_addr_reg_4_,n16357 );
   or U16703 ( n16359,n16357,instqueuerd_addr_reg_4_ );
   nand U16704 ( n16357,n16362,n16363 );
   nand U16705 ( n16363,n16364,n9788 );
   not U16706 ( n9788,instqueuewr_addr_reg_3_ );
   or U16707 ( n16364,n16349,instqueuerd_addr_reg_3_ );
   nand U16708 ( n16362,instqueuerd_addr_reg_3_,n16349 );
   nand U16709 ( n16349,n16365,n16366 );
   nand U16710 ( n16366,n16367,n9354 );
   not U16711 ( n9354,instqueuewr_addr_reg_2_ );
   or U16712 ( n16367,n16346,instqueuerd_addr_reg_2_ );
   nand U16713 ( n16365,instqueuerd_addr_reg_2_,n16346 );
   nand U16714 ( n16346,n16368,n16369 );
   nand U16715 ( n16369,n16370,n9356 );
   not U16716 ( n9356,instqueuewr_addr_reg_1_ );
   nand U16717 ( n16370,n9339,n16335 );
   nand U16718 ( n16368,n16371,instqueuerd_addr_reg_1_ );
   not U16719 ( n16371,n16335 );
   nand U16720 ( n16335,instqueuerd_addr_reg_0_,n15188 );
   not U16721 ( n15188,instqueuewr_addr_reg_0_ );
   nor U16722 ( n16358,n16304,n11732 );
   nand U16723 ( n11732,n16372,state2_reg_0_ );
   nor U16724 ( n16372,n11708,n9391 );
   nand U16725 ( n16304,n16373,n16374 );
   nor U16726 ( n16374,n8866,n12994 );
   nor U16727 ( n12994,n10808,n15063 );
   not U16728 ( n8866,n15215 );
   nand U16729 ( n15215,n14979,n10808 );
   not U16730 ( n14979,n15063 );
   nand U16731 ( n15063,n9391,state2_reg_0_ );
   not U16732 ( n9391,n10818 );
   nor U16733 ( n16373,n16375,n16376 );
   nor U16734 ( n16376,n12992,n16333 );
   nand U16735 ( n16333,n11708,state2_reg_0_ );
   not U16736 ( n11708,n10778 );
   nand U16737 ( n10778,n16377,n16378 );
   nor U16738 ( n16378,n16379,n16380 );
   nand U16739 ( n16380,n16381,n16382 );
   nor U16740 ( n16382,n16383,n16384 );
   nor U16741 ( n16384,n16169,n15306 );
   not U16742 ( n15306,instqueue_reg_10__4_ );
   nor U16743 ( n16383,n16170,n15326 );
   not U16744 ( n15326,instqueue_reg_8__4_ );
   nor U16745 ( n16381,n16385,n16386 );
   nor U16746 ( n16386,n16173,n15318 );
   not U16747 ( n15318,instqueue_reg_15__4_ );
   nor U16748 ( n16385,n16174,n15317 );
   not U16749 ( n15317,instqueue_reg_14__4_ );
   nand U16750 ( n16379,n16387,n16388 );
   nor U16751 ( n16388,n16389,n16390 );
   nor U16752 ( n16390,n16179,n10781 );
   not U16753 ( n10781,instqueue_reg_0__4_ );
   nor U16754 ( n16389,n16220,n15295 );
   not U16755 ( n15295,instqueue_reg_3__4_ );
   nor U16756 ( n16387,n16391,n16392 );
   nor U16757 ( n16392,n16183,n15327 );
   not U16758 ( n15327,instqueue_reg_12__4_ );
   nor U16759 ( n16391,n16184,n15313 );
   not U16760 ( n15313,instqueue_reg_11__4_ );
   nor U16761 ( n16377,n16393,n16394 );
   nand U16762 ( n16394,n16395,n16396 );
   nor U16763 ( n16396,n16397,n16398 );
   nor U16764 ( n16398,n16191,n15301 );
   not U16765 ( n15301,instqueue_reg_6__4_ );
   nor U16766 ( n16397,n16192,n15296 );
   not U16767 ( n15296,instqueue_reg_5__4_ );
   nor U16768 ( n16395,n16399,n16400 );
   nor U16769 ( n16400,n16195,n15323 );
   not U16770 ( n15323,instqueue_reg_4__4_ );
   nor U16771 ( n16399,n16196,n15292 );
   not U16772 ( n15292,instqueue_reg_2__4_ );
   nand U16773 ( n16393,n16401,n16402 );
   nor U16774 ( n16402,n16403,n16404 );
   nor U16775 ( n16404,n16201,n15305 );
   not U16776 ( n15305,instqueue_reg_9__4_ );
   nor U16777 ( n16403,n16202,n15314 );
   not U16778 ( n15314,instqueue_reg_13__4_ );
   nor U16779 ( n16401,n16405,n16406 );
   nor U16780 ( n16406,n16205,n15291 );
   not U16781 ( n15291,instqueue_reg_1__4_ );
   nor U16782 ( n16405,n15605,n15302 );
   not U16783 ( n15302,instqueue_reg_7__4_ );
   nand U16784 ( n12992,n10808,n10818 );
   nor U16785 ( n16375,n16407,n8863 );
   not U16786 ( n8863,state2_reg_0_ );
   nor U16787 ( n16407,n12386,n8874 );
   not U16788 ( n8874,n12359 );
   nand U16789 ( n12359,n10906,n10818 );
   nand U16790 ( n10818,n16408,n16409 );
   nor U16791 ( n16409,n16410,n16411 );
   nand U16792 ( n16411,n16412,n16413 );
   nor U16793 ( n16413,n16414,n16415 );
   nor U16794 ( n16415,n16169,n15019 );
   not U16795 ( n15019,instqueue_reg_10__0_ );
   nor U16796 ( n16414,n16170,n15046 );
   not U16797 ( n15046,instqueue_reg_8__0_ );
   nor U16798 ( n16412,n16416,n16417 );
   nor U16799 ( n16417,n16173,n15035 );
   not U16800 ( n15035,instqueue_reg_15__0_ );
   nor U16801 ( n16416,n16174,n15033 );
   not U16802 ( n15033,instqueue_reg_14__0_ );
   nand U16803 ( n16410,n16418,n16419 );
   nor U16804 ( n16419,n16420,n16421 );
   nor U16805 ( n16421,n16179,n10825 );
   not U16806 ( n10825,instqueue_reg_0__0_ );
   nor U16807 ( n16420,n16180,n15003 );
   not U16808 ( n15003,instqueue_reg_3__0_ );
   nor U16809 ( n16418,n16422,n16423 );
   nor U16810 ( n16423,n16183,n15048 );
   not U16811 ( n15048,instqueue_reg_12__0_ );
   nor U16812 ( n16422,n16184,n15027 );
   not U16813 ( n15027,instqueue_reg_11__0_ );
   nor U16814 ( n16408,n16424,n16425 );
   nand U16815 ( n16425,n16426,n16427 );
   nor U16816 ( n16427,n16428,n16429 );
   nor U16817 ( n16429,n16191,n15011 );
   not U16818 ( n15011,instqueue_reg_6__0_ );
   nor U16819 ( n16428,n16192,n15005 );
   not U16820 ( n15005,instqueue_reg_5__0_ );
   nor U16821 ( n16426,n16430,n16431 );
   nor U16822 ( n16431,n16195,n15042 );
   not U16823 ( n15042,instqueue_reg_4__0_ );
   nor U16824 ( n16430,n16196,n14999 );
   not U16825 ( n14999,instqueue_reg_2__0_ );
   nand U16826 ( n16424,n16432,n16433 );
   nor U16827 ( n16433,n16434,n16435 );
   nor U16828 ( n16435,n16201,n15017 );
   not U16829 ( n15017,instqueue_reg_9__0_ );
   nor U16830 ( n16434,n16202,n15029 );
   not U16831 ( n15029,instqueue_reg_13__0_ );
   nor U16832 ( n16432,n16436,n16437 );
   nor U16833 ( n16437,n16205,n14997 );
   not U16834 ( n14997,instqueue_reg_1__0_ );
   nor U16835 ( n16436,n15605,n15013 );
   not U16836 ( n15013,instqueue_reg_7__0_ );
   not U16837 ( n10906,n10808 );
   nand U16838 ( n10808,n16438,n16439 );
   nor U16839 ( n16439,n16440,n16441 );
   nand U16840 ( n16441,n16442,n16443 );
   nor U16841 ( n16443,n16444,n16445 );
   nor U16842 ( n16445,n16169,n14925 );
   not U16843 ( n14925,instqueue_reg_10__1_ );
   nor U16844 ( n16444,n16170,n14929 );
   not U16845 ( n14929,instqueue_reg_8__1_ );
   nor U16846 ( n16442,n16446,n16447 );
   nor U16847 ( n16447,n16173,n14916 );
   not U16848 ( n14916,instqueue_reg_15__1_ );
   nor U16849 ( n16446,n16174,n14915 );
   not U16850 ( n14915,instqueue_reg_14__1_ );
   nand U16851 ( n16440,n16448,n16449 );
   nor U16852 ( n16449,n16450,n16451 );
   nor U16853 ( n16451,n16179,n10811 );
   not U16854 ( n10811,instqueue_reg_0__1_ );
   nor U16855 ( n16450,n16180,n14948 );
   not U16856 ( n14948,instqueue_reg_3__1_ );
   nand U16857 ( n16180,n16452,n10861 );
   nor U16858 ( n16448,n16453,n16454 );
   nor U16859 ( n16454,n16183,n14919 );
   not U16860 ( n14919,instqueue_reg_12__1_ );
   nor U16861 ( n16453,n16184,n14926 );
   not U16862 ( n14926,instqueue_reg_11__1_ );
   nor U16863 ( n16438,n16455,n16456 );
   nand U16864 ( n16456,n16457,n16458 );
   nor U16865 ( n16458,n16459,n16460 );
   nor U16866 ( n16460,n16191,n14937 );
   not U16867 ( n14937,instqueue_reg_6__1_ );
   nor U16868 ( n16459,n16192,n14942 );
   not U16869 ( n14942,instqueue_reg_5__1_ );
   nor U16870 ( n16457,n16461,n16462 );
   nor U16871 ( n16462,n16195,n14941 );
   not U16872 ( n14941,instqueue_reg_4__1_ );
   nor U16873 ( n16461,n16196,n14947 );
   not U16874 ( n14947,instqueue_reg_2__1_ );
   nand U16875 ( n16455,n16463,n16464 );
   nor U16876 ( n16464,n16465,n16466 );
   nor U16877 ( n16466,n16201,n14930 );
   not U16878 ( n14930,instqueue_reg_9__1_ );
   nor U16879 ( n16465,n16202,n14920 );
   not U16880 ( n14920,instqueue_reg_13__1_ );
   nor U16881 ( n16463,n16467,n16468 );
   nor U16882 ( n16468,n16205,n14951 );
   not U16883 ( n14951,instqueue_reg_1__1_ );
   nor U16884 ( n16467,n15605,n14938 );
   not U16885 ( n14938,instqueue_reg_7__1_ );
   nor U16886 ( n12386,n15230,n16469 );
   nor U16887 ( n16469,n10771,n16179 );
   nand U16888 ( n16179,n15832,n14172 );
   not U16889 ( n10771,instqueue_reg_0__5_ );
   nand U16890 ( n15230,n16470,n16471 );
   nor U16891 ( n16471,n16472,n16473 );
   nand U16892 ( n16473,n16474,n16475 );
   nor U16893 ( n16475,n16476,n16477 );
   nor U16894 ( n16477,n16174,n15364 );
   not U16895 ( n15364,instqueue_reg_14__5_ );
   nand U16896 ( n16174,n15887,instqueuerd_addr_reg_3_ );
   nor U16897 ( n15887,n15878,n10864 );
   nor U16898 ( n16476,n16169,n15353 );
   not U16899 ( n15353,instqueue_reg_10__5_ );
   nand U16900 ( n16169,n15623,n15906 );
   nor U16901 ( n16474,n16478,n16479 );
   nor U16902 ( n16479,n16202,n15361 );
   not U16903 ( n15361,instqueue_reg_13__5_ );
   nand U16904 ( n16202,n15886,instqueuerd_addr_reg_3_ );
   nor U16905 ( n15886,n15876,n10864 );
   nor U16906 ( n16478,n16173,n15365 );
   not U16907 ( n15365,instqueue_reg_15__5_ );
   nand U16908 ( n16173,n15607,instqueuerd_addr_reg_3_ );
   nor U16909 ( n15607,n10864,n15830 );
   nand U16910 ( n16472,n16480,n16481 );
   nor U16911 ( n16481,n16482,n16483 );
   nor U16912 ( n16483,n16184,n15360 );
   not U16913 ( n15360,instqueue_reg_11__5_ );
   nand U16914 ( n16184,instqueuerd_addr_reg_3_,n15609 );
   nor U16915 ( n16482,n16220,n15342 );
   not U16916 ( n15342,instqueue_reg_3__5_ );
   nand U16917 ( n16220,n15609,n14172 );
   nor U16918 ( n15609,n15830,instqueuerd_addr_reg_2_ );
   nor U16919 ( n16480,n16484,n16485 );
   nor U16920 ( n16485,n16170,n15373 );
   not U16921 ( n15373,instqueue_reg_8__5_ );
   nand U16922 ( n16170,instqueuerd_addr_reg_3_,n15832 );
   nor U16923 ( n15832,n10868,instqueuerd_addr_reg_2_ );
   nor U16924 ( n16484,n16183,n15374 );
   not U16925 ( n15374,instqueue_reg_12__5_ );
   nand U16926 ( n16183,n15881,instqueuerd_addr_reg_3_ );
   nor U16927 ( n15881,n10864,n10868 );
   nor U16928 ( n16470,n16486,n16487 );
   nand U16929 ( n16487,n16488,n16489 );
   or U16930 ( n16489,n15370,n16195 );
   nand U16931 ( n16195,n15652,n15619 );
   not U16932 ( n15619,n10868 );
   nand U16933 ( n10868,n8968,n9339 );
   not U16934 ( n15370,instqueue_reg_4__5_ );
   nor U16935 ( n16488,n16490,n16491 );
   nor U16936 ( n16491,n16196,n15339 );
   not U16937 ( n15339,instqueue_reg_2__5_ );
   nand U16938 ( n16196,n15623,n16452 );
   nor U16939 ( n16490,n16191,n15348 );
   not U16940 ( n15348,instqueue_reg_6__5_ );
   nand U16941 ( n16191,n15652,n15623 );
   not U16942 ( n15623,n15878 );
   nand U16943 ( n15878,instqueuerd_addr_reg_1_,n8968 );
   not U16944 ( n8968,instqueuerd_addr_reg_0_ );
   nand U16945 ( n16486,n16492,n16493 );
   nor U16946 ( n16493,n16494,n16495 );
   nor U16947 ( n16495,n15605,n15349 );
   not U16948 ( n15349,instqueue_reg_7__5_ );
   nand U16949 ( n15605,n15652,n10861 );
   not U16950 ( n10861,n15830 );
   nand U16951 ( n15830,instqueuerd_addr_reg_1_,instqueuerd_addr_reg_0_ );
   nor U16952 ( n16494,n16201,n15352 );
   not U16953 ( n15352,instqueue_reg_9__5_ );
   nand U16954 ( n16201,n15620,n15906 );
   nor U16955 ( n15906,n14172,instqueuerd_addr_reg_2_ );
   nor U16956 ( n16492,n16496,n16497 );
   nor U16957 ( n16497,n16192,n15343 );
   not U16958 ( n15343,instqueue_reg_5__5_ );
   nand U16959 ( n16192,n15652,n15620 );
   nor U16960 ( n15652,n10864,instqueuerd_addr_reg_3_ );
   nor U16961 ( n16496,n16205,n15338 );
   not U16962 ( n15338,instqueue_reg_1__5_ );
   nand U16963 ( n16205,n15620,n16452 );
   not U16964 ( n16452,n10862 );
   nand U16965 ( n10862,n10864,n14172 );
   not U16966 ( n14172,instqueuerd_addr_reg_3_ );
   not U16967 ( n10864,instqueuerd_addr_reg_2_ );
   not U16968 ( n15620,n15876 );
   nand U16969 ( n15876,instqueuerd_addr_reg_0_,n9339 );
   not U16970 ( n9339,instqueuerd_addr_reg_1_ );
   not U16971 ( n9287,n9015 );
   nand U16972 ( n9015,state2_reg_0_,n9275 );
   not U16973 ( n9275,n12996 );
   nand U16974 ( n12996,state2_reg_2_,n8948 );
   not U16975 ( n8948,state2_reg_1_ );
endmodule
