
module b21 ( si_31_, si_30_, si_29_, si_28_, si_27_, si_26_, si_25_, si_24_,         si_23_, si_22_, si_21_, si_20_, si_19_, si_18_, si_17_, si_16_, si_15_,         si_14_, si_13_, si_12_, si_11_, si_10_, si_9_, si_8_, si_7_, si_6_,         si_5_, si_4_, si_3_, si_2_, si_1_, si_0_, p1_ir_reg_0_, p1_ir_reg_1_,         p1_ir_reg_2_, p1_ir_reg_3_, p1_ir_reg_4_, p1_ir_reg_5_, p1_ir_reg_6_,         p1_ir_reg_7_, p1_ir_reg_8_, p1_ir_reg_9_, p1_ir_reg_10_, p1_ir_reg_11_,         p1_ir_reg_12_, p1_ir_reg_13_, p1_ir_reg_14_, p1_ir_reg_15_,         p1_ir_reg_16_, p1_ir_reg_17_, p1_ir_reg_18_, p1_ir_reg_19_,         p1_ir_reg_20_, p1_ir_reg_21_, p1_ir_reg_22_, p1_ir_reg_23_,         p1_ir_reg_24_, p1_ir_reg_25_, p1_ir_reg_26_, p1_ir_reg_27_,         p1_ir_reg_28_, p1_ir_reg_29_, p1_ir_reg_30_, p1_ir_reg_31_,         p1_d_reg_0_, p1_d_reg_1_, p1_d_reg_2_, p1_d_reg_3_, p1_d_reg_4_,         p1_d_reg_5_, p1_d_reg_6_, p1_d_reg_7_, p1_d_reg_8_, p1_d_reg_9_,         p1_d_reg_10_, p1_d_reg_11_, p1_d_reg_12_, p1_d_reg_13_, p1_d_reg_14_,         p1_d_reg_15_, p1_d_reg_16_, p1_d_reg_17_, p1_d_reg_18_, p1_d_reg_19_,         p1_d_reg_20_, p1_d_reg_21_, p1_d_reg_22_, p1_d_reg_23_, p1_d_reg_24_,         p1_d_reg_25_, p1_d_reg_26_, p1_d_reg_27_, p1_d_reg_28_, p1_d_reg_29_,         p1_d_reg_30_, p1_d_reg_31_, p1_reg0_reg_0_, p1_reg0_reg_1_,         p1_reg0_reg_2_, p1_reg0_reg_3_, p1_reg0_reg_4_, p1_reg0_reg_5_,         p1_reg0_reg_6_, p1_reg0_reg_7_, p1_reg0_reg_8_, p1_reg0_reg_9_,         p1_reg0_reg_10_, p1_reg0_reg_11_, p1_reg0_reg_12_, p1_reg0_reg_13_,         p1_reg0_reg_14_, p1_reg0_reg_15_, p1_reg0_reg_16_, p1_reg0_reg_17_,         p1_reg0_reg_18_, p1_reg0_reg_19_, p1_reg0_reg_20_, p1_reg0_reg_21_,         p1_reg0_reg_22_, p1_reg0_reg_23_, p1_reg0_reg_24_, p1_reg0_reg_25_,         p1_reg0_reg_26_, p1_reg0_reg_27_, p1_reg0_reg_28_, p1_reg0_reg_29_,         p1_reg0_reg_30_, p1_reg0_reg_31_, p1_reg1_reg_0_, p1_reg1_reg_1_,         p1_reg1_reg_2_, p1_reg1_reg_3_, p1_reg1_reg_4_, p1_reg1_reg_5_,         p1_reg1_reg_6_, p1_reg1_reg_7_, p1_reg1_reg_8_, p1_reg1_reg_9_,         p1_reg1_reg_10_, p1_reg1_reg_11_, p1_reg1_reg_12_, p1_reg1_reg_13_,         p1_reg1_reg_14_, p1_reg1_reg_15_, p1_reg1_reg_16_, p1_reg1_reg_17_,         p1_reg1_reg_18_, p1_reg1_reg_19_, p1_reg1_reg_20_, p1_reg1_reg_21_,         p1_reg1_reg_22_, p1_reg1_reg_23_, p1_reg1_reg_24_, p1_reg1_reg_25_,         p1_reg1_reg_26_, p1_reg1_reg_27_, p1_reg1_reg_28_, p1_reg1_reg_29_,         p1_reg1_reg_30_, p1_reg1_reg_31_, p1_reg2_reg_0_, p1_reg2_reg_1_,         p1_reg2_reg_2_, p1_reg2_reg_3_, p1_reg2_reg_4_, p1_reg2_reg_5_,         p1_reg2_reg_6_, p1_reg2_reg_7_, p1_reg2_reg_8_, p1_reg2_reg_9_,         p1_reg2_reg_10_, p1_reg2_reg_11_, p1_reg2_reg_12_, p1_reg2_reg_13_,         p1_reg2_reg_14_, p1_reg2_reg_15_, p1_reg2_reg_16_, p1_reg2_reg_17_,         p1_reg2_reg_18_, p1_reg2_reg_19_, p1_reg2_reg_20_, p1_reg2_reg_21_,         p1_reg2_reg_22_, p1_reg2_reg_23_, p1_reg2_reg_24_, p1_reg2_reg_25_,         p1_reg2_reg_26_, p1_reg2_reg_27_, p1_reg2_reg_28_, p1_reg2_reg_29_,         p1_reg2_reg_30_, p1_reg2_reg_31_, p1_addr_reg_19_, p1_addr_reg_18_,         p1_addr_reg_17_, p1_addr_reg_16_, p1_addr_reg_15_, p1_addr_reg_14_,         p1_addr_reg_13_, p1_addr_reg_12_, p1_addr_reg_11_, p1_addr_reg_10_,         p1_addr_reg_9_, p1_addr_reg_8_, p1_addr_reg_7_, p1_addr_reg_6_,         p1_addr_reg_5_, p1_addr_reg_4_, p1_addr_reg_3_, p1_addr_reg_2_,         p1_addr_reg_1_, p1_addr_reg_0_, p1_datao_reg_0_, p1_datao_reg_1_,         p1_datao_reg_2_, p1_datao_reg_3_, p1_datao_reg_4_, p1_datao_reg_5_,         p1_datao_reg_6_, p1_datao_reg_7_, p1_datao_reg_8_, p1_datao_reg_9_,         p1_datao_reg_10_, p1_datao_reg_11_, p1_datao_reg_12_, p1_datao_reg_13_,         p1_datao_reg_14_, p1_datao_reg_15_, p1_datao_reg_16_, p1_datao_reg_17_,         p1_datao_reg_18_, p1_datao_reg_19_, p1_datao_reg_20_, p1_datao_reg_21_,         p1_datao_reg_22_, p1_datao_reg_23_, p1_datao_reg_24_, p1_datao_reg_25_,         p1_datao_reg_26_, p1_datao_reg_27_, p1_datao_reg_28_, p1_datao_reg_29_,         p1_datao_reg_30_, p1_datao_reg_31_, p1_b_reg, p1_reg3_reg_15_,         p1_reg3_reg_26_, p1_reg3_reg_6_, p1_reg3_reg_18_, p1_reg3_reg_2_,         p1_reg3_reg_11_, p1_reg3_reg_22_, p1_reg3_reg_13_, p1_reg3_reg_20_,         p1_reg3_reg_0_, p1_reg3_reg_9_, p1_reg3_reg_4_, p1_reg3_reg_24_,         p1_reg3_reg_17_, p1_reg3_reg_5_, p1_reg3_reg_16_, p1_reg3_reg_25_,         p1_reg3_reg_12_, p1_reg3_reg_21_, p1_reg3_reg_1_, p1_reg3_reg_8_,         p1_reg3_reg_28_, p1_reg3_reg_19_, p1_reg3_reg_3_, p1_reg3_reg_10_,         p1_reg3_reg_23_, p1_reg3_reg_14_, p1_reg3_reg_27_, p1_reg3_reg_7_,         p1_state_reg, p1_rd_reg, p1_wr_reg, p2_ir_reg_0_, p2_ir_reg_1_,         p2_ir_reg_2_, p2_ir_reg_3_, p2_ir_reg_4_, p2_ir_reg_5_, p2_ir_reg_6_,         p2_ir_reg_7_, p2_ir_reg_8_, p2_ir_reg_9_, p2_ir_reg_10_, p2_ir_reg_11_,         p2_ir_reg_12_, p2_ir_reg_13_, p2_ir_reg_14_, p2_ir_reg_15_,         p2_ir_reg_16_, p2_ir_reg_17_, p2_ir_reg_18_, p2_ir_reg_19_,         p2_ir_reg_20_, p2_ir_reg_21_, p2_ir_reg_22_, p2_ir_reg_23_,         p2_ir_reg_24_, p2_ir_reg_25_, p2_ir_reg_26_, p2_ir_reg_27_,         p2_ir_reg_28_, p2_ir_reg_29_, p2_ir_reg_30_, p2_ir_reg_31_,         p2_d_reg_0_, p2_d_reg_1_, p2_d_reg_2_, p2_d_reg_3_, p2_d_reg_4_,         p2_d_reg_5_, p2_d_reg_6_, p2_d_reg_7_, p2_d_reg_8_, p2_d_reg_9_,         p2_d_reg_10_, p2_d_reg_11_, p2_d_reg_12_, p2_d_reg_13_, p2_d_reg_14_,         p2_d_reg_15_, p2_d_reg_16_, p2_d_reg_17_, p2_d_reg_18_, p2_d_reg_19_,         p2_d_reg_20_, p2_d_reg_21_, p2_d_reg_22_, p2_d_reg_23_, p2_d_reg_24_,         p2_d_reg_25_, p2_d_reg_26_, p2_d_reg_27_, p2_d_reg_28_, p2_d_reg_29_,         p2_d_reg_30_, p2_d_reg_31_, p2_reg0_reg_0_, p2_reg0_reg_1_,         p2_reg0_reg_2_, p2_reg0_reg_3_, p2_reg0_reg_4_, p2_reg0_reg_5_,         p2_reg0_reg_6_, p2_reg0_reg_7_, p2_reg0_reg_8_, p2_reg0_reg_9_,         p2_reg0_reg_10_, p2_reg0_reg_11_, p2_reg0_reg_12_, p2_reg0_reg_13_,         p2_reg0_reg_14_, p2_reg0_reg_15_, p2_reg0_reg_16_, p2_reg0_reg_17_,         p2_reg0_reg_18_, p2_reg0_reg_19_, p2_reg0_reg_20_, p2_reg0_reg_21_,         p2_reg0_reg_22_, p2_reg0_reg_23_, p2_reg0_reg_24_, p2_reg0_reg_25_,         p2_reg0_reg_26_, p2_reg0_reg_27_, p2_reg0_reg_28_, p2_reg0_reg_29_,         p2_reg0_reg_30_, p2_reg0_reg_31_, p2_reg1_reg_0_, p2_reg1_reg_1_,         p2_reg1_reg_2_, p2_reg1_reg_3_, p2_reg1_reg_4_, p2_reg1_reg_5_,         p2_reg1_reg_6_, p2_reg1_reg_7_, p2_reg1_reg_8_, p2_reg1_reg_9_,         p2_reg1_reg_10_, p2_reg1_reg_11_, p2_reg1_reg_12_, p2_reg1_reg_13_,         p2_reg1_reg_14_, p2_reg1_reg_15_, p2_reg1_reg_16_, p2_reg1_reg_17_,         p2_reg1_reg_18_, p2_reg1_reg_19_, p2_reg1_reg_20_, p2_reg1_reg_21_,         p2_reg1_reg_22_, p2_reg1_reg_23_, p2_reg1_reg_24_, p2_reg1_reg_25_,         p2_reg1_reg_26_, p2_reg1_reg_27_, p2_reg1_reg_28_, p2_reg1_reg_29_,         p2_reg1_reg_30_, p2_reg1_reg_31_, p2_reg2_reg_0_, p2_reg2_reg_1_,         p2_reg2_reg_2_, p2_reg2_reg_3_, p2_reg2_reg_4_, p2_reg2_reg_5_,         p2_reg2_reg_6_, p2_reg2_reg_7_, p2_reg2_reg_8_, p2_reg2_reg_9_,         p2_reg2_reg_10_, p2_reg2_reg_11_, p2_reg2_reg_12_, p2_reg2_reg_13_,         p2_reg2_reg_14_, p2_reg2_reg_15_, p2_reg2_reg_16_, p2_reg2_reg_17_,         p2_reg2_reg_18_, p2_reg2_reg_19_, p2_reg2_reg_20_, p2_reg2_reg_21_,         p2_reg2_reg_22_, p2_reg2_reg_23_, p2_reg2_reg_24_, p2_reg2_reg_25_,         p2_reg2_reg_26_, p2_reg2_reg_27_, p2_reg2_reg_28_, p2_reg2_reg_29_,         p2_reg2_reg_30_, p2_reg2_reg_31_, p2_addr_reg_19_, p2_addr_reg_18_,         p2_addr_reg_17_, p2_addr_reg_16_, p2_addr_reg_15_, p2_addr_reg_14_,         p2_addr_reg_13_, p2_addr_reg_12_, p2_addr_reg_11_, p2_addr_reg_10_,         p2_addr_reg_9_, p2_addr_reg_8_, p2_addr_reg_7_, p2_addr_reg_6_,         p2_addr_reg_5_, p2_addr_reg_4_, p2_addr_reg_3_, p2_addr_reg_2_,         p2_addr_reg_1_, p2_addr_reg_0_, p2_datao_reg_0_, p2_datao_reg_1_,         p2_datao_reg_2_, p2_datao_reg_3_, p2_datao_reg_4_, p2_datao_reg_5_,         p2_datao_reg_6_, p2_datao_reg_7_, p2_datao_reg_8_, p2_datao_reg_9_,         p2_datao_reg_10_, p2_datao_reg_11_, p2_datao_reg_12_, p2_datao_reg_13_,         p2_datao_reg_14_, p2_datao_reg_15_, p2_datao_reg_16_, p2_datao_reg_17_,         p2_datao_reg_18_, p2_datao_reg_19_, p2_datao_reg_20_, p2_datao_reg_21_,         p2_datao_reg_22_, p2_datao_reg_23_, p2_datao_reg_24_, p2_datao_reg_25_,         p2_datao_reg_26_, p2_datao_reg_27_, p2_datao_reg_28_, p2_datao_reg_29_,         p2_datao_reg_30_, p2_datao_reg_31_, p2_b_reg, p2_reg3_reg_15_,         p2_reg3_reg_26_, p2_reg3_reg_6_, p2_reg3_reg_18_, p2_reg3_reg_2_,         p2_reg3_reg_11_, p2_reg3_reg_22_, p2_reg3_reg_13_, p2_reg3_reg_20_,         p2_reg3_reg_0_, p2_reg3_reg_9_, p2_reg3_reg_4_, p2_reg3_reg_24_,         p2_reg3_reg_17_, p2_reg3_reg_5_, p2_reg3_reg_16_, p2_reg3_reg_25_,         p2_reg3_reg_12_, p2_reg3_reg_21_, p2_reg3_reg_1_, p2_reg3_reg_8_,         p2_reg3_reg_28_, p2_reg3_reg_19_, p2_reg3_reg_3_, p2_reg3_reg_10_,         p2_reg3_reg_23_, p2_reg3_reg_14_, p2_reg3_reg_27_, p2_reg3_reg_7_,         p2_state_reg, p2_rd_reg, p2_wr_reg, add_1071_u4, add_1071_u55,         add_1071_u56, add_1071_u57, add_1071_u58, add_1071_u59, add_1071_u60,         add_1071_u61, add_1071_u62, add_1071_u63, add_1071_u47, add_1071_u48,         add_1071_u49, add_1071_u50, add_1071_u51, add_1071_u52, add_1071_u53,         add_1071_u54, add_1071_u5, add_1071_u46, u126, u123, p1_u3353,         p1_u3352, p1_u3351, p1_u3350, p1_u3349, p1_u3348, p1_u3347, p1_u3346,         p1_u3345, p1_u3344, p1_u3343, p1_u3342, p1_u3341, p1_u3340, p1_u3339,         p1_u3338, p1_u3337, p1_u3336, p1_u3335, p1_u3334, p1_u3333, p1_u3332,         p1_u3331, p1_u3330, p1_u3329, p1_u3328, p1_u3327, p1_u3326, p1_u3325,         p1_u3324, p1_u3323, p1_u3322, p1_u3440, p1_u3441, p1_u3321, p1_u3320,         p1_u3319, p1_u3318, p1_u3317, p1_u3316, p1_u3315, p1_u3314, p1_u3313,         p1_u3312, p1_u3311, p1_u3310, p1_u3309, p1_u3308, p1_u3307, p1_u3306,         p1_u3305, p1_u3304, p1_u3303, p1_u3302, p1_u3301, p1_u3300, p1_u3299,         p1_u3298, p1_u3297, p1_u3296, p1_u3295, p1_u3294, p1_u3293, p1_u3292,         p1_u3454, p1_u3457, p1_u3460, p1_u3463, p1_u3466, p1_u3469, p1_u3472,         p1_u3475, p1_u3478, p1_u3481, p1_u3484, p1_u3487, p1_u3490, p1_u3493,         p1_u3496, p1_u3499, p1_u3502, p1_u3505, p1_u3508, p1_u3510, p1_u3511,         p1_u3512, p1_u3513, p1_u3514, p1_u3515, p1_u3516, p1_u3517, p1_u3518,         p1_u3519, p1_u3520, p1_u3521, p1_u3522, p1_u3523, p1_u3524, p1_u3525,         p1_u3526, p1_u3527, p1_u3528, p1_u3529, p1_u3530, p1_u3531, p1_u3532,         p1_u3533, p1_u3534, p1_u3535, p1_u3536, p1_u3537, p1_u3538, p1_u3539,         p1_u3540, p1_u3541, p1_u3542, p1_u3543, p1_u3544, p1_u3545, p1_u3546,         p1_u3547, p1_u3548, p1_u3549, p1_u3550, p1_u3551, p1_u3552, p1_u3553,         p1_u3554, p1_u3291, p1_u3290, p1_u3289, p1_u3288, p1_u3287, p1_u3286,         p1_u3285, p1_u3284, p1_u3283, p1_u3282, p1_u3281, p1_u3280, p1_u3279,         p1_u3278, p1_u3277, p1_u3276, p1_u3275, p1_u3274, p1_u3273, p1_u3272,         p1_u3271, p1_u3270, p1_u3269, p1_u3268, p1_u3267, p1_u3266, p1_u3265,         p1_u3264, p1_u3263, p1_u3355, p1_u3262, p1_u3261, p1_u3260, p1_u3259,         p1_u3258, p1_u3257, p1_u3256, p1_u3255, p1_u3254, p1_u3253, p1_u3252,         p1_u3251, p1_u3250, p1_u3249, p1_u3248, p1_u3247, p1_u3246, p1_u3245,         p1_u3244, p1_u3243, p1_u3242, p1_u3241, p1_u3555, p1_u3556, p1_u3557,         p1_u3558, p1_u3559, p1_u3560, p1_u3561, p1_u3562, p1_u3563, p1_u3564,         p1_u3565, p1_u3566, p1_u3567, p1_u3568, p1_u3569, p1_u3570, p1_u3571,         p1_u3572, p1_u3573, p1_u3574, p1_u3575, p1_u3576, p1_u3577, p1_u3578,         p1_u3579, p1_u3580, p1_u3581, p1_u3582, p1_u3583, p1_u3584, p1_u3585,         p1_u3586, p1_u3240, p1_u3239, p1_u3238, p1_u3237, p1_u3236, p1_u3235,         p1_u3234, p1_u3233, p1_u3232, p1_u3231, p1_u3230, p1_u3229, p1_u3228,         p1_u3227, p1_u3226, p1_u3225, p1_u3224, p1_u3223, p1_u3222, p1_u3221,         p1_u3220, p1_u3219, p1_u3218, p1_u3217, p1_u3216, p1_u3215, p1_u3214,         p1_u3213, p1_u3212, p1_u3211, p1_u3084, p1_u3083, p1_u4006, p2_u3358,         p2_u3357, p2_u3356, p2_u3355, p2_u3354, p2_u3353, p2_u3352, p2_u3351,         p2_u3350, p2_u3349, p2_u3348, p2_u3347, p2_u3346, p2_u3345, p2_u3344,         p2_u3343, p2_u3342, p2_u3341, p2_u3340, p2_u3339, p2_u3338, p2_u3337,         p2_u3336, p2_u3335, p2_u3334, p2_u3333, p2_u3332, p2_u3331, p2_u3330,         p2_u3329, p2_u3328, p2_u3327, p2_u3437, p2_u3438, p2_u3326, p2_u3325,         p2_u3324, p2_u3323, p2_u3322, p2_u3321, p2_u3320, p2_u3319, p2_u3318,         p2_u3317, p2_u3316, p2_u3315, p2_u3314, p2_u3313, p2_u3312, p2_u3311,         p2_u3310, p2_u3309, p2_u3308, p2_u3307, p2_u3306, p2_u3305, p2_u3304,         p2_u3303, p2_u3302, p2_u3301, p2_u3300, p2_u3299, p2_u3298, p2_u3297,         p2_u3451, p2_u3454, p2_u3457, p2_u3460, p2_u3463, p2_u3466, p2_u3469,         p2_u3472, p2_u3475, p2_u3478, p2_u3481, p2_u3484, p2_u3487, p2_u3490,         p2_u3493, p2_u3496, p2_u3499, p2_u3502, p2_u3505, p2_u3507, p2_u3508,         p2_u3509, p2_u3510, p2_u3511, p2_u3512, p2_u3513, p2_u3514, p2_u3515,         p2_u3516, p2_u3517, p2_u3518, p2_u3519, p2_u3520, p2_u3521, p2_u3522,         p2_u3523, p2_u3524, p2_u3525, p2_u3526, p2_u3527, p2_u3528, p2_u3529,         p2_u3530, p2_u3531, p2_u3532, p2_u3533, p2_u3534, p2_u3535, p2_u3536,         p2_u3537, p2_u3538, p2_u3539, p2_u3540, p2_u3541, p2_u3542, p2_u3543,         p2_u3544, p2_u3545, p2_u3546, p2_u3547, p2_u3548, p2_u3549, p2_u3550,         p2_u3551, p2_u3296, p2_u3295, p2_u3294, p2_u3293, p2_u3292, p2_u3291,         p2_u3290, p2_u3289, p2_u3288, p2_u3287, p2_u3286, p2_u3285, p2_u3284,         p2_u3283, p2_u3282, p2_u3281, p2_u3280, p2_u3279, p2_u3278, p2_u3277,         p2_u3276, p2_u3275, p2_u3274, p2_u3273, p2_u3272, p2_u3271, p2_u3270,         p2_u3269, p2_u3268, p2_u3267, p2_u3266, p2_u3265, p2_u3264, p2_u3263,         p2_u3262, p2_u3261, p2_u3260, p2_u3259, p2_u3258, p2_u3257, p2_u3256,         p2_u3255, p2_u3254, p2_u3253, p2_u3252, p2_u3251, p2_u3250, p2_u3249,         p2_u3248, p2_u3247, p2_u3246, p2_u3245, p2_u3552, p2_u3553, p2_u3554,         p2_u3555, p2_u3556, p2_u3557, p2_u3558, p2_u3559, p2_u3560, p2_u3561,         p2_u3562, p2_u3563, p2_u3564, p2_u3565, p2_u3566, p2_u3567, p2_u3568,         p2_u3569, p2_u3570, p2_u3571, p2_u3572, p2_u3573, p2_u3574, p2_u3575,         p2_u3576, p2_u3577, p2_u3578, p2_u3579, p2_u3580, p2_u3581, p2_u3582,         p2_u3583, p2_u3244, p2_u3243, p2_u3242, p2_u3241, p2_u3240, p2_u3239,         p2_u3238, p2_u3237, p2_u3236, p2_u3235, p2_u3234, p2_u3233, p2_u3232,         p2_u3231, p2_u3230, p2_u3229, p2_u3228, p2_u3227, p2_u3226, p2_u3225,         p2_u3224, p2_u3223, p2_u3222, p2_u3221, p2_u3220, p2_u3219, p2_u3218,         p2_u3217, p2_u3216, p2_u3215, p2_u3152, p2_u3151, p2_u3966 );
input si_31_, si_30_, si_29_, si_28_, si_27_, si_26_, si_25_, si_24_, si_23_,         si_22_, si_21_, si_20_, si_19_, si_18_, si_17_, si_16_, si_15_,         si_14_, si_13_, si_12_, si_11_, si_10_, si_9_, si_8_, si_7_, si_6_,         si_5_, si_4_, si_3_, si_2_, si_1_, si_0_, p1_ir_reg_0_, p1_ir_reg_1_,         p1_ir_reg_2_, p1_ir_reg_3_, p1_ir_reg_4_, p1_ir_reg_5_, p1_ir_reg_6_,         p1_ir_reg_7_, p1_ir_reg_8_, p1_ir_reg_9_, p1_ir_reg_10_,         p1_ir_reg_11_, p1_ir_reg_12_, p1_ir_reg_13_, p1_ir_reg_14_,         p1_ir_reg_15_, p1_ir_reg_16_, p1_ir_reg_17_, p1_ir_reg_18_,         p1_ir_reg_19_, p1_ir_reg_20_, p1_ir_reg_21_, p1_ir_reg_22_,         p1_ir_reg_23_, p1_ir_reg_24_, p1_ir_reg_25_, p1_ir_reg_26_,         p1_ir_reg_27_, p1_ir_reg_28_, p1_ir_reg_29_, p1_ir_reg_30_,         p1_ir_reg_31_, p1_d_reg_0_, p1_d_reg_1_, p1_d_reg_2_, p1_d_reg_3_,         p1_d_reg_4_, p1_d_reg_5_, p1_d_reg_6_, p1_d_reg_7_, p1_d_reg_8_,         p1_d_reg_9_, p1_d_reg_10_, p1_d_reg_11_, p1_d_reg_12_, p1_d_reg_13_,         p1_d_reg_14_, p1_d_reg_15_, p1_d_reg_16_, p1_d_reg_17_, p1_d_reg_18_,         p1_d_reg_19_, p1_d_reg_20_, p1_d_reg_21_, p1_d_reg_22_, p1_d_reg_23_,         p1_d_reg_24_, p1_d_reg_25_, p1_d_reg_26_, p1_d_reg_27_, p1_d_reg_28_,         p1_d_reg_29_, p1_d_reg_30_, p1_d_reg_31_, p1_reg0_reg_0_,         p1_reg0_reg_1_, p1_reg0_reg_2_, p1_reg0_reg_3_, p1_reg0_reg_4_,         p1_reg0_reg_5_, p1_reg0_reg_6_, p1_reg0_reg_7_, p1_reg0_reg_8_,         p1_reg0_reg_9_, p1_reg0_reg_10_, p1_reg0_reg_11_, p1_reg0_reg_12_,         p1_reg0_reg_13_, p1_reg0_reg_14_, p1_reg0_reg_15_, p1_reg0_reg_16_,         p1_reg0_reg_17_, p1_reg0_reg_18_, p1_reg0_reg_19_, p1_reg0_reg_20_,         p1_reg0_reg_21_, p1_reg0_reg_22_, p1_reg0_reg_23_, p1_reg0_reg_24_,         p1_reg0_reg_25_, p1_reg0_reg_26_, p1_reg0_reg_27_, p1_reg0_reg_28_,         p1_reg0_reg_29_, p1_reg0_reg_30_, p1_reg0_reg_31_, p1_reg1_reg_0_,         p1_reg1_reg_1_, p1_reg1_reg_2_, p1_reg1_reg_3_, p1_reg1_reg_4_,         p1_reg1_reg_5_, p1_reg1_reg_6_, p1_reg1_reg_7_, p1_reg1_reg_8_,         p1_reg1_reg_9_, p1_reg1_reg_10_, p1_reg1_reg_11_, p1_reg1_reg_12_,         p1_reg1_reg_13_, p1_reg1_reg_14_, p1_reg1_reg_15_, p1_reg1_reg_16_,         p1_reg1_reg_17_, p1_reg1_reg_18_, p1_reg1_reg_19_, p1_reg1_reg_20_,         p1_reg1_reg_21_, p1_reg1_reg_22_, p1_reg1_reg_23_, p1_reg1_reg_24_,         p1_reg1_reg_25_, p1_reg1_reg_26_, p1_reg1_reg_27_, p1_reg1_reg_28_,         p1_reg1_reg_29_, p1_reg1_reg_30_, p1_reg1_reg_31_, p1_reg2_reg_0_,         p1_reg2_reg_1_, p1_reg2_reg_2_, p1_reg2_reg_3_, p1_reg2_reg_4_,         p1_reg2_reg_5_, p1_reg2_reg_6_, p1_reg2_reg_7_, p1_reg2_reg_8_,         p1_reg2_reg_9_, p1_reg2_reg_10_, p1_reg2_reg_11_, p1_reg2_reg_12_,         p1_reg2_reg_13_, p1_reg2_reg_14_, p1_reg2_reg_15_, p1_reg2_reg_16_,         p1_reg2_reg_17_, p1_reg2_reg_18_, p1_reg2_reg_19_, p1_reg2_reg_20_,         p1_reg2_reg_21_, p1_reg2_reg_22_, p1_reg2_reg_23_, p1_reg2_reg_24_,         p1_reg2_reg_25_, p1_reg2_reg_26_, p1_reg2_reg_27_, p1_reg2_reg_28_,         p1_reg2_reg_29_, p1_reg2_reg_30_, p1_reg2_reg_31_, p1_addr_reg_19_,         p1_addr_reg_18_, p1_addr_reg_17_, p1_addr_reg_16_, p1_addr_reg_15_,         p1_addr_reg_14_, p1_addr_reg_13_, p1_addr_reg_12_, p1_addr_reg_11_,         p1_addr_reg_10_, p1_addr_reg_9_, p1_addr_reg_8_, p1_addr_reg_7_,         p1_addr_reg_6_, p1_addr_reg_5_, p1_addr_reg_4_, p1_addr_reg_3_,         p1_addr_reg_2_, p1_addr_reg_1_, p1_addr_reg_0_, p1_datao_reg_0_,         p1_datao_reg_1_, p1_datao_reg_2_, p1_datao_reg_3_, p1_datao_reg_4_,         p1_datao_reg_5_, p1_datao_reg_6_, p1_datao_reg_7_, p1_datao_reg_8_,         p1_datao_reg_9_, p1_datao_reg_10_, p1_datao_reg_11_, p1_datao_reg_12_,         p1_datao_reg_13_, p1_datao_reg_14_, p1_datao_reg_15_,         p1_datao_reg_16_, p1_datao_reg_17_, p1_datao_reg_18_,         p1_datao_reg_19_, p1_datao_reg_20_, p1_datao_reg_21_,         p1_datao_reg_22_, p1_datao_reg_23_, p1_datao_reg_24_,         p1_datao_reg_25_, p1_datao_reg_26_, p1_datao_reg_27_,         p1_datao_reg_28_, p1_datao_reg_29_, p1_datao_reg_30_,         p1_datao_reg_31_, p1_b_reg, p1_reg3_reg_15_, p1_reg3_reg_26_,         p1_reg3_reg_6_, p1_reg3_reg_18_, p1_reg3_reg_2_, p1_reg3_reg_11_,         p1_reg3_reg_22_, p1_reg3_reg_13_, p1_reg3_reg_20_, p1_reg3_reg_0_,         p1_reg3_reg_9_, p1_reg3_reg_4_, p1_reg3_reg_24_, p1_reg3_reg_17_,         p1_reg3_reg_5_, p1_reg3_reg_16_, p1_reg3_reg_25_, p1_reg3_reg_12_,         p1_reg3_reg_21_, p1_reg3_reg_1_, p1_reg3_reg_8_, p1_reg3_reg_28_,         p1_reg3_reg_19_, p1_reg3_reg_3_, p1_reg3_reg_10_, p1_reg3_reg_23_,         p1_reg3_reg_14_, p1_reg3_reg_27_, p1_reg3_reg_7_, p1_state_reg,         p1_rd_reg, p1_wr_reg, p2_ir_reg_0_, p2_ir_reg_1_, p2_ir_reg_2_,         p2_ir_reg_3_, p2_ir_reg_4_, p2_ir_reg_5_, p2_ir_reg_6_, p2_ir_reg_7_,         p2_ir_reg_8_, p2_ir_reg_9_, p2_ir_reg_10_, p2_ir_reg_11_,         p2_ir_reg_12_, p2_ir_reg_13_, p2_ir_reg_14_, p2_ir_reg_15_,         p2_ir_reg_16_, p2_ir_reg_17_, p2_ir_reg_18_, p2_ir_reg_19_,         p2_ir_reg_20_, p2_ir_reg_21_, p2_ir_reg_22_, p2_ir_reg_23_,         p2_ir_reg_24_, p2_ir_reg_25_, p2_ir_reg_26_, p2_ir_reg_27_,         p2_ir_reg_28_, p2_ir_reg_29_, p2_ir_reg_30_, p2_ir_reg_31_,         p2_d_reg_0_, p2_d_reg_1_, p2_d_reg_2_, p2_d_reg_3_, p2_d_reg_4_,         p2_d_reg_5_, p2_d_reg_6_, p2_d_reg_7_, p2_d_reg_8_, p2_d_reg_9_,         p2_d_reg_10_, p2_d_reg_11_, p2_d_reg_12_, p2_d_reg_13_, p2_d_reg_14_,         p2_d_reg_15_, p2_d_reg_16_, p2_d_reg_17_, p2_d_reg_18_, p2_d_reg_19_,         p2_d_reg_20_, p2_d_reg_21_, p2_d_reg_22_, p2_d_reg_23_, p2_d_reg_24_,         p2_d_reg_25_, p2_d_reg_26_, p2_d_reg_27_, p2_d_reg_28_, p2_d_reg_29_,         p2_d_reg_30_, p2_d_reg_31_, p2_reg0_reg_0_, p2_reg0_reg_1_,         p2_reg0_reg_2_, p2_reg0_reg_3_, p2_reg0_reg_4_, p2_reg0_reg_5_,         p2_reg0_reg_6_, p2_reg0_reg_7_, p2_reg0_reg_8_, p2_reg0_reg_9_,         p2_reg0_reg_10_, p2_reg0_reg_11_, p2_reg0_reg_12_, p2_reg0_reg_13_,         p2_reg0_reg_14_, p2_reg0_reg_15_, p2_reg0_reg_16_, p2_reg0_reg_17_,         p2_reg0_reg_18_, p2_reg0_reg_19_, p2_reg0_reg_20_, p2_reg0_reg_21_,         p2_reg0_reg_22_, p2_reg0_reg_23_, p2_reg0_reg_24_, p2_reg0_reg_25_,         p2_reg0_reg_26_, p2_reg0_reg_27_, p2_reg0_reg_28_, p2_reg0_reg_29_,         p2_reg0_reg_30_, p2_reg0_reg_31_, p2_reg1_reg_0_, p2_reg1_reg_1_,         p2_reg1_reg_2_, p2_reg1_reg_3_, p2_reg1_reg_4_, p2_reg1_reg_5_,         p2_reg1_reg_6_, p2_reg1_reg_7_, p2_reg1_reg_8_, p2_reg1_reg_9_,         p2_reg1_reg_10_, p2_reg1_reg_11_, p2_reg1_reg_12_, p2_reg1_reg_13_,         p2_reg1_reg_14_, p2_reg1_reg_15_, p2_reg1_reg_16_, p2_reg1_reg_17_,         p2_reg1_reg_18_, p2_reg1_reg_19_, p2_reg1_reg_20_, p2_reg1_reg_21_,         p2_reg1_reg_22_, p2_reg1_reg_23_, p2_reg1_reg_24_, p2_reg1_reg_25_,         p2_reg1_reg_26_, p2_reg1_reg_27_, p2_reg1_reg_28_, p2_reg1_reg_29_,         p2_reg1_reg_30_, p2_reg1_reg_31_, p2_reg2_reg_0_, p2_reg2_reg_1_,         p2_reg2_reg_2_, p2_reg2_reg_3_, p2_reg2_reg_4_, p2_reg2_reg_5_,         p2_reg2_reg_6_, p2_reg2_reg_7_, p2_reg2_reg_8_, p2_reg2_reg_9_,         p2_reg2_reg_10_, p2_reg2_reg_11_, p2_reg2_reg_12_, p2_reg2_reg_13_,         p2_reg2_reg_14_, p2_reg2_reg_15_, p2_reg2_reg_16_, p2_reg2_reg_17_,         p2_reg2_reg_18_, p2_reg2_reg_19_, p2_reg2_reg_20_, p2_reg2_reg_21_,         p2_reg2_reg_22_, p2_reg2_reg_23_, p2_reg2_reg_24_, p2_reg2_reg_25_,         p2_reg2_reg_26_, p2_reg2_reg_27_, p2_reg2_reg_28_, p2_reg2_reg_29_,         p2_reg2_reg_30_, p2_reg2_reg_31_, p2_addr_reg_19_, p2_addr_reg_18_,         p2_addr_reg_17_, p2_addr_reg_16_, p2_addr_reg_15_, p2_addr_reg_14_,         p2_addr_reg_13_, p2_addr_reg_12_, p2_addr_reg_11_, p2_addr_reg_10_,         p2_addr_reg_9_, p2_addr_reg_8_, p2_addr_reg_7_, p2_addr_reg_6_,         p2_addr_reg_5_, p2_addr_reg_4_, p2_addr_reg_3_, p2_addr_reg_2_,         p2_addr_reg_1_, p2_addr_reg_0_, p2_datao_reg_0_, p2_datao_reg_1_,         p2_datao_reg_2_, p2_datao_reg_3_, p2_datao_reg_4_, p2_datao_reg_5_,         p2_datao_reg_6_, p2_datao_reg_7_, p2_datao_reg_8_, p2_datao_reg_9_,         p2_datao_reg_10_, p2_datao_reg_11_, p2_datao_reg_12_,         p2_datao_reg_13_, p2_datao_reg_14_, p2_datao_reg_15_,         p2_datao_reg_16_, p2_datao_reg_17_, p2_datao_reg_18_,         p2_datao_reg_19_, p2_datao_reg_20_, p2_datao_reg_21_,         p2_datao_reg_22_, p2_datao_reg_23_, p2_datao_reg_24_,         p2_datao_reg_25_, p2_datao_reg_26_, p2_datao_reg_27_,         p2_datao_reg_28_, p2_datao_reg_29_, p2_datao_reg_30_,         p2_datao_reg_31_, p2_b_reg, p2_reg3_reg_15_, p2_reg3_reg_26_,         p2_reg3_reg_6_, p2_reg3_reg_18_, p2_reg3_reg_2_, p2_reg3_reg_11_,         p2_reg3_reg_22_, p2_reg3_reg_13_, p2_reg3_reg_20_, p2_reg3_reg_0_,         p2_reg3_reg_9_, p2_reg3_reg_4_, p2_reg3_reg_24_, p2_reg3_reg_17_,         p2_reg3_reg_5_, p2_reg3_reg_16_, p2_reg3_reg_25_, p2_reg3_reg_12_,         p2_reg3_reg_21_, p2_reg3_reg_1_, p2_reg3_reg_8_, p2_reg3_reg_28_,         p2_reg3_reg_19_, p2_reg3_reg_3_, p2_reg3_reg_10_, p2_reg3_reg_23_,         p2_reg3_reg_14_, p2_reg3_reg_27_, p2_reg3_reg_7_, p2_state_reg,         p2_rd_reg, p2_wr_reg;
output add_1071_u4, add_1071_u55, add_1071_u56, add_1071_u57, add_1071_u58,         add_1071_u59, add_1071_u60, add_1071_u61, add_1071_u62, add_1071_u63,         add_1071_u47, add_1071_u48, add_1071_u49, add_1071_u50, add_1071_u51,         add_1071_u52, add_1071_u53, add_1071_u54, add_1071_u5, add_1071_u46,         u126, u123, p1_u3353, p1_u3352, p1_u3351, p1_u3350, p1_u3349,         p1_u3348, p1_u3347, p1_u3346, p1_u3345, p1_u3344, p1_u3343, p1_u3342,         p1_u3341, p1_u3340, p1_u3339, p1_u3338, p1_u3337, p1_u3336, p1_u3335,         p1_u3334, p1_u3333, p1_u3332, p1_u3331, p1_u3330, p1_u3329, p1_u3328,         p1_u3327, p1_u3326, p1_u3325, p1_u3324, p1_u3323, p1_u3322, p1_u3440,         p1_u3441, p1_u3321, p1_u3320, p1_u3319, p1_u3318, p1_u3317, p1_u3316,         p1_u3315, p1_u3314, p1_u3313, p1_u3312, p1_u3311, p1_u3310, p1_u3309,         p1_u3308, p1_u3307, p1_u3306, p1_u3305, p1_u3304, p1_u3303, p1_u3302,         p1_u3301, p1_u3300, p1_u3299, p1_u3298, p1_u3297, p1_u3296, p1_u3295,         p1_u3294, p1_u3293, p1_u3292, p1_u3454, p1_u3457, p1_u3460, p1_u3463,         p1_u3466, p1_u3469, p1_u3472, p1_u3475, p1_u3478, p1_u3481, p1_u3484,         p1_u3487, p1_u3490, p1_u3493, p1_u3496, p1_u3499, p1_u3502, p1_u3505,         p1_u3508, p1_u3510, p1_u3511, p1_u3512, p1_u3513, p1_u3514, p1_u3515,         p1_u3516, p1_u3517, p1_u3518, p1_u3519, p1_u3520, p1_u3521, p1_u3522,         p1_u3523, p1_u3524, p1_u3525, p1_u3526, p1_u3527, p1_u3528, p1_u3529,         p1_u3530, p1_u3531, p1_u3532, p1_u3533, p1_u3534, p1_u3535, p1_u3536,         p1_u3537, p1_u3538, p1_u3539, p1_u3540, p1_u3541, p1_u3542, p1_u3543,         p1_u3544, p1_u3545, p1_u3546, p1_u3547, p1_u3548, p1_u3549, p1_u3550,         p1_u3551, p1_u3552, p1_u3553, p1_u3554, p1_u3291, p1_u3290, p1_u3289,         p1_u3288, p1_u3287, p1_u3286, p1_u3285, p1_u3284, p1_u3283, p1_u3282,         p1_u3281, p1_u3280, p1_u3279, p1_u3278, p1_u3277, p1_u3276, p1_u3275,         p1_u3274, p1_u3273, p1_u3272, p1_u3271, p1_u3270, p1_u3269, p1_u3268,         p1_u3267, p1_u3266, p1_u3265, p1_u3264, p1_u3263, p1_u3355, p1_u3262,         p1_u3261, p1_u3260, p1_u3259, p1_u3258, p1_u3257, p1_u3256, p1_u3255,         p1_u3254, p1_u3253, p1_u3252, p1_u3251, p1_u3250, p1_u3249, p1_u3248,         p1_u3247, p1_u3246, p1_u3245, p1_u3244, p1_u3243, p1_u3242, p1_u3241,         p1_u3555, p1_u3556, p1_u3557, p1_u3558, p1_u3559, p1_u3560, p1_u3561,         p1_u3562, p1_u3563, p1_u3564, p1_u3565, p1_u3566, p1_u3567, p1_u3568,         p1_u3569, p1_u3570, p1_u3571, p1_u3572, p1_u3573, p1_u3574, p1_u3575,         p1_u3576, p1_u3577, p1_u3578, p1_u3579, p1_u3580, p1_u3581, p1_u3582,         p1_u3583, p1_u3584, p1_u3585, p1_u3586, p1_u3240, p1_u3239, p1_u3238,         p1_u3237, p1_u3236, p1_u3235, p1_u3234, p1_u3233, p1_u3232, p1_u3231,         p1_u3230, p1_u3229, p1_u3228, p1_u3227, p1_u3226, p1_u3225, p1_u3224,         p1_u3223, p1_u3222, p1_u3221, p1_u3220, p1_u3219, p1_u3218, p1_u3217,         p1_u3216, p1_u3215, p1_u3214, p1_u3213, p1_u3212, p1_u3211, p1_u3084,         p1_u3083, p1_u4006, p2_u3358, p2_u3357, p2_u3356, p2_u3355, p2_u3354,         p2_u3353, p2_u3352, p2_u3351, p2_u3350, p2_u3349, p2_u3348, p2_u3347,         p2_u3346, p2_u3345, p2_u3344, p2_u3343, p2_u3342, p2_u3341, p2_u3340,         p2_u3339, p2_u3338, p2_u3337, p2_u3336, p2_u3335, p2_u3334, p2_u3333,         p2_u3332, p2_u3331, p2_u3330, p2_u3329, p2_u3328, p2_u3327, p2_u3437,         p2_u3438, p2_u3326, p2_u3325, p2_u3324, p2_u3323, p2_u3322, p2_u3321,         p2_u3320, p2_u3319, p2_u3318, p2_u3317, p2_u3316, p2_u3315, p2_u3314,         p2_u3313, p2_u3312, p2_u3311, p2_u3310, p2_u3309, p2_u3308, p2_u3307,         p2_u3306, p2_u3305, p2_u3304, p2_u3303, p2_u3302, p2_u3301, p2_u3300,         p2_u3299, p2_u3298, p2_u3297, p2_u3451, p2_u3454, p2_u3457, p2_u3460,         p2_u3463, p2_u3466, p2_u3469, p2_u3472, p2_u3475, p2_u3478, p2_u3481,         p2_u3484, p2_u3487, p2_u3490, p2_u3493, p2_u3496, p2_u3499, p2_u3502,         p2_u3505, p2_u3507, p2_u3508, p2_u3509, p2_u3510, p2_u3511, p2_u3512,         p2_u3513, p2_u3514, p2_u3515, p2_u3516, p2_u3517, p2_u3518, p2_u3519,         p2_u3520, p2_u3521, p2_u3522, p2_u3523, p2_u3524, p2_u3525, p2_u3526,         p2_u3527, p2_u3528, p2_u3529, p2_u3530, p2_u3531, p2_u3532, p2_u3533,         p2_u3534, p2_u3535, p2_u3536, p2_u3537, p2_u3538, p2_u3539, p2_u3540,         p2_u3541, p2_u3542, p2_u3543, p2_u3544, p2_u3545, p2_u3546, p2_u3547,         p2_u3548, p2_u3549, p2_u3550, p2_u3551, p2_u3296, p2_u3295, p2_u3294,         p2_u3293, p2_u3292, p2_u3291, p2_u3290, p2_u3289, p2_u3288, p2_u3287,         p2_u3286, p2_u3285, p2_u3284, p2_u3283, p2_u3282, p2_u3281, p2_u3280,         p2_u3279, p2_u3278, p2_u3277, p2_u3276, p2_u3275, p2_u3274, p2_u3273,         p2_u3272, p2_u3271, p2_u3270, p2_u3269, p2_u3268, p2_u3267, p2_u3266,         p2_u3265, p2_u3264, p2_u3263, p2_u3262, p2_u3261, p2_u3260, p2_u3259,         p2_u3258, p2_u3257, p2_u3256, p2_u3255, p2_u3254, p2_u3253, p2_u3252,         p2_u3251, p2_u3250, p2_u3249, p2_u3248, p2_u3247, p2_u3246, p2_u3245,         p2_u3552, p2_u3553, p2_u3554, p2_u3555, p2_u3556, p2_u3557, p2_u3558,         p2_u3559, p2_u3560, p2_u3561, p2_u3562, p2_u3563, p2_u3564, p2_u3565,         p2_u3566, p2_u3567, p2_u3568, p2_u3569, p2_u3570, p2_u3571, p2_u3572,         p2_u3573, p2_u3574, p2_u3575, p2_u3576, p2_u3577, p2_u3578, p2_u3579,         p2_u3580, p2_u3581, p2_u3582, p2_u3583, p2_u3244, p2_u3243, p2_u3242,         p2_u3241, p2_u3240, p2_u3239, p2_u3238, p2_u3237, p2_u3236, p2_u3235,         p2_u3234, p2_u3233, p2_u3232, p2_u3231, p2_u3230, p2_u3229, p2_u3228,         p2_u3227, p2_u3226, p2_u3225, p2_u3224, p2_u3223, p2_u3222, p2_u3221,         p2_u3220, p2_u3219, p2_u3218, p2_u3217, p2_u3216, p2_u3215, p2_u3152,         p2_u3151, p2_u3966;
wire   n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,         n19378, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,         n10009, n10010, n10011, n10012, n10032, n10034, n10037, n10040,         n10043, n10046, n10049, n10052, n10055, n10058, n10061, n10068,         n10069, n10071, n10072, n10076, n10077, n10079, n10080, n10084,         n10085, n10087, n10089, n10090, n10092, n10093, n10097, n10098,         n10100, n10101, n10103, n10104, n10106, n10107, n10147, n10150,         n10155, n10160, n10163, n10166, n10169, n10172, n10175, n10178,         n10189, n10192, n10197, n10200, n10205, n10208, n10211, n10216,         n10219, n10222, n10492, n10493, n10565, n10566, n10567, n10568,         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,         n18913;

   nand U9546 ( n16678,n16693,n16694,n16461 );
   nand U9547 ( n16604,n16619,n16620,n16461 );
   nand U9548 ( n16500,n16521,n16522,n16461 );
   nand U9549 ( n16435,n16459,n16460,n16461 );
   nand U9550 ( n16969,n16970,p1_state_reg,n16963 );
   or U9551 ( n9952,n12048,n12049,n12050,n12051 );
   or U9552 ( n9953,n12081,n12082,n12083,n12084 );
   or U9553 ( n9954,n12157,n12158,n12159,n12160 );
   or U9554 ( n9955,n12213,n12214,n12215,n12216 );
   or U9555 ( n9956,n12237,n12238,n12239,n12240 );
   or U9556 ( n9957,n12277,n12278,n12279,n12280 );
   or U9557 ( n9958,n11707,n11708,n11709,n11710 );
   or U9558 ( n9959,n11748,n11749,n11750,n11751 );
   or U9559 ( n9960,n11816,n11817,n11818,n11819 );
   or U9560 ( n9961,n11850,n11851,n11852,n11853 );
   or U9561 ( n9962,n11997,n11998,n11999,n12000 );
   or U9562 ( n9963,n12023,n12024,n12025,n12026 );
   or U9563 ( n9964,n9958,n9977 );
   or U9564 ( n9965,n9959,n9978 );
   or U9565 ( n9966,n9960,n9979 );
   or U9566 ( n9967,n9961,n9980 );
   or U9567 ( n9968,n9962,n9981 );
   or U9568 ( n9969,n9963,n9982 );
   or U9569 ( n9970,n9952,n9983 );
   or U9570 ( n9971,n9953,n9984 );
   or U9571 ( n9972,n9954,n9985 );
   or U9572 ( n9973,n9955,n9986 );
   or U9573 ( n9974,n9956,n9987 );
   or U9574 ( n9975,n9957,n9988 );
   nor U9575 ( n9976,n11460,n10908 );
   and U9576 ( n9977,n11461,n10630 );
   and U9577 ( n9978,n11461,n10627 );
   and U9578 ( n9979,n11461,n10621 );
   and U9579 ( n9980,n11461,n10618 );
   and U9580 ( n9981,n11461,n10606 );
   and U9581 ( n9982,n11461,n10603 );
   and U9582 ( n9983,n11461,n10600 );
   and U9583 ( n9984,n11461,n10597 );
   and U9584 ( n9985,n11461,n10591 );
   and U9585 ( n9986,n11461,n10585 );
   and U9586 ( n9987,n11461,n10582 );
   and U9587 ( n9988,n11461,n10579 );
   and U9588 ( n9989,n11479,n10974 );
   nor U9589 ( n9990,n11460,n11008 );
   nor U9590 ( n9991,n11460,n10996 );
   nor U9591 ( n9992,n11460,n10964 );
   nor U9592 ( n9993,n11460,n10898 );
   nor U9593 ( n9994,n11460,n10886 );
   nor U9594 ( n9995,n11460,n10864 );
   nor U9595 ( n9996,n11460,n10830 );
   nor U9596 ( n9997,n11460,n10818 );
   nor U9597 ( n9998,n11460,n10920 );
   nor U9598 ( n9999,n11460,n10839 );
   nor U9599 ( n10000,n11456,n10909 );
   or U9600 ( n10001,n9989,n10077 );
   or U9601 ( n10002,n10085,n9998 );
   or U9602 ( n10003,n9976,n10000 );
   or U9603 ( n10004,n10101,n9999 );
   or U9604 ( n10005,n9990,n10069 );
   or U9605 ( n10006,n9991,n10072 );
   or U9606 ( n10007,n9992,n10080 );
   or U9607 ( n10008,n9993,n10090 );
   or U9608 ( n10009,n9994,n10093 );
   or U9609 ( n10010,n9995,n10098 );
   or U9610 ( n10011,n9996,n10104 );
   or U9611 ( n10012,n9997,n10107 );
   nand U9612 ( n12563,n13060,n12365 );
   not U9613 ( n13589,n13574 );
   not U9614 ( n17500,n17575 );
   not U9615 ( n13572,n13591 );
   not U9616 ( n17515,n17507 );
   not U9617 ( n17497,n17576 );
   not U9618 ( n12572,n12538 );
   buf U9619 ( p2_u3319,n19199 );
   nor U9620 ( n19199,n11146,n11424 );
   buf U9621 ( p2_u3315,n19200 );
   nor U9622 ( n19200,n11146,n11425 );
   buf U9623 ( p2_u3320,n19198 );
   nor U9624 ( n19198,n11146,n11423 );
   buf U9625 ( p2_u3314,n19201 );
   nor U9626 ( n19201,n11146,n11426 );
   buf U9627 ( p2_u3321,n19197 );
   nor U9628 ( n19197,n11146,n11422 );
   buf U9629 ( p2_u3313,n19202 );
   nor U9630 ( n19202,n11146,n11427 );
   buf U9631 ( p2_u3322,n19196 );
   nor U9632 ( n19196,n11146,n11421 );
   buf U9633 ( p2_u3312,n19203 );
   nor U9634 ( n19203,n11146,n11428 );
   buf U9635 ( p2_u3323,n19195 );
   nor U9636 ( n19195,n11146,n11420 );
   buf U9637 ( p2_u3303,n19204 );
   nor U9638 ( n19204,n11146,n11429 );
   buf U9639 ( p2_u3298,n19209 );
   nor U9640 ( n19209,n11146,n11434 );
   buf U9641 ( p2_u3302,n19205 );
   nor U9642 ( n19205,n11146,n11430 );
   buf U9643 ( p2_u3297,n19210 );
   nor U9644 ( n19210,n11146,n11435 );
   buf U9645 ( p2_u3301,n19206 );
   nor U9646 ( n19206,n11146,n11431 );
   buf U9647 ( p2_u3324,n19194 );
   nor U9648 ( n19194,n11146,n11419 );
   buf U9649 ( p2_u3300,n19207 );
   nor U9650 ( n19207,n11146,n11432 );
   buf U9651 ( p2_u3326,n19192 );
   nor U9652 ( n19192,n11146,n11417 );
   buf U9653 ( p2_u3299,n19208 );
   nor U9654 ( n19208,n11146,n11433 );
   buf U9655 ( p2_u3325,n19193 );
   nor U9656 ( n19193,n11146,n11418 );
   nand U9657 ( n10032,n11145,p2_d_reg_10_ );
   not U9658 ( p2_u3318,n10032 );
   nand U9659 ( n10034,n11145,p2_d_reg_11_ );
   not U9660 ( p2_u3317,n10034 );
   buf U9661 ( p2_u3438,n19191 );
   nand U9662 ( n19191,n11143,n11144 );
   nand U9663 ( n10037,n11145,p2_d_reg_12_ );
   not U9664 ( p2_u3316,n10037 );
   buf U9665 ( p2_u3437,n19190 );
   nand U9666 ( n19190,n11148,n11149 );
   nand U9667 ( n10040,n11145,p2_d_reg_17_ );
   not U9668 ( p2_u3311,n10040 );
   buf U9669 ( p2_u3328,n19188 );
   nand U9670 ( n19188,n11401,n11402,n11403,n11404 );
   nand U9671 ( n10043,n11145,p2_d_reg_18_ );
   not U9672 ( p2_u3310,n10043 );
   buf U9673 ( p2_u3329,n19187 );
   nand U9674 ( n19187,n11391,n11392,n11393,n11394 );
   nand U9675 ( n10046,n11145,p2_d_reg_19_ );
   not U9676 ( p2_u3309,n10046 );
   buf U9677 ( p2_u3330,n19186 );
   nand U9678 ( n19186,n11381,n11382,n11383,n11384 );
   nand U9679 ( n10049,n11145,p2_d_reg_20_ );
   not U9680 ( p2_u3308,n10049 );
   buf U9681 ( p2_u3331,n19185 );
   nand U9682 ( n19185,n11372,n11373,n11374,n11375 );
   nand U9683 ( n10052,n11145,p2_d_reg_21_ );
   not U9684 ( p2_u3307,n10052 );
   buf U9685 ( p2_u3333,n19183 );
   nand U9686 ( n19183,n11355,n11356,n11357,n11358 );
   nand U9687 ( n10055,n11145,p2_d_reg_22_ );
   not U9688 ( p2_u3306,n10055 );
   buf U9689 ( p2_u3334,n19182 );
   nand U9690 ( n19182,n11346,n11347,n11348,n11349 );
   nand U9691 ( n10058,n11145,p2_d_reg_23_ );
   not U9692 ( p2_u3305,n10058 );
   buf U9693 ( p2_u3336,n19180 );
   nand U9694 ( n19180,n11329,n11330,n11331,n11332 );
   nand U9695 ( n10061,n11145,p2_d_reg_24_ );
   not U9696 ( p2_u3304,n10061 );
   buf U9697 ( p2_u3337,n19179 );
   nand U9698 ( n19179,n11320,n11321,n11322,n11323 );
   buf U9699 ( p2_u3296,n19275 );
   nand U9700 ( n19275,n11438,n11439,n11440,n11441 );
   nand U9701 ( n11439,n11458,n11125 );
   buf U9702 ( p2_u3340,n19176 );
   nand U9703 ( n19176,n11296,n11297,n11298,n11299 );
   buf U9704 ( p2_u3288,n19283 );
   nand U9705 ( n19283,n11645,n11646,n11647,n11648 );
   nor U9706 ( n11648,n11649,n11650,n11651,n11652 );
   buf U9707 ( p2_u3341,n19175 );
   nand U9708 ( n19175,n11286,n11287,n11288,n11289 );
   not U9709 ( p2_u3286,n10068 );
   not U9710 ( n10069,n11706 );
   nor U9711 ( n10068,n9964,n10005 );
   or U9712 ( n11706,n11456,n11006 );
   buf U9713 ( p2_u3342,n19174 );
   nand U9714 ( n19174,n11279,n11280,n11281,n11282 );
   not U9715 ( p2_u3285,n10071 );
   not U9716 ( n10072,n11747 );
   nor U9717 ( n10071,n9965,n10006 );
   or U9718 ( n11747,n11456,n10997 );
   buf U9719 ( p2_u3343,n19173 );
   nand U9720 ( n19173,n11269,n11270,n11271,n11272 );
   buf U9721 ( p2_u3284,n19285 );
   nand U9722 ( n19285,n11785,n11786,n11787,n11788 );
   nor U9723 ( n11788,n11789,n11790,n11791,n11792 );
   buf U9724 ( p2_u3344,n19172 );
   nand U9725 ( n19172,n11262,n11263,n11264,n11265 );
   not U9726 ( p2_u3283,n10076 );
   not U9727 ( n10077,n11815 );
   nor U9728 ( n10076,n9966,n10001 );
   or U9729 ( n11815,n11456,n10975 );
   buf U9730 ( p2_u3345,n19171 );
   nand U9731 ( n19171,n11252,n11253,n11254,n11255 );
   not U9732 ( p2_u3282,n10079 );
   not U9733 ( n10080,n11849 );
   nor U9734 ( n10079,n9967,n10007 );
   or U9735 ( n11849,n11456,n10962 );
   buf U9736 ( p2_u3346,n19170 );
   nand U9737 ( n19170,n11245,n11246,n11247,n11248 );
   buf U9738 ( p2_u3280,n19287 );
   nand U9739 ( n19287,n11916,n11917,n11918,n11919 );
   nor U9740 ( n11919,n11920,n11921,n11922,n11923 );
   buf U9741 ( p2_u3347,n19169 );
   nand U9742 ( n19169,n11235,n11236,n11237,n11238 );
   not U9743 ( p2_u3278,n10084 );
   not U9744 ( n10085,n11996 );
   nor U9745 ( n10084,n9968,n10002 );
   or U9746 ( n11996,n11456,n10919 );
   buf U9747 ( p2_u3348,n19168 );
   nand U9748 ( n19168,n11228,n11229,n11230,n11231 );
   not U9749 ( p2_u3277,n10087 );
   nor U9750 ( n10087,n9969,n10003 );
   buf U9751 ( p2_u3349,n19167 );
   nand U9752 ( n19167,n11219,n11220,n11221,n11222 );
   not U9753 ( p2_u3276,n10089 );
   not U9754 ( n10090,n12047 );
   nor U9755 ( n10089,n9970,n10008 );
   or U9756 ( n12047,n11456,n10896 );
   buf U9757 ( p2_u3351,n19165 );
   nand U9758 ( n19165,n11203,n11204,n11205,n11206 );
   not U9759 ( p2_u3275,n10092 );
   not U9760 ( n10093,n12080 );
   nor U9761 ( n10092,n9971,n10009 );
   or U9762 ( n12080,n11456,n10887 );
   buf U9763 ( p2_u3353,n19163 );
   nand U9764 ( n19163,n11186,n11187,n11188,n11189 );
   buf U9765 ( p2_u3274,n19289 );
   nand U9766 ( n19289,n12122,n12123,n12124,n12125 );
   buf U9767 ( p2_u3355,n19161 );
   nand U9768 ( n19161,n11173,n11174,n11175,n11176 );
   not U9769 ( p2_u3273,n10097 );
   not U9770 ( n10098,n12156 );
   nor U9771 ( n10097,n9972,n10010 );
   or U9772 ( n12156,n11456,n10865 );
   buf U9773 ( p2_u3356,n19160 );
   nand U9774 ( n19160,n11166,n11167,n11168,n11169 );
   not U9775 ( p2_u3271,n10100 );
   not U9776 ( n10101,n12212 );
   nor U9777 ( n10100,n9973,n10004 );
   or U9778 ( n12212,n11456,n10840 );
   buf U9779 ( p2_u3357,n19159 );
   nand U9780 ( n19159,n11160,n11161,n11162,n11163 );
   not U9781 ( p2_u3270,n10103 );
   not U9782 ( n10104,n12236 );
   nor U9783 ( n10103,n9974,n10011 );
   or U9784 ( n12236,n11456,n10828 );
   buf U9785 ( p2_u3358,n19158 );
   nand U9786 ( n19158,n11151,n11152,n11153 );
   not U9787 ( p2_u3269,n10106 );
   not U9788 ( n10107,n12276 );
   nor U9789 ( n10106,n9975,n10012 );
   or U9790 ( n12276,n11456,n10819 );
   not U9791 ( p1_u3083,n16965 );
   nand U9792 ( n16965,n18784,n14496 );
   buf U9793 ( p2_u3267,n19292 );
   nand U9794 ( n19292,n12340,n12341,n12342,n12343 );
   nor U9795 ( n12343,n12344,n12345,n12346 );
   buf U9796 ( p1_u3211,n19156 );
   nand U9797 ( n19156,n18476,n18477,n18478,n18479 );
   buf U9798 ( p2_u3266,n19293 );
   nand U9799 ( n19293,n12508,n12509,n12510,n12511 );
   buf U9800 ( p1_u3215,n19152 );
   nand U9801 ( n19152,n17857,n17858,n17859,n17860 );
   or U9802 ( n17858,n17865,n17502 );
   buf U9803 ( p2_u3265,n19294 );
   nand U9804 ( n19294,n12514,n12515,n12516,n12511 );
   buf U9805 ( p1_u3216,n19151 );
   nand U9806 ( n19151,n17843,n17844,n17845,n17846 );
   buf U9807 ( p2_u3264,n19295 );
   nand U9808 ( n19295,n12532,n12533,n12534 );
   nor U9809 ( n12534,n12535,n12536,n12537 );
   buf U9810 ( p1_u3217,n19150 );
   nand U9811 ( n19150,n17830,n17831,n17832,n17833 );
   nand U9812 ( n17831,n17838,n17517 );
   buf U9813 ( p2_u3262,n19297 );
   nand U9814 ( n19297,n12596,n12597,n12598 );
   nor U9815 ( n12598,n12599,n12600,n12601 );
   buf U9816 ( p1_u3220,n19147 );
   nand U9817 ( n19147,n17757,n17758,n17759,n17760 );
   buf U9818 ( p2_u3258,n19301 );
   nand U9819 ( n19301,n12702,n12703,n12704 );
   nor U9820 ( n12704,n12705,n12706,n12707 );
   buf U9821 ( p1_u3222,n19145 );
   nand U9822 ( n19145,n17729,n17730,n17731,n17732 );
   buf U9823 ( p2_u3255,n19304 );
   nand U9824 ( n19304,n12788,n12789,n12790 );
   nor U9825 ( n12790,n12791,n12792,n12793 );
   buf U9826 ( p1_u3225,n19142 );
   nand U9827 ( n19142,n17687,n17688,n17689,n17690 );
   buf U9828 ( p2_u3253,n19306 );
   nand U9829 ( n19306,n12839,n12840,n12841 );
   nor U9830 ( n12841,n12842,n12843,n12844 );
   buf U9831 ( p1_u3226,n19141 );
   nand U9832 ( n19141,n17672,n17673,n17674,n17675 );
   nand U9833 ( n17673,n17680,n17681,n17517 );
   buf U9834 ( p2_u3247,n19312 );
   nand U9835 ( n19312,n13019,n13020,n13021 );
   nor U9836 ( n13021,n13022,n13023,n13024 );
   buf U9837 ( p1_u3229,n19138 );
   nand U9838 ( n19138,n17634,n17635,n17636,n17637 );
   buf U9839 ( p2_u3552,n19315 );
   nand U9840 ( n19315,n10661,n10662 );
   nand U9841 ( n10662,p2_datao_reg_0_,n10569 );
   buf U9842 ( p1_u3232,n19135 );
   nand U9843 ( n19135,n17596,n17597,n17598,n17599 );
   nand U9844 ( n17597,n17604,n17605,n17517 );
   buf U9845 ( p2_u3553,n19316 );
   nand U9846 ( n19316,n10658,n10659 );
   nand U9847 ( n10659,p2_datao_reg_1_,n10569 );
   buf U9848 ( p1_u3233,n19134 );
   nand U9849 ( n19134,n17582,n17583,n17584,n17585 );
   buf U9850 ( p2_u3554,n19317 );
   nand U9851 ( n19317,n10655,n10656 );
   nand U9852 ( n10656,p2_datao_reg_2_,n10569 );
   buf U9853 ( p1_u3237,n19130 );
   nand U9854 ( n19130,n17527,n17528,n17529,n17530 );
   buf U9855 ( p2_u3555,n19318 );
   nand U9856 ( n19318,n10652,n10653 );
   nand U9857 ( n10653,p2_datao_reg_3_,n10569 );
   buf U9858 ( p1_u3238,n19129 );
   nand U9859 ( n19129,n17508,n17509,n17510,n17511 );
   buf U9860 ( p2_u3556,n19319 );
   nand U9861 ( n19319,n10649,n10650 );
   nand U9862 ( n10650,p2_datao_reg_4_,n10569 );
   buf U9863 ( p1_u3239,n19128 );
   nand U9864 ( n19128,n17490,n17491,n17492,n17493 );
   or U9865 ( n17491,n17501,n17502 );
   buf U9866 ( p2_u3557,n19320 );
   nand U9867 ( n19320,n10646,n10647 );
   nand U9868 ( n10647,p2_datao_reg_5_,n10569 );
   buf U9869 ( p1_u3274,n19060 );
   nand U9870 ( n19060,n15882,n15883,n15884,n15885 );
   nor U9871 ( n15885,n15886,n15887,n15888,n15889 );
   buf U9872 ( p2_u3558,n19321 );
   nand U9873 ( n19321,n10643,n10644 );
   nand U9874 ( n10644,p2_datao_reg_6_,n10569 );
   buf U9875 ( p1_u3278,n19056 );
   nand U9876 ( n19056,n15754,n15755,n15756,n15757 );
   nor U9877 ( n15757,n15758,n15759,n15760,n15761 );
   buf U9878 ( p2_u3559,n19322 );
   nand U9879 ( n19322,n10640,n10641 );
   nand U9880 ( n10641,p2_datao_reg_7_,n10569 );
   buf U9881 ( p1_u3283,n19051 );
   nand U9882 ( n19051,n15590,n15591,n15592,n15593 );
   nor U9883 ( n15593,n15594,n15595,n15596,n15597 );
   buf U9884 ( p2_u3560,n19323 );
   nand U9885 ( n19323,n10637,n10638 );
   nand U9886 ( n10638,p2_datao_reg_8_,n10569 );
   buf U9887 ( p1_u3286,n19048 );
   nand U9888 ( n19048,n15473,n15474,n15475,n15476 );
   nor U9889 ( n15476,n15477,n15478,n15479,n15480 );
   buf U9890 ( p2_u3561,n19324 );
   nand U9891 ( n19324,n10634,n10635 );
   nand U9892 ( n10635,p2_datao_reg_9_,n10569 );
   buf U9893 ( p1_u3289,n19045 );
   nand U9894 ( n19045,n15388,n15389,n15390,n15391 );
   nor U9895 ( n15391,n15392,n15393,n15394,n15395 );
   buf U9896 ( p2_u3562,n19325 );
   nand U9897 ( n19325,n10631,n10632 );
   nand U9898 ( n10632,p2_datao_reg_10_,n10569 );
   nand U9899 ( n10147,n15069,p1_d_reg_31_ );
   not U9900 ( p1_u3292,n10147 );
   buf U9901 ( p2_u3563,n19326 );
   nand U9902 ( n19326,n10628,n10629 );
   nand U9903 ( n10629,p2_datao_reg_11_,n10569 );
   nand U9904 ( n10150,n15069,p1_d_reg_30_ );
   not U9905 ( p1_u3293,n10150 );
   buf U9906 ( p2_u3564,n19327 );
   nand U9907 ( n19327,n10625,n10626 );
   nand U9908 ( n10626,p2_datao_reg_12_,n10569 );
   buf U9909 ( p1_u3294,n18978 );
   nor U9910 ( n18978,n15070,n15347 );
   buf U9911 ( p2_u3565,n19328 );
   nand U9912 ( n19328,n10622,n10623 );
   nand U9913 ( n10623,p2_datao_reg_13_,n10569 );
   nand U9914 ( n10155,n15069,p1_d_reg_28_ );
   not U9915 ( p1_u3295,n10155 );
   buf U9916 ( p2_u3566,n19329 );
   nand U9917 ( n19329,n10619,n10620 );
   nand U9918 ( n10620,p2_datao_reg_14_,n10569 );
   buf U9919 ( p1_u3296,n18977 );
   nor U9920 ( n18977,n15070,n15346 );
   buf U9921 ( p2_u3567,n19330 );
   nand U9922 ( n19330,n10616,n10617 );
   nand U9923 ( n10617,p2_datao_reg_15_,n10569 );
   nand U9924 ( n10160,n15069,p1_d_reg_26_ );
   not U9925 ( p1_u3297,n10160 );
   buf U9926 ( p2_u3568,n19331 );
   nand U9927 ( n19331,n10613,n10614 );
   nand U9928 ( n10614,p2_datao_reg_16_,n10569 );
   nand U9929 ( n10163,n15069,p1_d_reg_25_ );
   not U9930 ( p1_u3298,n10163 );
   buf U9931 ( p2_u3569,n19332 );
   nand U9932 ( n19332,n10610,n10611 );
   nand U9933 ( n10611,p2_datao_reg_17_,n10569 );
   nand U9934 ( n10166,n15069,p1_d_reg_24_ );
   not U9935 ( p1_u3299,n10166 );
   buf U9936 ( p2_u3570,n19333 );
   nand U9937 ( n19333,n10607,n10608 );
   nand U9938 ( n10608,p2_datao_reg_18_,n10569 );
   nand U9939 ( n10169,n15069,p1_d_reg_23_ );
   not U9940 ( p1_u3300,n10169 );
   buf U9941 ( p2_u3571,n19334 );
   nand U9942 ( n19334,n10604,n10605 );
   nand U9943 ( n10605,p2_datao_reg_19_,n10569 );
   nand U9944 ( n10172,n15069,p1_d_reg_22_ );
   not U9945 ( p1_u3301,n10172 );
   buf U9946 ( p2_u3572,n19335 );
   nand U9947 ( n19335,n10601,n10602 );
   nand U9948 ( n10602,p2_datao_reg_20_,n10569 );
   nand U9949 ( n10175,n15069,p1_d_reg_21_ );
   not U9950 ( p1_u3302,n10175 );
   buf U9951 ( p2_u3573,n19336 );
   nand U9952 ( n19336,n10598,n10599 );
   nand U9953 ( n10599,p2_datao_reg_21_,n10569 );
   nand U9954 ( n10178,n15069,p1_d_reg_20_ );
   not U9955 ( p1_u3303,n10178 );
   buf U9956 ( p2_u3574,n19337 );
   nand U9957 ( n19337,n10595,n10596 );
   nand U9958 ( n10596,p2_datao_reg_22_,n10569 );
   buf U9959 ( p1_u3304,n18976 );
   nor U9960 ( n18976,n15070,n15345 );
   buf U9961 ( p2_u3575,n19338 );
   nand U9962 ( n19338,n10592,n10593 );
   nand U9963 ( n10593,p2_datao_reg_23_,n10569 );
   buf U9964 ( p1_u3305,n18975 );
   nor U9965 ( n18975,n15070,n15344 );
   buf U9966 ( p2_u3576,n19339 );
   nand U9967 ( n19339,n10589,n10590 );
   nand U9968 ( n10590,p2_datao_reg_24_,n10569 );
   buf U9969 ( p1_u3306,n18974 );
   nor U9970 ( n18974,n15070,n15343 );
   buf U9971 ( p2_u3577,n19340 );
   nand U9972 ( n19340,n10586,n10587 );
   nand U9973 ( n10587,p2_datao_reg_25_,n10569 );
   buf U9974 ( p1_u3307,n18973 );
   nor U9975 ( n18973,n15070,n15342 );
   buf U9976 ( p2_u3578,n19341 );
   nand U9977 ( n19341,n10583,n10584 );
   nand U9978 ( n10584,p2_datao_reg_26_,n10569 );
   nand U9979 ( n10189,n15069,p1_d_reg_15_ );
   not U9980 ( p1_u3308,n10189 );
   buf U9981 ( p2_u3579,n19342 );
   nand U9982 ( n19342,n10580,n10581 );
   nand U9983 ( n10581,p2_datao_reg_27_,n10569 );
   nand U9984 ( n10192,n15069,p1_d_reg_14_ );
   not U9985 ( p1_u3309,n10192 );
   buf U9986 ( p2_u3580,n19343 );
   nand U9987 ( n19343,n10577,n10578 );
   nand U9988 ( n10578,p2_datao_reg_28_,n10569 );
   buf U9989 ( p1_u3310,n18972 );
   nor U9990 ( n18972,n15070,n15341 );
   buf U9991 ( p2_u3581,n19344 );
   nand U9992 ( n19344,n10574,n10575 );
   nand U9993 ( n10575,p2_datao_reg_29_,n10569 );
   nand U9994 ( n10197,n15069,p1_d_reg_12_ );
   not U9995 ( p1_u3311,n10197 );
   buf U9996 ( p2_u3582,n19345 );
   nand U9997 ( n19345,n10571,n10572 );
   nand U9998 ( n10572,p2_datao_reg_30_,n10569 );
   nand U9999 ( n10200,n15069,p1_d_reg_11_ );
   not U10000 ( p1_u3312,n10200 );
   buf U10001 ( p2_u3583,n19346 );
   nand U10002 ( n19346,n10567,n10568 );
   nand U10003 ( n10568,p2_datao_reg_31_,n10569 );
   buf U10004 ( p1_u3313,n18971 );
   nor U10005 ( n18971,n15070,n15340 );
   buf U10006 ( p2_u3242,n19349 );
   nand U10007 ( n19349,n13582,n13583,n13584,n13585 );
   nand U10008 ( n10205,n15069,p1_d_reg_9_ );
   not U10009 ( p1_u3314,n10205 );
   buf U10010 ( p2_u3241,n19350 );
   nand U10011 ( n19350,n13606,n13607,n13608,n13609 );
   nand U10012 ( n10208,n15069,p1_d_reg_8_ );
   not U10013 ( p1_u3315,n10208 );
   buf U10014 ( p2_u3238,n19353 );
   nand U10015 ( n19353,n13651,n13652,n13653,n13654 );
   nand U10016 ( n10211,n15069,p1_d_reg_7_ );
   not U10017 ( p1_u3316,n10211 );
   buf U10018 ( p2_u3237,n19354 );
   nand U10019 ( n19354,n13671,n13672,n13673,n13674 );
   buf U10020 ( p1_u3317,n18970 );
   nor U10021 ( n18970,n15070,n15339 );
   buf U10022 ( p2_u3235,n19356 );
   nand U10023 ( n19356,n13703,n13704,n13705,n13706 );
   nand U10024 ( n10216,n15069,p1_d_reg_5_ );
   not U10025 ( p1_u3318,n10216 );
   buf U10026 ( p2_u3234,n19357 );
   nand U10027 ( n19357,n13717,n13718,n13719,n13720 );
   nand U10028 ( n10219,n15069,p1_d_reg_4_ );
   not U10029 ( p1_u3319,n10219 );
   buf U10030 ( p2_u3233,n19358 );
   nand U10031 ( n19358,n13730,n13731,n13732,n13733 );
   or U10032 ( n13731,n13737,n13576 );
   nand U10033 ( n10222,n15069,p1_d_reg_3_ );
   not U10034 ( p1_u3320,n10222 );
   buf U10035 ( p2_u3231,n19360 );
   nand U10036 ( n19360,n13754,n13755,n13756,n13757 );
   buf U10037 ( p1_u3321,n18969 );
   nor U10038 ( n18969,n15070,n15338 );
   not U10039 ( n15070,n15069 );
   buf U10040 ( p2_u3228,n19363 );
   nand U10041 ( n19363,n13797,n13798,n13799,n13800 );
   nand U10042 ( n13798,n13806,n13807,n13594 );
   buf U10043 ( u126,n18934 );
   xor U10044 ( n18934,n10565,p1_rd_reg );
   buf U10045 ( p2_u3226,n19365 );
   nand U10046 ( n19365,n13824,n13825,n13826,n13827 );
   buf U10047 ( add_1071_u46,n18933 );
   xor U10048 ( n18933,p2_addr_reg_0_,p1_addr_reg_0_ );
   buf U10049 ( p2_u3215,n19376 );
   nand U10050 ( n19376,n14298,n14299,n14300,n14301 );
   and U10051 ( n17827,n18694,n18695 );
   and U10052 ( n13906,n14439,n14438 );
   nor U10053 ( n15384,n15089,n14733 );
   not U10054 ( n11460,n11479 );
   nand U10055 ( n11145,n11436,n11437 );
   not U10056 ( n11146,n11145 );
   not U10057 ( n10790,n10773 );
   not U10058 ( n17013,n17012 );
   nor U10059 ( n17012,n16454,n16979 );
   not U10060 ( p2_u3966,n10569 );
   not U10061 ( n10569,n19378 );
   nor U10062 ( n19378,n13072,p2_u3152 );
   nand U10063 ( n16506,n16964,n16965 );
   not U10064 ( n12574,n12551 );
   not U10065 ( n16446,n16735 );
   buf U10066 ( p2_u3246,n19313 );
   nand U10067 ( n19313,n13037,n13038,n13039 );
   nor U10068 ( n13039,n13040,n13041,n13042 );
   buf U10069 ( p2_u3354,n19162 );
   nand U10070 ( n19162,n11179,n11180,n11181,n11182 );
   buf U10071 ( p2_u3224,n19367 );
   nand U10072 ( n19367,n13849,n13850,n13851,n13852 );
   buf U10073 ( p1_u3270,n19064 );
   nand U10074 ( n19064,n15993,n15994,n15995,n15996 );
   buf U10075 ( p1_u3290,n19044 );
   nand U10076 ( n19044,n15368,n15369,n15370,n15371 );
   nor U10077 ( n15371,n15372,n15373,n15374,n15375 );
   buf U10078 ( p2_u3295,n19276 );
   nand U10079 ( n19276,n11462,n11463,n11464,n11465 );
   nor U10080 ( n11465,n11466,n11467,n11468,n11469 );
   buf U10081 ( p1_u3231,n19136 );
   nand U10082 ( n19136,n17611,n17612,n17613,n17614 );
   buf U10083 ( p2_u3225,n19366 );
   nand U10084 ( n19366,n13834,n13835,n13836,n13837 );
   not U10085 ( n15376,n15088 );
   buf U10086 ( p2_u3352,n19164 );
   nand U10087 ( n19164,n11196,n11197,n11198,n11199 );
   buf U10088 ( p1_u3245,n19090 );
   nand U10089 ( n19090,n16842,n16843,n16844,n16845 );
   nand U10090 ( n16843,n16852,n16860 );
   nor U10091 ( n16845,n16846,n16847,n16848 );
   buf U10092 ( p2_u3261,n19298 );
   nand U10093 ( n19298,n12627,n12628,n12629,n12630 );
   nand U10094 ( n12630,n12612,n12631 );
   buf U10095 ( p1_u3268,n19066 );
   nand U10096 ( n19066,n16065,n16066,n16067,n16068 );
   nor U10097 ( n16068,n16069,n16070,n16071,n16072 );
   buf U10098 ( p1_u3277,n19057 );
   nand U10099 ( n19057,n15790,n15791,n15792,n15793 );
   nor U10100 ( n15793,n15794,n15795,n15796,n15797 );
   buf U10101 ( p1_u3219,n19148 );
   nand U10102 ( n19148,n17768,n17769,n17770,n17771 );
   buf U10103 ( p2_u3294,n19277 );
   nand U10104 ( n19277,n11482,n11483,n11484,n11485 );
   nor U10105 ( n11485,n11486,n11487,n11488,n11489 );
   buf U10106 ( p1_u3227,n19140 );
   nand U10107 ( n19140,n17659,n17660,n17661,n17662 );
   buf U10108 ( p2_u3227,n19364 );
   nand U10109 ( n19364,n13812,n13813,n13814,n13815 );
   buf U10110 ( p2_u3223,n19368 );
   nand U10111 ( n19368,n13860,n13861,n13862,n13863 );
   or U10112 ( n13861,n13868,n13576 );
   nor U10113 ( n11461,n10851,n11445 );
   buf U10114 ( p2_u3350,n19166 );
   nand U10115 ( n19166,n11212,n11213,n11214,n11215 );
   buf U10116 ( p1_u3267,n19067 );
   nand U10117 ( n19067,n16108,n16109,n16110,n16111 );
   buf U10118 ( p1_u3288,n19046 );
   nand U10119 ( n19046,n15424,n15425,n15426,n15427 );
   nor U10120 ( n15427,n15428,n15429,n15430,n15431 );
   buf U10121 ( p1_u3255,n19080 );
   nand U10122 ( n19080,n16579,n16580,n16581,n16582 );
   nand U10123 ( n16582,n16573,n16583 );
   buf U10124 ( p1_u3244,n19091 );
   nand U10125 ( n19091,n16872,n16873,n16874,n16875 );
   nand U10126 ( n16872,n16461,n16885 );
   buf U10127 ( p2_u3292,n19279 );
   nand U10128 ( n19279,n11538,n11539,n11540,n11541 );
   nor U10129 ( n11541,n11542,n11543,n11544,n11545 );
   buf U10130 ( p1_u3224,n19143 );
   nand U10131 ( n19143,n17699,n17700,n17701,n17702 );
   nand U10132 ( n17700,n17707,n17517 );
   buf U10133 ( p2_u3248,n19311 );
   nand U10134 ( n19311,n12986,n12987,n12988,n12989 );
   buf U10135 ( p2_u3243,n19348 );
   nand U10136 ( n19348,n13564,n13565,n13566,n13567 );
   buf U10137 ( p2_u3222,n19369 );
   nand U10138 ( n19369,n13873,n13874,n13875,n13876 );
   nand U10139 ( n13874,n13881,n13882,n13594 );
   not U10140 ( n11721,n11672 );
   buf U10141 ( p2_u3339,n19177 );
   nand U10142 ( n19177,n11306,n11307,n11308,n11309 );
   buf U10143 ( p1_u3285,n19049 );
   nand U10144 ( n19049,n15513,n15514,n15515,n15516 );
   nor U10145 ( n15516,n15517,n15518,n15519,n15520 );
   buf U10146 ( p1_u3266,n19068 );
   nand U10147 ( n19068,n16138,n16139,n16140,n16141 );
   buf U10148 ( p1_u3282,n19052 );
   nand U10149 ( n19052,n15628,n15629,n15630,n15631 );
   nor U10150 ( n15631,n15632,n15633,n15634,n15635 );
   buf U10151 ( p1_u3260,n19075 );
   nand U10152 ( n19075,n16435,n16436,n16437,n16438 );
   buf U10153 ( p2_u3293,n19278 );
   nand U10154 ( n19278,n11512,n11513,n11514,n11515 );
   nor U10155 ( n11515,n11516,n11517,n11518,n11519 );
   buf U10156 ( p2_u3232,n19359 );
   nand U10157 ( n19359,n13742,n13743,n13744,n13745 );
   buf U10158 ( p1_u3236,n19131 );
   nand U10159 ( n19131,n17541,n17542,n17543,n17544 );
   buf U10160 ( p1_u3223,n19144 );
   nand U10161 ( n19144,n17712,n17713,n17714,n17715 );
   buf U10162 ( p1_u3257,n19078 );
   nand U10163 ( n19078,n16530,n16531,n16532,n16533 );
   nand U10164 ( n16533,n16519,n16534 );
   buf U10165 ( p2_u3221,n19370 );
   nand U10166 ( n19370,n13909,n13910,n13911,n13912 );
   nand U10167 ( n13910,n13594,n13917 );
   buf U10168 ( p2_u3263,n19296 );
   nand U10169 ( n19296,n12565,n12566,n12567,n12568 );
   nand U10170 ( n12568,n12547,n12569 );
   nand U10171 ( n11630,n13209,n13153 );
   not U10172 ( n11722,n11676 );
   not U10173 ( n15491,n15616 );
   buf U10174 ( p2_u3338,n19178 );
   nand U10175 ( n19178,n11313,n11314,n11315,n11316 );
   buf U10176 ( p2_u3239,n19352 );
   nand U10177 ( n19352,n13635,n13636,n13637,n13638 );
   buf U10178 ( p1_u3284,n19050 );
   nand U10179 ( n19050,n15550,n15551,n15552,n15553 );
   nor U10180 ( n15553,n15554,n15555,n15556,n15557 );
   buf U10181 ( p1_u3264,n19070 );
   nand U10182 ( n19070,n16208,n16209,n16210,n16211 );
   buf U10183 ( p1_u3276,n19058 );
   nand U10184 ( n19058,n15815,n15816,n15817,n15818 );
   nor U10185 ( n15818,n15819,n15820,n15821,n15822 );
   buf U10186 ( p1_u3258,n19077 );
   nand U10187 ( n19077,n16500,n16501,n16502,n16503 );
   buf U10188 ( p2_u3290,n19281 );
   nand U10189 ( n19281,n11588,n11589,n11590,n11591 );
   nor U10190 ( n11591,n11592,n11593,n11594,n11595 );
   buf U10191 ( p1_u3252,n19083 );
   nand U10192 ( n19083,n16654,n16655,n16656,n16657 );
   nand U10193 ( n16657,n16644,n16658 );
   buf U10194 ( p1_u3235,n19132 );
   nand U10195 ( n19132,n17555,n17556,n17557,n17558 );
   buf U10196 ( p1_u3221,n19146 );
   nand U10197 ( n19146,n17742,n17743,n17744,n17745 );
   buf U10198 ( p2_u3217,n19374 );
   nand U10199 ( n19374,n13970,n13971,n13972,n13973 );
   nand U10200 ( n13971,n13594,n13979 );
   buf U10201 ( p2_u3259,n19300 );
   nand U10202 ( n19300,n12676,n12677,n12678,n12679 );
   not U10203 ( n11631,n11724 );
   nor U10204 ( n16427,n16913,n16426 );
   not U10205 ( n15404,n15573 );
   nor U10206 ( n10808,n12366,n12520 );
   not U10207 ( n14699,n14756 );
   buf U10208 ( p2_u3335,n19181 );
   nand U10209 ( n19181,n11339,n11340,n11341,n11342 );
   buf U10210 ( p1_u3262,n19073 );
   nand U10211 ( n19073,n16414,n16415,n16416,n16417 );
   buf U10212 ( p1_u3275,n19059 );
   nand U10213 ( n19059,n15838,n15839,n15840,n15841 );
   nor U10214 ( n15841,n15842,n15843,n15844,n15845 );
   buf U10215 ( p2_u3281,n19286 );
   nand U10216 ( n19286,n11885,n11886,n11887,n11888 );
   or U10217 ( n11886,n11460,n10952 );
   nor U10218 ( n11888,n11889,n11890,n11891,n11892 );
   buf U10219 ( p1_u3254,n19081 );
   nand U10220 ( n19081,n16604,n16605,n16606,n16607 );
   buf U10221 ( p1_u3287,n19047 );
   nand U10222 ( n19047,n15448,n15449,n15450,n15451 );
   nor U10223 ( n15451,n15452,n15453,n15454,n15455 );
   buf U10224 ( p1_u3281,n19053 );
   nand U10225 ( n19053,n15648,n15649,n15650,n15651 );
   nor U10226 ( n15651,n15652,n15653,n15654,n15655 );
   buf U10227 ( p2_u3289,n19282 );
   nand U10228 ( n19282,n11615,n11616,n11617,n11618 );
   nor U10229 ( n11618,n11619,n11620,n11621,n11622 );
   buf U10230 ( p1_u3218,n19149 );
   nand U10231 ( n19149,n17780,n17781,n17782,n17783 );
   nand U10232 ( n17781,n17788,n17789,n17517 );
   buf U10233 ( p2_u3219,n19372 );
   nand U10234 ( n19372,n13944,n13945,n13946,n13947 );
   buf U10235 ( p2_u3216,n19375 );
   nand U10236 ( n19375,n13984,n13985,n13986,n13987 );
   buf U10237 ( p1_u3259,n19076 );
   nand U10238 ( n19076,n16470,n16471,n16472,n16473 );
   nand U10239 ( n16473,n16458,n16474 );
   buf U10240 ( p2_u3256,n19303 );
   nand U10241 ( n19303,n12759,n12760,n12761,n12762 );
   nand U10242 ( n12762,n12750,n12763 );
   not U10243 ( n15403,n15437 );
   nor U10244 ( n17399,n18695,n18696 );
   nor U10245 ( n13550,n14440,n14438 );
   nand U10246 ( n11629,n12349,n11132 );
   not U10247 ( n10792,n10805 );
   buf U10248 ( p2_u3327,n19189 );
   nand U10249 ( n19189,n11411,n11412,n11413 );
   nand U10250 ( n11411,n11415,n11158 );
   buf U10251 ( p1_u3454,n18979 );
   nand U10252 ( n18979,n15049,n15050 );
   nand U10253 ( n15050,n14693,n14688 );
   buf U10254 ( p1_u3457,n18980 );
   nand U10255 ( n18980,n15037,n15038 );
   nand U10256 ( n15038,n14693,n14685 );
   buf U10257 ( p1_u3460,n18981 );
   nand U10258 ( n18981,n15025,n15026 );
   nand U10259 ( n15026,n14693,n14682 );
   buf U10260 ( p1_u3463,n18982 );
   nand U10261 ( n18982,n15014,n15015 );
   nand U10262 ( n15015,n14693,n14679 );
   buf U10263 ( p1_u3466,n18983 );
   nand U10264 ( n18983,n15003,n15004 );
   nand U10265 ( n15004,n14693,n14676 );
   buf U10266 ( p1_u3469,n18984 );
   nand U10267 ( n18984,n14991,n14992 );
   nand U10268 ( n14992,n14693,n14673 );
   buf U10269 ( p1_u3472,n18985 );
   nand U10270 ( n18985,n14979,n14980 );
   nand U10271 ( n14980,n14693,n14670 );
   buf U10272 ( p1_u3475,n18986 );
   nand U10273 ( n18986,n14967,n14968 );
   nand U10274 ( n14968,n14693,n14667 );
   buf U10275 ( p1_u3478,n18987 );
   nand U10276 ( n18987,n14955,n14956 );
   nand U10277 ( n14956,n14693,n14664 );
   buf U10278 ( p1_u3481,n18988 );
   nand U10279 ( n18988,n14944,n14945 );
   nand U10280 ( n14945,n14693,n14661 );
   buf U10281 ( p1_u3484,n18989 );
   nand U10282 ( n18989,n14933,n14934 );
   nand U10283 ( n14934,n14693,n14658 );
   buf U10284 ( p1_u3487,n18990 );
   nand U10285 ( n18990,n14921,n14922 );
   nand U10286 ( n14922,n14693,n14655 );
   buf U10287 ( p1_u3490,n18991 );
   nand U10288 ( n18991,n14910,n14911 );
   nand U10289 ( n14911,n14693,n14652 );
   buf U10290 ( p1_u3493,n18992 );
   nand U10291 ( n18992,n14898,n14899 );
   nand U10292 ( n14899,n14693,n14649 );
   buf U10293 ( p1_u3496,n18993 );
   nand U10294 ( n18993,n14887,n14888 );
   nand U10295 ( n14888,n14693,n14646 );
   buf U10296 ( p1_u3499,n18994 );
   nand U10297 ( n18994,n14876,n14877 );
   nand U10298 ( n14877,n14693,n14643 );
   buf U10299 ( p1_u3502,n18995 );
   nand U10300 ( n18995,n14865,n14866 );
   nand U10301 ( n14866,n14693,n14640 );
   buf U10302 ( p1_u3505,n18996 );
   nand U10303 ( n18996,n14853,n14854 );
   nand U10304 ( n14854,n14693,n14637 );
   buf U10305 ( p1_u3508,n18997 );
   nand U10306 ( n18997,n14842,n14843 );
   nand U10307 ( n14843,n14693,n14634 );
   buf U10308 ( p1_u3510,n18998 );
   nand U10309 ( n18998,n14831,n14832 );
   nand U10310 ( n14832,n14693,n14631 );
   buf U10311 ( p1_u3511,n18999 );
   nand U10312 ( n18999,n14820,n14821 );
   nand U10313 ( n14821,n14693,n14628 );
   buf U10314 ( p1_u3512,n19000 );
   nand U10315 ( n19000,n14808,n14809 );
   nand U10316 ( n14809,n14693,n14625 );
   buf U10317 ( p1_u3513,n19001 );
   nand U10318 ( n19001,n14795,n14796 );
   nand U10319 ( n14796,n14693,n14622 );
   buf U10320 ( p1_u3514,n19002 );
   nand U10321 ( n19002,n14783,n14784 );
   nand U10322 ( n14784,n14693,n14619 );
   buf U10323 ( p1_u3515,n19003 );
   nand U10324 ( n19003,n14772,n14773 );
   nand U10325 ( n14773,n14693,n14616 );
   buf U10326 ( p1_u3516,n19004 );
   nand U10327 ( n19004,n14760,n14761 );
   nand U10328 ( n14761,n14693,n14613 );
   buf U10329 ( p1_u3517,n19005 );
   nand U10330 ( n19005,n14747,n14748 );
   nand U10331 ( n14748,n14693,n14610 );
   buf U10332 ( p1_u3518,n19006 );
   nand U10333 ( n19006,n14735,n14736 );
   nand U10334 ( n14736,n14693,n14607 );
   buf U10335 ( p1_u3519,n19007 );
   nand U10336 ( n19007,n14721,n14722 );
   nand U10337 ( n14722,n14693,n14604 );
   buf U10338 ( p1_u3520,n19008 );
   nand U10339 ( n19008,n14710,n14711 );
   nand U10340 ( n14711,n14693,n14601 );
   buf U10341 ( p1_u3521,n19009 );
   nand U10342 ( n19009,n14702,n14703 );
   nand U10343 ( n14703,n14693,n14598 );
   buf U10344 ( p1_u3522,n19010 );
   nand U10345 ( n19010,n14691,n14692 );
   nand U10346 ( n14692,n14693,n14594 );
   buf U10347 ( p1_u3440,n18967 );
   nand U10348 ( n18967,n15072,n15073 );
   nand U10349 ( n15073,p1_d_reg_0_,n15069 );
   buf U10350 ( p1_u3565,n19105 );
   nand U10351 ( n19105,n14558,n14559 );
   nand U10352 ( n14559,p1_datao_reg_10_,n14496 );
   buf U10353 ( p1_u3567,n19107 );
   nand U10354 ( n19107,n14552,n14553 );
   nand U10355 ( n14553,p1_datao_reg_12_,n14496 );
   buf U10356 ( p1_u3574,n19114 );
   nand U10357 ( n19114,n14531,n14532 );
   nand U10358 ( n14532,p1_datao_reg_19_,n14496 );
   buf U10359 ( p1_u3576,n19116 );
   nand U10360 ( n19116,n14525,n14526 );
   nand U10361 ( n14526,p1_datao_reg_21_,n14496 );
   buf U10362 ( p1_u3584,n19124 );
   nand U10363 ( n19124,n14501,n14502 );
   nand U10364 ( n14502,p1_datao_reg_29_,n14496 );
   buf U10365 ( p2_u3332,n19184 );
   nand U10366 ( n19184,n11365,n11366,n11367,n11368 );
   buf U10367 ( p1_u3261,n19074 );
   nand U10368 ( n19074,n16419,n16420,n16416,n16421 );
   buf U10369 ( p1_u3265,n19069 );
   nand U10370 ( n19069,n16164,n16165,n16166,n16167 );
   buf U10371 ( p2_u3279,n19288 );
   nand U10372 ( n19288,n11961,n11962,n11963,n11964 );
   or U10373 ( n11962,n11460,n10930 );
   nor U10374 ( n11964,n11965,n11966,n11967,n11968 );
   buf U10375 ( p1_u3272,n19062 );
   nand U10376 ( n19062,n15937,n15938,n15939,n15940 );
   buf U10377 ( p1_u3279,n19055 );
   nand U10378 ( n19055,n15734,n15735,n15736,n15737 );
   nor U10379 ( n15737,n15738,n15739,n15740,n15741 );
   buf U10380 ( p1_u3251,n19084 );
   nand U10381 ( n19084,n16678,n16679,n16680,n16681 );
   buf U10382 ( p2_u3229,n19362 );
   nand U10383 ( n19362,n13785,n13786,n13787,n13788 );
   buf U10384 ( p2_u3287,n19284 );
   nand U10385 ( n19284,n11683,n11684,n11685,n11686 );
   nor U10386 ( n11686,n11687,n11688,n11689,n11690 );
   buf U10387 ( p1_u3228,n19139 );
   nand U10388 ( n19139,n17646,n17647,n17648,n17649 );
   or U10389 ( n17646,n17654,n17502 );
   buf U10390 ( p1_u3212,n19155 );
   nand U10391 ( n19155,n17896,n17897,n17898,n17899 );
   buf U10392 ( p2_u3236,n19355 );
   nand U10393 ( n19355,n13685,n13686,n13687,n13688 );
   nand U10394 ( n13686,n13693,n13694,n13594 );
   buf U10395 ( p1_u3256,n19079 );
   nand U10396 ( n19079,n16554,n16555,n16556,n16557 );
   nand U10397 ( n16557,n16558,n16559 );
   buf U10398 ( p2_u3260,n19299 );
   nand U10399 ( n19299,n12651,n12652,n12653,n12654 );
   nand U10400 ( n12654,n12655,n12656 );
   not U10401 ( n11670,n11477 );
   not U10402 ( n15493,n15572 );
   nor U10403 ( n14057,n11416,n12521 );
   nor U10404 ( n14059,n11414,n12521 );
   nor U10405 ( n12521,n12520,n13068 );
   not U10406 ( n11632,n12329 );
   nor U10407 ( n17398,n18695,n18694 );
   nor U10408 ( n13549,n14438,n14439 );
   nand U10409 ( n17811,n18339,n18687 );
   nand U10410 ( n11459,n12526,n11455 );
   nor U10411 ( n11157,n11156,p2_u3152 );
   buf U10412 ( p1_u3322,n18966 );
   nand U10413 ( n18966,n15335,n15336,n15337 );
   buf U10414 ( p1_u3554,n19042 );
   nand U10415 ( n19042,n14591,n14592 );
   nand U10416 ( n14592,n14593,n14594 );
   buf U10417 ( p2_u3551,n19274 );
   nand U10418 ( n19274,n10664,n10665 );
   buf U10419 ( p1_u3441,n18968 );
   nand U10420 ( n18968,n15067,n15068 );
   nand U10421 ( n15068,p1_d_reg_1_,n15069 );
   buf U10422 ( p1_u3523,n19011 );
   nand U10423 ( n19011,n14686,n14687 );
   buf U10424 ( p1_u3524,n19012 );
   nand U10425 ( n19012,n14683,n14684 );
   buf U10426 ( p1_u3525,n19013 );
   nand U10427 ( n19013,n14680,n14681 );
   buf U10428 ( p1_u3526,n19014 );
   nand U10429 ( n19014,n14677,n14678 );
   buf U10430 ( p1_u3527,n19015 );
   nand U10431 ( n19015,n14674,n14675 );
   buf U10432 ( p1_u3528,n19016 );
   nand U10433 ( n19016,n14671,n14672 );
   buf U10434 ( p1_u3529,n19017 );
   nand U10435 ( n19017,n14668,n14669 );
   buf U10436 ( p1_u3530,n19018 );
   nand U10437 ( n19018,n14665,n14666 );
   buf U10438 ( p1_u3531,n19019 );
   nand U10439 ( n19019,n14662,n14663 );
   buf U10440 ( p1_u3532,n19020 );
   nand U10441 ( n19020,n14659,n14660 );
   buf U10442 ( p1_u3533,n19021 );
   nand U10443 ( n19021,n14656,n14657 );
   buf U10444 ( p1_u3534,n19022 );
   nand U10445 ( n19022,n14653,n14654 );
   buf U10446 ( p1_u3535,n19023 );
   nand U10447 ( n19023,n14650,n14651 );
   buf U10448 ( p1_u3536,n19024 );
   nand U10449 ( n19024,n14647,n14648 );
   buf U10450 ( p1_u3537,n19025 );
   nand U10451 ( n19025,n14644,n14645 );
   buf U10452 ( p1_u3538,n19026 );
   nand U10453 ( n19026,n14641,n14642 );
   buf U10454 ( p1_u3539,n19027 );
   nand U10455 ( n19027,n14638,n14639 );
   buf U10456 ( p1_u3540,n19028 );
   nand U10457 ( n19028,n14635,n14636 );
   buf U10458 ( p1_u3541,n19029 );
   nand U10459 ( n19029,n14632,n14633 );
   buf U10460 ( p1_u3542,n19030 );
   nand U10461 ( n19030,n14629,n14630 );
   buf U10462 ( p1_u3543,n19031 );
   nand U10463 ( n19031,n14626,n14627 );
   buf U10464 ( p1_u3544,n19032 );
   nand U10465 ( n19032,n14623,n14624 );
   buf U10466 ( p1_u3545,n19033 );
   nand U10467 ( n19033,n14620,n14621 );
   buf U10468 ( p1_u3546,n19034 );
   nand U10469 ( n19034,n14617,n14618 );
   buf U10470 ( p1_u3547,n19035 );
   nand U10471 ( n19035,n14614,n14615 );
   buf U10472 ( p1_u3548,n19036 );
   nand U10473 ( n19036,n14611,n14612 );
   buf U10474 ( p1_u3549,n19037 );
   nand U10475 ( n19037,n14608,n14609 );
   buf U10476 ( p1_u3550,n19038 );
   nand U10477 ( n19038,n14605,n14606 );
   buf U10478 ( p1_u3551,n19039 );
   nand U10479 ( n19039,n14602,n14603 );
   buf U10480 ( p1_u3552,n19040 );
   nand U10481 ( n19040,n14599,n14600 );
   buf U10482 ( p1_u3553,n19041 );
   nand U10483 ( n19041,n14596,n14597 );
   buf U10484 ( p1_u3555,n19095 );
   nand U10485 ( n19095,n14588,n14589 );
   nand U10486 ( n14589,p1_datao_reg_0_,n14496 );
   buf U10487 ( p1_u3556,n19096 );
   nand U10488 ( n19096,n14585,n14586 );
   nand U10489 ( n14586,p1_datao_reg_1_,n14496 );
   buf U10490 ( p1_u3557,n19097 );
   nand U10491 ( n19097,n14582,n14583 );
   nand U10492 ( n14583,p1_datao_reg_2_,n14496 );
   buf U10493 ( p1_u3558,n19098 );
   nand U10494 ( n19098,n14579,n14580 );
   nand U10495 ( n14580,p1_datao_reg_3_,n14496 );
   buf U10496 ( p1_u3559,n19099 );
   nand U10497 ( n19099,n14576,n14577 );
   nand U10498 ( n14577,p1_datao_reg_4_,n14496 );
   buf U10499 ( p1_u3560,n19100 );
   nand U10500 ( n19100,n14573,n14574 );
   nand U10501 ( n14574,p1_datao_reg_5_,n14496 );
   buf U10502 ( p1_u3561,n19101 );
   nand U10503 ( n19101,n14570,n14571 );
   nand U10504 ( n14571,p1_datao_reg_6_,n14496 );
   buf U10505 ( p1_u3562,n19102 );
   nand U10506 ( n19102,n14567,n14568 );
   nand U10507 ( n14568,p1_datao_reg_7_,n14496 );
   buf U10508 ( p1_u3563,n19103 );
   nand U10509 ( n19103,n14564,n14565 );
   nand U10510 ( n14565,p1_datao_reg_8_,n14496 );
   buf U10511 ( p1_u3564,n19104 );
   nand U10512 ( n19104,n14561,n14562 );
   nand U10513 ( n14562,p1_datao_reg_9_,n14496 );
   buf U10514 ( p1_u3566,n19106 );
   nand U10515 ( n19106,n14555,n14556 );
   nand U10516 ( n14556,p1_datao_reg_11_,n14496 );
   buf U10517 ( p1_u3568,n19108 );
   nand U10518 ( n19108,n14549,n14550 );
   nand U10519 ( n14550,p1_datao_reg_13_,n14496 );
   buf U10520 ( p1_u3569,n19109 );
   nand U10521 ( n19109,n14546,n14547 );
   nand U10522 ( n14547,p1_datao_reg_14_,n14496 );
   buf U10523 ( p1_u3570,n19110 );
   nand U10524 ( n19110,n14543,n14544 );
   nand U10525 ( n14544,p1_datao_reg_15_,n14496 );
   buf U10526 ( p1_u3571,n19111 );
   nand U10527 ( n19111,n14540,n14541 );
   nand U10528 ( n14541,p1_datao_reg_16_,n14496 );
   buf U10529 ( p1_u3572,n19112 );
   nand U10530 ( n19112,n14537,n14538 );
   nand U10531 ( n14538,p1_datao_reg_17_,n14496 );
   buf U10532 ( p1_u3573,n19113 );
   nand U10533 ( n19113,n14534,n14535 );
   nand U10534 ( n14535,p1_datao_reg_18_,n14496 );
   buf U10535 ( p1_u3575,n19115 );
   nand U10536 ( n19115,n14528,n14529 );
   nand U10537 ( n14529,p1_datao_reg_20_,n14496 );
   buf U10538 ( p1_u3577,n19117 );
   nand U10539 ( n19117,n14522,n14523 );
   nand U10540 ( n14523,p1_datao_reg_22_,n14496 );
   buf U10541 ( p1_u3578,n19118 );
   nand U10542 ( n19118,n14519,n14520 );
   nand U10543 ( n14520,p1_datao_reg_23_,n14496 );
   buf U10544 ( p1_u3579,n19119 );
   nand U10545 ( n19119,n14516,n14517 );
   nand U10546 ( n14517,p1_datao_reg_24_,n14496 );
   buf U10547 ( p1_u3580,n19120 );
   nand U10548 ( n19120,n14513,n14514 );
   nand U10549 ( n14514,p1_datao_reg_25_,n14496 );
   buf U10550 ( p1_u3581,n19121 );
   nand U10551 ( n19121,n14510,n14511 );
   nand U10552 ( n14511,p1_datao_reg_26_,n14496 );
   buf U10553 ( p1_u3582,n19122 );
   nand U10554 ( n19122,n14507,n14508 );
   nand U10555 ( n14508,p1_datao_reg_27_,n14496 );
   buf U10556 ( p1_u3583,n19123 );
   nand U10557 ( n19123,n14504,n14505 );
   nand U10558 ( n14505,p1_datao_reg_28_,n14496 );
   buf U10559 ( p1_u3585,n19125 );
   nand U10560 ( n19125,n14498,n14499 );
   nand U10561 ( n14499,p1_datao_reg_30_,n14496 );
   buf U10562 ( p1_u3586,n19126 );
   nand U10563 ( n19126,n14494,n14495 );
   nand U10564 ( n14495,p1_datao_reg_31_,n14496 );
   buf U10565 ( p2_u3520,n19243 );
   nand U10566 ( n19243,n10759,n10760 );
   nand U10567 ( n10760,p2_reg1_reg_0_,n10668 );
   buf U10568 ( p2_u3521,n19244 );
   nand U10569 ( n19244,n10756,n10757 );
   nand U10570 ( n10757,p2_reg1_reg_1_,n10668 );
   buf U10571 ( p2_u3522,n19245 );
   nand U10572 ( n19245,n10753,n10754 );
   nand U10573 ( n10754,p2_reg1_reg_2_,n10668 );
   buf U10574 ( p2_u3523,n19246 );
   nand U10575 ( n19246,n10750,n10751 );
   nand U10576 ( n10751,p2_reg1_reg_3_,n10668 );
   buf U10577 ( p2_u3524,n19247 );
   nand U10578 ( n19247,n10747,n10748 );
   buf U10579 ( p2_u3525,n19248 );
   nand U10580 ( n19248,n10744,n10745 );
   buf U10581 ( p2_u3526,n19249 );
   nand U10582 ( n19249,n10741,n10742 );
   buf U10583 ( p2_u3527,n19250 );
   nand U10584 ( n19250,n10738,n10739 );
   buf U10585 ( p2_u3528,n19251 );
   nand U10586 ( n19251,n10735,n10736 );
   buf U10587 ( p2_u3529,n19252 );
   nand U10588 ( n19252,n10732,n10733 );
   buf U10589 ( p2_u3530,n19253 );
   nand U10590 ( n19253,n10729,n10730 );
   buf U10591 ( p2_u3531,n19254 );
   nand U10592 ( n19254,n10726,n10727 );
   buf U10593 ( p2_u3532,n19255 );
   nand U10594 ( n19255,n10723,n10724 );
   buf U10595 ( p2_u3533,n19256 );
   nand U10596 ( n19256,n10720,n10721 );
   buf U10597 ( p2_u3534,n19257 );
   nand U10598 ( n19257,n10717,n10718 );
   buf U10599 ( p2_u3535,n19258 );
   nand U10600 ( n19258,n10714,n10715 );
   buf U10601 ( p2_u3536,n19259 );
   nand U10602 ( n19259,n10711,n10712 );
   buf U10603 ( p2_u3537,n19260 );
   nand U10604 ( n19260,n10708,n10709 );
   buf U10605 ( p2_u3538,n19261 );
   nand U10606 ( n19261,n10705,n10706 );
   buf U10607 ( p2_u3539,n19262 );
   nand U10608 ( n19262,n10702,n10703 );
   buf U10609 ( p2_u3540,n19263 );
   nand U10610 ( n19263,n10699,n10700 );
   buf U10611 ( p2_u3541,n19264 );
   nand U10612 ( n19264,n10696,n10697 );
   buf U10613 ( p2_u3542,n19265 );
   nand U10614 ( n19265,n10693,n10694 );
   buf U10615 ( p2_u3543,n19266 );
   nand U10616 ( n19266,n10690,n10691 );
   buf U10617 ( p2_u3544,n19267 );
   nand U10618 ( n19267,n10687,n10688 );
   buf U10619 ( p2_u3545,n19268 );
   nand U10620 ( n19268,n10684,n10685 );
   buf U10621 ( p2_u3546,n19269 );
   nand U10622 ( n19269,n10681,n10682 );
   buf U10623 ( p2_u3547,n19270 );
   nand U10624 ( n19270,n10678,n10679 );
   buf U10625 ( p2_u3548,n19271 );
   nand U10626 ( n19271,n10675,n10676 );
   buf U10627 ( p2_u3549,n19272 );
   nand U10628 ( n19272,n10672,n10673 );
   buf U10629 ( p2_u3550,n19273 );
   nand U10630 ( n19273,n10669,n10670 );
   buf U10631 ( p1_u3352,n18936 );
   nand U10632 ( n18936,n15131,n15132,n15133,n15134 );
   buf U10633 ( p1_u3353,n18935 );
   nand U10634 ( n18935,n15123,n15124,n15125 );
   nand U10635 ( n15124,p1_ir_reg_0_,n15127 );
   buf U10636 ( p1_u3350,n18938 );
   nand U10637 ( n18938,n15142,n15143,n15144,n15145 );
   buf U10638 ( p1_u3344,n18944 );
   nand U10639 ( n18944,n15182,n15183,n15184,n15185 );
   buf U10640 ( p1_u3343,n18945 );
   nand U10641 ( n18945,n15187,n15188,n15189,n15190 );
   buf U10642 ( p1_u3342,n18946 );
   nand U10643 ( n18946,n15193,n15194,n15195,n15196 );
   buf U10644 ( p1_u3339,n18949 );
   nand U10645 ( n18949,n15212,n15213,n15214,n15215 );
   buf U10646 ( p1_u3351,n18937 );
   nand U10647 ( n18937,n15136,n15137,n15138,n15139 );
   buf U10648 ( p1_u3349,n18939 );
   nand U10649 ( n18939,n15147,n15148,n15149,n15150 );
   buf U10650 ( p1_u3347,n18941 );
   nand U10651 ( n18941,n15162,n15163,n15164,n15165 );
   buf U10652 ( p1_u3345,n18943 );
   nand U10653 ( n18943,n15176,n15177,n15178,n15179 );
   buf U10654 ( p1_u3341,n18947 );
   nand U10655 ( n18947,n15198,n15199,n15200,n15201 );
   buf U10656 ( p1_u3337,n18951 );
   nand U10657 ( n18951,n15227,n15228,n15229,n15230 );
   buf U10658 ( p1_u3334,n18954 );
   nand U10659 ( n18954,n15250,n15251,n15252,n15253 );
   buf U10660 ( p1_u3333,n18955 );
   nand U10661 ( n18955,n15256,n15257,n15258,n15259 );
   buf U10662 ( p1_u3331,n18957 );
   nand U10663 ( n18957,n15270,n15271,n15272,n15273 );
   buf U10664 ( p1_u3329,n18959 );
   nand U10665 ( n18959,n15284,n15285,n15286,n15287 );
   buf U10666 ( p1_u3327,n18961 );
   nand U10667 ( n18961,n15298,n15299,n15300,n15301 );
   buf U10668 ( p1_u3325,n18963 );
   nand U10669 ( n18963,n15312,n15313,n15314,n15315 );
   buf U10670 ( p1_u3263,n19071 );
   nand U10671 ( n19071,n16254,n16255,n16256,n16257 );
   buf U10672 ( p2_u3291,n19280 );
   nand U10673 ( n19280,n11563,n11564,n11565,n11566 );
   or U10674 ( n11564,n11460,n11067 );
   nor U10675 ( n11566,n11567,n11568,n11569,n11570 );
   buf U10676 ( p1_u3273,n19061 );
   nand U10677 ( n19061,n15916,n15917,n15918,n15919 );
   buf U10678 ( p1_u3249,n19086 );
   nand U10679 ( n19086,n16726,n16727,n16728,n16729 );
   buf U10680 ( p2_u3272,n19290 );
   nand U10681 ( n19290,n12191,n12192,n12193,n12194 );
   buf U10682 ( p1_u3271,n19063 );
   nand U10683 ( n19063,n15955,n15956,n15957,n15958 );
   buf U10684 ( p1_u3291,n19043 );
   nand U10685 ( n19043,n15349,n15350,n15351,n15352 );
   nor U10686 ( n15352,n15353,n15354,n15355 );
   nand U10687 ( n15350,p1_reg2_reg_0_,n15089 );
   buf U10688 ( p1_u3213,n19154 );
   nand U10689 ( n19154,n17883,n17884,n17885,n17886 );
   buf U10690 ( p2_u3240,n19351 );
   nand U10691 ( n19351,n13621,n13622,n13623,n13624 );
   buf U10692 ( p1_u3234,n19133 );
   nand U10693 ( n19133,n17567,n17568,n17569,n17570 );
   nand U10694 ( n17568,n17577,n17517 );
   buf U10695 ( p1_u3243,n19092 );
   nand U10696 ( n19092,n16892,n16854,n16893,n16894 );
   nor U10697 ( n16894,n16895,n16896,n16897 );
   buf U10698 ( p2_u3230,n19361 );
   nand U10699 ( n19361,n13767,n13768,n13769,n13770 );
   nand U10700 ( n13768,n13775,n13776,n13594 );
   buf U10701 ( p1_u3348,n18940 );
   nand U10702 ( n18940,n15153,n15154,n15155,n15156 );
   buf U10703 ( p1_u3346,n18942 );
   nand U10704 ( n18942,n15168,n15169,n15170,n15171 );
   buf U10705 ( p1_u3340,n18948 );
   nand U10706 ( n18948,n15204,n15205,n15206,n15207 );
   buf U10707 ( p1_u3338,n18950 );
   nand U10708 ( n18950,n15218,n15219,n15220,n15221 );
   buf U10709 ( p1_u3336,n18952 );
   nand U10710 ( n18952,n15233,n15234,n15235,n15236 );
   buf U10711 ( p1_u3335,n18953 );
   nand U10712 ( n18953,n15241,n15242,n15243,n15244 );
   buf U10713 ( p1_u3332,n18956 );
   nand U10714 ( n18956,n15262,n15263,n15264,n15265 );
   buf U10715 ( p1_u3330,n18958 );
   nand U10716 ( n18958,n15276,n15277,n15278,n15279 );
   buf U10717 ( p1_u3328,n18960 );
   nand U10718 ( n18960,n15290,n15291,n15292,n15293 );
   buf U10719 ( p1_u3326,n18962 );
   nand U10720 ( n18962,n15304,n15305,n15306,n15307 );
   buf U10721 ( p1_u3324,n18964 );
   nand U10722 ( n18964,n15318,n15319,n15320,n15321 );
   buf U10723 ( p1_u3323,n18965 );
   nand U10724 ( n18965,n15326,n15327,n15328,n15329 );
   buf U10725 ( p2_u3245,n19314 );
   nand U10726 ( n19314,n13053,n13054,n13055,n13056 );
   nand U10727 ( n13056,p2_ir_reg_0_,n13057 );
   buf U10728 ( p1_u3355,n19072 );
   nand U10729 ( n19072,n15075,n15076,n15077,n15078 );
   nor U10730 ( n15078,n15079,n15080,n15081 );
   buf U10731 ( p1_u3241,n19094 );
   nand U10732 ( n19094,n16942,n16943,n16944,n16945 );
   nand U10733 ( n16943,p1_addr_reg_0_,n16441 );
   buf U10734 ( p2_u3244,n19347 );
   nor U10735 ( n19347,n13076,n13077 );
   buf U10736 ( add_1071_u4,n18914 );
   xor U10737 ( n18914,n18846,n18847 );
   nor U10738 ( n10666,n10762,n10763,n10764 );
   not U10739 ( n10764,n11436 );
   buf U10740 ( p1_u4006,n19157 );
   not U10741 ( n14496,p1_u4006 );
   nor U10742 ( n19157,n16963,p1_u3084,n17488 );
   not U10743 ( n11472,n11457 );
   nor U10744 ( n11457,n11130,n11445,n10790 );
   nor U10745 ( n14766,n16426,n16274 );
   not U10746 ( n14803,n14698 );
   not U10747 ( n15378,n15086 );
   not U10748 ( n14729,n14717 );
   nor U10749 ( n14717,n17013,n17289 );
   not U10750 ( n15492,n16059 );
   nand U10751 ( n15495,n16443,n16979,n17286 );
   not U10752 ( n10668,n10666 );
   and U10753 ( n13548,n14438,n14440 );
   and U10754 ( n17397,n18696,n18695 );
   buf U10755 ( n10492,n15348 );
   nand U10756 ( n15069,n15061,n10492 );
   nor U10757 ( n18752,n18756,n10492 );
   nor U10758 ( n18767,n18772,n10492 );
   nor U10759 ( n18766,n18773,n10492 );
   nor U10760 ( n18758,n18761,n10492 );
   nor U10761 ( n18769,n18770,n10492 );
   nor U10762 ( n18768,n18771,n10492 );
   nor U10763 ( n18763,n10492,n15346 );
   nor U10764 ( n18765,n10492,n15347 );
   nor U10765 ( n18759,n10492,n15342 );
   nor U10766 ( n18760,n10492,n15345 );
   nor U10767 ( n18753,n10492,n15343 );
   nor U10768 ( n18754,n10492,n15341 );
   nor U10769 ( n18755,n10492,n15339 );
   nor U10770 ( n18757,n10492,n15340 );
   nor U10771 ( n18764,n10492,n15338 );
   nor U10772 ( n18762,n10492,n15344 );
   or U10773 ( n18745,n10492,p1_d_reg_1_ );
   or U10774 ( n18774,n10492,p1_d_reg_0_ );
   not U10775 ( n16461,n16855 );
   nor U10776 ( n11158,n11416,p2_state_reg );
   nand U10777 ( n11669,n13209,n11131 );
   not U10778 ( n17806,n18339 );
   nor U10779 ( n11154,n11414,p2_state_reg );
   nor U10780 ( n10803,n11126,n11127 );
   not U10781 ( n14693,n14701 );
   nand U10782 ( n14701,n14690,n15059 );
   not U10783 ( n14593,n14595 );
   nand U10784 ( n14595,n14689,n14690 );
   nor U10785 ( n15126,n11414,p1_state_reg );
   nor U10786 ( n15130,n11416,p1_state_reg );
   nor U10787 ( n17402,n11414,n16427 );
   nor U10788 ( n17407,n11416,n16427 );
   nor U10789 ( n15082,n16430,n15089 );
   not U10790 ( n10493,n17631 );
   not U10791 ( n17631,n17808 );
   xor U10792 ( n17801,n17807,n10493 );
   xor U10793 ( n17912,n17914,n17808 );
   xor U10794 ( n17949,n17948,n10493 );
   xor U10795 ( n18532,n18531,n17808 );
   xor U10796 ( n18684,n18683,n17808 );
   xor U10797 ( n17980,n17979,n17808 );
   xor U10798 ( n18041,n18040,n17808 );
   xor U10799 ( n18329,n18326,n10493 );
   nand U10800 ( n17808,n16980,n18687,n17288 );
   nand U10801 ( n14001,n11141,n14328,n14433 );
   not U10802 ( n15090,n15089 );
   nand U10803 ( n15089,n15061,n16432 );
   not U10804 ( n11445,n11455 );
   nand U10805 ( n11455,n12527,n12528 );
   not U10806 ( n13726,n13728 );
   nand U10807 ( n13728,n13214,n14425 );
   not U10808 ( n11414,n11416 );
   nand U10809 ( n11416,n18739,n18740 );
   not U10810 ( n17805,n18332 );
   nand U10811 ( n13265,n12349,n12366 );
   not U10812 ( n13297,n13361 );
   not U10813 ( u123,n10566 );
   buf U10814 ( p2_u3451,n19211 );
   nand U10815 ( n19211,n11118,n11119 );
   nand U10816 ( n11118,p2_reg0_reg_0_,n10775 );
   buf U10817 ( p2_u3454,n19212 );
   nand U10818 ( n19212,n11105,n11106 );
   nand U10819 ( n11105,p2_reg0_reg_1_,n10775 );
   buf U10820 ( p2_u3457,n19213 );
   nand U10821 ( n19213,n11093,n11094 );
   buf U10822 ( p2_u3460,n19214 );
   nand U10823 ( n19214,n11081,n11082 );
   buf U10824 ( p2_u3463,n19215 );
   nand U10825 ( n19215,n11069,n11070 );
   buf U10826 ( p2_u3466,n19216 );
   nand U10827 ( n19216,n11058,n11059 );
   buf U10828 ( p2_u3469,n19217 );
   nand U10829 ( n19217,n11046,n11047 );
   buf U10830 ( p2_u3472,n19218 );
   nand U10831 ( n19218,n11033,n11034 );
   buf U10832 ( p2_u3475,n19219 );
   nand U10833 ( n19219,n11022,n11023 );
   buf U10834 ( p2_u3478,n19220 );
   nand U10835 ( n19220,n11009,n11010 );
   buf U10836 ( p2_u3481,n19221 );
   nand U10837 ( n19221,n10998,n10999 );
   buf U10838 ( p2_u3484,n19222 );
   nand U10839 ( n19222,n10987,n10988 );
   buf U10840 ( p2_u3487,n19223 );
   nand U10841 ( n19223,n10976,n10977 );
   buf U10842 ( p2_u3490,n19224 );
   nand U10843 ( n19224,n10965,n10966 );
   buf U10844 ( p2_u3493,n19225 );
   nand U10845 ( n19225,n10954,n10955 );
   buf U10846 ( p2_u3496,n19226 );
   nand U10847 ( n19226,n10943,n10944 );
   buf U10848 ( p2_u3499,n19227 );
   nand U10849 ( n19227,n10932,n10933 );
   buf U10850 ( p2_u3502,n19228 );
   nand U10851 ( n19228,n10921,n10922 );
   buf U10852 ( p2_u3505,n19229 );
   nand U10853 ( n19229,n10910,n10911 );
   buf U10854 ( p2_u3507,n19230 );
   nand U10855 ( n19230,n10899,n10900 );
   buf U10856 ( p2_u3508,n19231 );
   nand U10857 ( n19231,n10888,n10889 );
   buf U10858 ( p2_u3509,n19232 );
   nand U10859 ( n19232,n10877,n10878 );
   buf U10860 ( p2_u3510,n19233 );
   nand U10861 ( n19233,n10866,n10867 );
   buf U10862 ( p2_u3511,n19234 );
   nand U10863 ( n19234,n10855,n10856 );
   buf U10864 ( p2_u3512,n19235 );
   nand U10865 ( n19235,n10842,n10843 );
   buf U10866 ( p2_u3513,n19236 );
   nand U10867 ( n19236,n10831,n10832 );
   buf U10868 ( p2_u3514,n19237 );
   nand U10869 ( n19237,n10820,n10821 );
   buf U10870 ( p2_u3515,n19238 );
   nand U10871 ( n19238,n10809,n10810 );
   buf U10872 ( p2_u3516,n19239 );
   nand U10873 ( n19239,n10795,n10796 );
   buf U10874 ( p2_u3517,n19240 );
   nand U10875 ( n19240,n10783,n10784 );
   buf U10876 ( p2_u3518,n19241 );
   nand U10877 ( n19241,n10776,n10777 );
   buf U10878 ( p2_u3519,n19242 );
   nand U10879 ( n19242,n10765,n10766 );
   buf U10880 ( p2_u3151,n19377 );
   nand U10881 ( n19377,n13074,n14472 );
   or U10882 ( n14472,n14318,n12522,n12521 );
   buf U10883 ( p1_u3240,n19127 );
   nand U10884 ( n19127,n16968,n16969 );
   buf U10885 ( p1_u3280,n19054 );
   nand U10886 ( n19054,n15690,n15691,n15692,n15693 );
   nor U10887 ( n15693,n15694,n15695,n15696,n15697 );
   buf U10888 ( p2_u3268,n19291 );
   nand U10889 ( n19291,n12307,n12308,n12309,n12310 );
   or U10890 ( n12309,n11460,n10807 );
   buf U10891 ( p1_u3269,n19065 );
   nand U10892 ( n19065,n16038,n16039,n16040,n16041 );
   buf U10893 ( p1_u3253,n19082 );
   nand U10894 ( n19082,n16625,n16626,n16627,n16628 );
   buf U10895 ( p1_u3250,n19085 );
   nand U10896 ( n19085,n16699,n16700,n16701,n16702 );
   buf U10897 ( p1_u3248,n19087 );
   nand U10898 ( n19087,n16752,n16753,n16754,n16755 );
   buf U10899 ( p1_u3247,n19088 );
   nand U10900 ( n19088,n16781,n16782,n16783,n16784 );
   buf U10901 ( p1_u3246,n19089 );
   nand U10902 ( n19089,n16811,n16812,n16813,n16814 );
   buf U10903 ( p2_u3257,n19302 );
   nand U10904 ( n19302,n12729,n12730,n12731,n12732 );
   buf U10905 ( p2_u3254,n19305 );
   nand U10906 ( n19305,n12813,n12814,n12815,n12816 );
   buf U10907 ( p2_u3252,n19307 );
   nand U10908 ( n19307,n12865,n12866,n12867,n12868 );
   buf U10909 ( p2_u3251,n19308 );
   nand U10910 ( n19308,n12894,n12895,n12896,n12897 );
   buf U10911 ( p2_u3250,n19309 );
   nand U10912 ( n19309,n12924,n12925,n12926,n12927 );
   buf U10913 ( p2_u3249,n19310 );
   nand U10914 ( n19310,n12953,n12954,n12955,n12956 );
   buf U10915 ( p1_u3242,n19093 );
   nand U10916 ( n19093,n16928,n16929,n16930,n16931 );
   buf U10917 ( p1_u3214,n19153 );
   nand U10918 ( n19153,n17870,n17871,n17872,n17873 );
   buf U10919 ( p2_u3218,n19373 );
   nand U10920 ( n19373,n13957,n13958,n13959,n13960 );
   buf U10921 ( p2_u3220,n19371 );
   nand U10922 ( n19371,n13928,n13929,n13930,n13931 );
   buf U10923 ( p1_u3230,n19137 );
   nand U10924 ( n19137,n17625,n17626,n17627,n17628 );
   buf U10925 ( add_1071_u55,n18915 );
   xor U10926 ( n18915,n18824,n18825 );
   buf U10927 ( add_1071_u56,n18916 );
   xor U10928 ( n18916,n18822,n18823 );
   buf U10929 ( add_1071_u57,n18917 );
   xor U10930 ( n18917,n18819,n18820 );
   buf U10931 ( add_1071_u58,n18918 );
   xor U10932 ( n18918,n18816,n18817 );
   buf U10933 ( add_1071_u59,n18919 );
   xor U10934 ( n18919,n18813,n18814 );
   buf U10935 ( add_1071_u60,n18920 );
   xor U10936 ( n18920,n18811,n18812 );
   buf U10937 ( add_1071_u61,n18921 );
   xor U10938 ( n18921,n18809,n18810 );
   buf U10939 ( add_1071_u62,n18922 );
   xor U10940 ( n18922,n18806,n18807 );
   buf U10941 ( add_1071_u63,n18923 );
   xor U10942 ( n18923,n18804,n18805 );
   buf U10943 ( add_1071_u47,n18924 );
   xor U10944 ( n18924,n18844,n18845 );
   buf U10945 ( add_1071_u48,n18925 );
   xor U10946 ( n18925,n18842,n18843 );
   buf U10947 ( add_1071_u49,n18926 );
   xor U10948 ( n18926,n18840,n18841 );
   buf U10949 ( add_1071_u50,n18927 );
   xor U10950 ( n18927,n18835,n18836 );
   buf U10951 ( add_1071_u51,n18928 );
   xor U10952 ( n18928,n18833,n18834 );
   buf U10953 ( add_1071_u52,n18929 );
   xor U10954 ( n18929,n18831,n18832 );
   buf U10955 ( add_1071_u53,n18930 );
   xor U10956 ( n18930,n18829,n18830 );
   buf U10957 ( add_1071_u54,n18931 );
   xor U10958 ( n18931,n18827,n18828 );
   buf U10959 ( add_1071_u5,n18932 );
   xor U10960 ( n18932,n18837,n18838 );
   xor U10961 ( n18838,n18839,n16934 );
   not U10962 ( n10775,n10767 );
   nor U10963 ( n10767,n10762,n11133,n10764 );
   nor U10964 ( n15128,p1_u3084,p1_ir_reg_31_ );
   nor U10965 ( n15129,n15128,p1_u3084 );
   not U10966 ( p1_u3084,p1_state_reg );
   nor U10967 ( n11156,p2_u3152,p2_ir_reg_31_ );
   not U10968 ( p2_u3152,p2_state_reg );
   xor U10969 ( n10566,p2_wr_reg,p1_wr_reg );
   nand U10970 ( n10567,n19378,n10570 );
   nand U10971 ( n10571,n19378,n10573 );
   nand U10972 ( n10574,n19378,n10576 );
   nand U10973 ( n10577,n19378,n10579 );
   nand U10974 ( n10580,n19378,n10582 );
   nand U10975 ( n10583,n19378,n10585 );
   nand U10976 ( n10586,n19378,n10588 );
   nand U10977 ( n10589,n19378,n10591 );
   nand U10978 ( n10592,n19378,n10594 );
   nand U10979 ( n10595,n19378,n10597 );
   nand U10980 ( n10598,n19378,n10600 );
   nand U10981 ( n10601,n19378,n10603 );
   nand U10982 ( n10604,n19378,n10606 );
   nand U10983 ( n10607,n19378,n10609 );
   nand U10984 ( n10610,n19378,n10612 );
   nand U10985 ( n10613,n19378,n10615 );
   nand U10986 ( n10616,n19378,n10618 );
   nand U10987 ( n10619,n19378,n10621 );
   nand U10988 ( n10622,n19378,n10624 );
   nand U10989 ( n10625,n19378,n10627 );
   nand U10990 ( n10628,n19378,n10630 );
   nand U10991 ( n10631,n19378,n10633 );
   nand U10992 ( n10634,n19378,n10636 );
   nand U10993 ( n10637,n19378,n10639 );
   nand U10994 ( n10640,n19378,n10642 );
   nand U10995 ( n10643,n19378,n10645 );
   nand U10996 ( n10646,n19378,n10648 );
   nand U10997 ( n10649,n19378,n10651 );
   nand U10998 ( n10652,n19378,n10654 );
   nand U10999 ( n10655,n19378,n10657 );
   nand U11000 ( n10658,n19378,n10660 );
   nand U11001 ( n10661,n19378,n10663 );
   nand U11002 ( n10665,n10666,n10667 );
   nand U11003 ( n10664,p2_reg1_reg_31_,n10668 );
   nand U11004 ( n10670,p2_reg1_reg_30_,n10668 );
   nand U11005 ( n10669,n10666,n10671 );
   nand U11006 ( n10673,p2_reg1_reg_29_,n10668 );
   nand U11007 ( n10672,n10666,n10674 );
   nand U11008 ( n10676,p2_reg1_reg_28_,n10668 );
   nand U11009 ( n10675,n10666,n10677 );
   nand U11010 ( n10679,p2_reg1_reg_27_,n10668 );
   nand U11011 ( n10678,n10666,n10680 );
   nand U11012 ( n10682,p2_reg1_reg_26_,n10668 );
   nand U11013 ( n10681,n10666,n10683 );
   nand U11014 ( n10685,p2_reg1_reg_25_,n10668 );
   nand U11015 ( n10684,n10666,n10686 );
   nand U11016 ( n10688,p2_reg1_reg_24_,n10668 );
   nand U11017 ( n10687,n10666,n10689 );
   nand U11018 ( n10691,p2_reg1_reg_23_,n10668 );
   nand U11019 ( n10690,n10666,n10692 );
   nand U11020 ( n10694,p2_reg1_reg_22_,n10668 );
   nand U11021 ( n10693,n10666,n10695 );
   nand U11022 ( n10697,p2_reg1_reg_21_,n10668 );
   nand U11023 ( n10696,n10666,n10698 );
   nand U11024 ( n10700,p2_reg1_reg_20_,n10668 );
   nand U11025 ( n10699,n10666,n10701 );
   nand U11026 ( n10703,p2_reg1_reg_19_,n10668 );
   nand U11027 ( n10702,n10666,n10704 );
   nand U11028 ( n10706,p2_reg1_reg_18_,n10668 );
   nand U11029 ( n10705,n10666,n10707 );
   nand U11030 ( n10709,p2_reg1_reg_17_,n10668 );
   nand U11031 ( n10708,n10666,n10710 );
   nand U11032 ( n10712,p2_reg1_reg_16_,n10668 );
   nand U11033 ( n10711,n10666,n10713 );
   nand U11034 ( n10715,p2_reg1_reg_15_,n10668 );
   nand U11035 ( n10714,n10666,n10716 );
   nand U11036 ( n10718,p2_reg1_reg_14_,n10668 );
   nand U11037 ( n10717,n10666,n10719 );
   nand U11038 ( n10721,p2_reg1_reg_13_,n10668 );
   nand U11039 ( n10720,n10666,n10722 );
   nand U11040 ( n10724,p2_reg1_reg_12_,n10668 );
   nand U11041 ( n10723,n10666,n10725 );
   nand U11042 ( n10727,p2_reg1_reg_11_,n10668 );
   nand U11043 ( n10726,n10666,n10728 );
   nand U11044 ( n10730,p2_reg1_reg_10_,n10668 );
   nand U11045 ( n10729,n10666,n10731 );
   nand U11046 ( n10733,p2_reg1_reg_9_,n10668 );
   nand U11047 ( n10732,n10666,n10734 );
   nand U11048 ( n10736,p2_reg1_reg_8_,n10668 );
   nand U11049 ( n10735,n10666,n10737 );
   nand U11050 ( n10739,p2_reg1_reg_7_,n10668 );
   nand U11051 ( n10738,n10666,n10740 );
   nand U11052 ( n10742,p2_reg1_reg_6_,n10668 );
   nand U11053 ( n10741,n10666,n10743 );
   nand U11054 ( n10745,p2_reg1_reg_5_,n10668 );
   nand U11055 ( n10744,n10666,n10746 );
   nand U11056 ( n10748,p2_reg1_reg_4_,n10668 );
   nand U11057 ( n10747,n10666,n10749 );
   nand U11058 ( n10750,n10666,n10752 );
   nand U11059 ( n10753,n10666,n10755 );
   nand U11060 ( n10756,n10666,n10758 );
   nand U11061 ( n10759,n10666,n10761 );
   nand U11062 ( n10766,n10767,n10667 );
   nand U11063 ( n10667,n10768,n10769,n10770 );
   nand U11064 ( n10770,n10771,n10772 );
   nand U11065 ( n10768,n10773,n10774 );
   nand U11066 ( n10765,p2_reg0_reg_31_,n10775 );
   nand U11067 ( n10777,n10767,n10671 );
   nand U11068 ( n10671,n10778,n10769,n10779 );
   nand U11069 ( n10779,n10780,n10772 );
   nand U11070 ( n10778,n10781,n10782,n10773 );
   nand U11071 ( n10776,p2_reg0_reg_30_,n10775 );
   nand U11072 ( n10784,n10767,n10674 );
   nand U11073 ( n10674,n10785,n10786,n10787,n10788 );
   or U11074 ( n10788,n10789,n10790 );
   nand U11075 ( n10787,n10791,n10772 );
   or U11076 ( n10786,n10792,n10793 );
   not U11077 ( n10785,n10794 );
   nand U11078 ( n10783,p2_reg0_reg_29_,n10775 );
   nand U11079 ( n10796,n10767,n10677 );
   nand U11080 ( n10677,n10797,n10798,n10799 );
   nor U11081 ( n10799,n10800,n10801,n10802 );
   nor U11082 ( n10802,n10803,n10804 );
   and U11083 ( n10801,n10805,n10806 );
   nor U11084 ( n10800,n10790,n10807 );
   nand U11085 ( n10798,n10808,n10576 );
   nand U11086 ( n10795,p2_reg0_reg_28_,n10775 );
   nand U11087 ( n10810,n10767,n10680 );
   nand U11088 ( n10680,n10811,n10812,n10813 );
   nor U11089 ( n10813,n10814,n10815,n10816 );
   nor U11090 ( n10816,n10803,n10817 );
   nor U11091 ( n10815,n10790,n10818 );
   nor U11092 ( n10814,n10792,n10819 );
   nand U11093 ( n10812,n10808,n10579 );
   nand U11094 ( n10809,p2_reg0_reg_27_,n10775 );
   nand U11095 ( n10821,n10767,n10683 );
   nand U11096 ( n10683,n10822,n10823,n10824 );
   nor U11097 ( n10824,n10825,n10826,n10827 );
   nor U11098 ( n10827,n10792,n10828 );
   nor U11099 ( n10826,n10803,n10829 );
   nor U11100 ( n10825,n10790,n10830 );
   nand U11101 ( n10823,n10808,n10582 );
   nand U11102 ( n10820,p2_reg0_reg_26_,n10775 );
   nand U11103 ( n10832,n10767,n10686 );
   nand U11104 ( n10686,n10833,n10834,n10835 );
   nor U11105 ( n10835,n10836,n10837,n10838 );
   nor U11106 ( n10838,n10790,n10839 );
   nor U11107 ( n10837,n10840,n10792 );
   nor U11108 ( n10836,n10803,n10841 );
   nand U11109 ( n10834,n10808,n10585 );
   nand U11110 ( n10831,p2_reg0_reg_25_,n10775 );
   nand U11111 ( n10843,n10767,n10689 );
   nand U11112 ( n10689,n10844,n10845,n10846,n10847 );
   nor U11113 ( n10847,n10848,n10849 );
   nor U11114 ( n10848,n10850,n10851 );
   nand U11115 ( n10846,n10852,n10773 );
   nand U11116 ( n10845,n10853,n10772 );
   nand U11117 ( n10844,n10805,n10854 );
   nand U11118 ( n10842,p2_reg0_reg_24_,n10775 );
   nand U11119 ( n10856,n10767,n10692 );
   nand U11120 ( n10692,n10857,n10858,n10859 );
   nor U11121 ( n10859,n10860,n10861,n10862 );
   nor U11122 ( n10862,n10803,n10863 );
   nor U11123 ( n10861,n10790,n10864 );
   nor U11124 ( n10860,n10865,n10792 );
   nand U11125 ( n10858,n10808,n10591 );
   nand U11126 ( n10855,p2_reg0_reg_23_,n10775 );
   nand U11127 ( n10867,n10767,n10695 );
   nand U11128 ( n10695,n10868,n10869,n10870 );
   nor U11129 ( n10870,n10871,n10872,n10873 );
   nor U11130 ( n10873,n10792,n10874 );
   nor U11131 ( n10872,n10803,n10875 );
   nor U11132 ( n10871,n10790,n10876 );
   nand U11133 ( n10869,n10808,n10594 );
   nand U11134 ( n10866,p2_reg0_reg_22_,n10775 );
   nand U11135 ( n10878,n10767,n10698 );
   nand U11136 ( n10698,n10879,n10880,n10881 );
   nor U11137 ( n10881,n10882,n10883,n10884 );
   nor U11138 ( n10884,n10803,n10885 );
   nor U11139 ( n10883,n10790,n10886 );
   nor U11140 ( n10882,n10792,n10887 );
   nand U11141 ( n10880,n10808,n10597 );
   nand U11142 ( n10877,p2_reg0_reg_21_,n10775 );
   nand U11143 ( n10889,n10767,n10701 );
   nand U11144 ( n10701,n10890,n10891,n10892 );
   nor U11145 ( n10892,n10893,n10894,n10895 );
   nor U11146 ( n10895,n10792,n10896 );
   nor U11147 ( n10894,n10803,n10897 );
   nor U11148 ( n10893,n10790,n10898 );
   nand U11149 ( n10891,n10808,n10600 );
   nand U11150 ( n10888,p2_reg0_reg_20_,n10775 );
   nand U11151 ( n10900,n10767,n10704 );
   nand U11152 ( n10704,n10901,n10902,n10903 );
   nor U11153 ( n10903,n10904,n10905,n10906 );
   nor U11154 ( n10906,n10803,n10907 );
   nor U11155 ( n10905,n10790,n10908 );
   nor U11156 ( n10904,n10792,n10909 );
   nand U11157 ( n10902,n10808,n10603 );
   nand U11158 ( n10899,p2_reg0_reg_19_,n10775 );
   nand U11159 ( n10911,n10767,n10707 );
   nand U11160 ( n10707,n10912,n10913,n10914 );
   nor U11161 ( n10914,n10915,n10916,n10917 );
   nor U11162 ( n10917,n10803,n10918 );
   nor U11163 ( n10916,n10792,n10919 );
   nor U11164 ( n10915,n10790,n10920 );
   nand U11165 ( n10913,n10808,n10606 );
   nand U11166 ( n10910,p2_reg0_reg_18_,n10775 );
   nand U11167 ( n10922,n10767,n10710 );
   nand U11168 ( n10710,n10923,n10924,n10925 );
   nor U11169 ( n10925,n10926,n10927,n10928 );
   nor U11170 ( n10928,n10803,n10929 );
   nor U11171 ( n10927,n10790,n10930 );
   nor U11172 ( n10926,n10792,n10931 );
   nand U11173 ( n10924,n10808,n10609 );
   nand U11174 ( n10921,p2_reg0_reg_17_,n10775 );
   nand U11175 ( n10933,n10767,n10713 );
   nand U11176 ( n10713,n10934,n10935,n10936,n10937 );
   nand U11177 ( n10937,n10938,n10773 );
   nor U11178 ( n10936,n10939,n10940 );
   nor U11179 ( n10940,n10803,n10941 );
   nor U11180 ( n10939,n10942,n10792 );
   nand U11181 ( n10935,n10808,n10612 );
   nand U11182 ( n10932,p2_reg0_reg_16_,n10775 );
   nand U11183 ( n10944,n10767,n10716 );
   nand U11184 ( n10716,n10945,n10946,n10947 );
   nor U11185 ( n10947,n10948,n10949,n10950 );
   nor U11186 ( n10950,n10803,n10951 );
   nor U11187 ( n10949,n10790,n10952 );
   nor U11188 ( n10948,n10792,n10953 );
   nand U11189 ( n10946,n10808,n10615 );
   nand U11190 ( n10943,p2_reg0_reg_15_,n10775 );
   nand U11191 ( n10955,n10767,n10719 );
   nand U11192 ( n10719,n10956,n10957,n10958 );
   nor U11193 ( n10958,n10959,n10960,n10961 );
   nor U11194 ( n10961,n10792,n10962 );
   nor U11195 ( n10960,n10803,n10963 );
   nor U11196 ( n10959,n10790,n10964 );
   nand U11197 ( n10957,n10808,n10618 );
   nand U11198 ( n10954,p2_reg0_reg_14_,n10775 );
   nand U11199 ( n10966,n10767,n10722 );
   nand U11200 ( n10722,n10967,n10968,n10969 );
   nor U11201 ( n10969,n10970,n10971,n10972 );
   nor U11202 ( n10972,n10803,n10973 );
   and U11203 ( n10971,n10974,n10773 );
   nor U11204 ( n10970,n10792,n10975 );
   nand U11205 ( n10968,n10808,n10621 );
   nand U11206 ( n10965,p2_reg0_reg_13_,n10775 );
   nand U11207 ( n10977,n10767,n10725 );
   nand U11208 ( n10725,n10978,n10979,n10980 );
   nor U11209 ( n10980,n10981,n10982,n10983 );
   nor U11210 ( n10983,n10792,n10984 );
   nor U11211 ( n10982,n10803,n10985 );
   nor U11212 ( n10981,n10790,n10986 );
   nand U11213 ( n10979,n10808,n10624 );
   nand U11214 ( n10976,p2_reg0_reg_12_,n10775 );
   nand U11215 ( n10988,n10767,n10728 );
   nand U11216 ( n10728,n10989,n10990,n10991 );
   nor U11217 ( n10991,n10992,n10993,n10994 );
   nor U11218 ( n10994,n10803,n10995 );
   nor U11219 ( n10993,n10790,n10996 );
   nor U11220 ( n10992,n10792,n10997 );
   nand U11221 ( n10990,n10808,n10627 );
   nand U11222 ( n10987,p2_reg0_reg_11_,n10775 );
   nand U11223 ( n10999,n10767,n10731 );
   nand U11224 ( n10731,n11000,n11001,n11002 );
   nor U11225 ( n11002,n11003,n11004,n11005 );
   nor U11226 ( n11005,n10792,n11006 );
   nor U11227 ( n11004,n10803,n11007 );
   nor U11228 ( n11003,n10790,n11008 );
   nand U11229 ( n11001,n10808,n10630 );
   nand U11230 ( n10998,p2_reg0_reg_10_,n10775 );
   nand U11231 ( n11010,n10767,n10734 );
   nand U11232 ( n10734,n11011,n11012,n11013,n11014 );
   nor U11233 ( n11014,n11015,n11016 );
   nor U11234 ( n11015,n11017,n10851 );
   nand U11235 ( n11013,n11018,n10772 );
   nand U11236 ( n11012,n11019,n10773 );
   nand U11237 ( n11011,n11020,n11021 );
   nand U11238 ( n11009,p2_reg0_reg_9_,n10775 );
   nand U11239 ( n11023,n10767,n10737 );
   nand U11240 ( n10737,n11024,n11025,n11026 );
   nor U11241 ( n11026,n11027,n11028,n11029 );
   nor U11242 ( n11029,n10792,n11030 );
   nor U11243 ( n11028,n10803,n11031 );
   nor U11244 ( n11027,n10790,n11032 );
   nand U11245 ( n11025,n10808,n10636 );
   nand U11246 ( n11022,p2_reg0_reg_8_,n10775 );
   nand U11247 ( n11034,n10767,n10740 );
   nand U11248 ( n10740,n11035,n11036,n11037,n11038 );
   nor U11249 ( n11038,n11039,n11040 );
   nor U11250 ( n11039,n11041,n10851 );
   nand U11251 ( n11037,n11042,n10772 );
   nand U11252 ( n11036,n11043,n11021,n11044 );
   nand U11253 ( n11035,n11045,n10773 );
   nand U11254 ( n11033,p2_reg0_reg_7_,n10775 );
   nand U11255 ( n11047,n10767,n10743 );
   nand U11256 ( n10743,n11048,n11049,n11050,n11051 );
   nor U11257 ( n11051,n11052,n11053 );
   nor U11258 ( n11052,n11054,n10851 );
   nand U11259 ( n11050,n11055,n10773 );
   nand U11260 ( n11049,n11056,n11021 );
   nand U11261 ( n11048,n11057,n10772 );
   nand U11262 ( n11046,p2_reg0_reg_6_,n10775 );
   nand U11263 ( n11059,n10767,n10746 );
   nand U11264 ( n10746,n11060,n11061,n11062 );
   nor U11265 ( n11062,n11063,n11064,n11065 );
   and U11266 ( n11065,n11021,n11066 );
   nor U11267 ( n11064,n10790,n11067 );
   nor U11268 ( n11063,n10803,n11068 );
   nand U11269 ( n11061,n10808,n10645 );
   nand U11270 ( n11058,p2_reg0_reg_5_,n10775 );
   nand U11271 ( n11070,n10767,n10749 );
   nand U11272 ( n10749,n11071,n11072,n11073,n11074 );
   nor U11273 ( n11074,n11075,n11076 );
   nor U11274 ( n11075,n11077,n10851 );
   nand U11275 ( n11073,n11078,n10773 );
   nand U11276 ( n11072,n11079,n11021 );
   nand U11277 ( n11071,n11080,n10772 );
   nand U11278 ( n11069,p2_reg0_reg_4_,n10775 );
   nand U11279 ( n11082,n10767,n10752 );
   nand U11280 ( n10752,n11083,n11084,n11085,n11086 );
   nor U11281 ( n11086,n11087,n11088 );
   nor U11282 ( n11087,n11089,n10851 );
   nand U11283 ( n11085,n11090,n10772 );
   nand U11284 ( n11084,n10773,n11091 );
   nand U11285 ( n11083,n11092,n11021 );
   nand U11286 ( n11081,p2_reg0_reg_3_,n10775 );
   nand U11287 ( n11094,n10767,n10755 );
   nand U11288 ( n10755,n11095,n11096,n11097,n11098 );
   nor U11289 ( n11098,n11099,n11100 );
   nor U11290 ( n11099,n11101,n10851 );
   nand U11291 ( n11097,n11102,n10773 );
   nand U11292 ( n11096,n11103,n11021 );
   nand U11293 ( n11095,n11104,n10772 );
   nand U11294 ( n11093,p2_reg0_reg_2_,n10775 );
   nand U11295 ( n11106,n10767,n10758 );
   nand U11296 ( n10758,n11107,n11108,n11109,n11110 );
   nor U11297 ( n11110,n11111,n11112 );
   nor U11298 ( n11111,n11113,n10851 );
   nand U11299 ( n11109,n11114,n10772 );
   not U11300 ( n10772,n10803 );
   nand U11301 ( n11108,n10773,n11115 );
   nand U11302 ( n11107,n11116,n11021 );
   or U11303 ( n11021,n11117,n10805 );
   nand U11304 ( n11119,n10767,n10761 );
   nand U11305 ( n10761,n11120,n11121,n11122,n11123 );
   nand U11306 ( n11123,n11124,n11125 );
   nand U11307 ( n11124,n10803,n10790 );
   not U11308 ( n11126,n11128 );
   nand U11309 ( n11122,n11129,n10805 );
   nor U11310 ( n10805,n11130,n11131,n11132 );
   nand U11311 ( n11121,n10808,n10660 );
   not U11312 ( n11133,n10763 );
   nand U11313 ( n10762,n11134,n11135,n11136 );
   nand U11314 ( n11136,n11137,n11138,n11139,n11140 );
   nand U11315 ( n11140,n11131,n11141 );
   nand U11316 ( n11139,n11132,n11142 );
   nand U11317 ( n11144,p2_d_reg_1_,n11145 );
   nand U11318 ( n11143,n11146,n11147 );
   nand U11319 ( n11149,p2_d_reg_0_,n11145 );
   nand U11320 ( n11148,n11146,n11150 );
   nand U11321 ( n11153,n11154,p1_datao_reg_0_ );
   nand U11322 ( n11152,p2_ir_reg_0_,n11155 );
   or U11323 ( n11155,n11156,n11157 );
   nand U11324 ( n11151,n11158,n11159 );
   nand U11325 ( n11163,n11157,n11164 );
   nand U11326 ( n11162,n11158,n11165 );
   nand U11327 ( n11161,n11154,p1_datao_reg_1_ );
   nand U11328 ( n11160,n11156,p2_ir_reg_1_ );
   nand U11329 ( n11169,n11170,n11157 );
   not U11330 ( n11170,n11171 );
   nand U11331 ( n11168,n11158,n11172 );
   nand U11332 ( n11167,n11154,p1_datao_reg_2_ );
   nand U11333 ( n11166,n11156,p2_ir_reg_2_ );
   nand U11334 ( n11176,n11177,n11157 );
   nand U11335 ( n11175,n11158,n11178 );
   nand U11336 ( n11174,n11154,p1_datao_reg_3_ );
   nand U11337 ( n11173,n11156,p2_ir_reg_3_ );
   nand U11338 ( n11182,n11183,n11184,n11157 );
   nand U11339 ( n11181,n11185,n11158 );
   nand U11340 ( n11180,n11154,p1_datao_reg_4_ );
   nand U11341 ( n11179,n11156,p2_ir_reg_4_ );
   nand U11342 ( n11189,p2_ir_reg_5_,n11190 );
   nand U11343 ( n11190,n11191,n11192 );
   nand U11344 ( n11192,n11157,n11193 );
   nand U11345 ( n11188,n11157,n11184,n11194 );
   nand U11346 ( n11187,n11195,n11158 );
   nand U11347 ( n11186,n11154,p1_datao_reg_5_ );
   nand U11348 ( n11199,n11200,n11201,n11157 );
   nand U11349 ( n11198,n11158,n11202 );
   nand U11350 ( n11197,n11154,p1_datao_reg_6_ );
   nand U11351 ( n11196,n11156,p2_ir_reg_6_ );
   nand U11352 ( n11206,p2_ir_reg_7_,n11207 );
   nand U11353 ( n11207,n11191,n11208 );
   nand U11354 ( n11208,n11157,n11209 );
   nand U11355 ( n11205,n11157,n11201,n11210 );
   nand U11356 ( n11204,n11211,n11158 );
   nand U11357 ( n11203,n11154,p1_datao_reg_7_ );
   nand U11358 ( n11215,n11216,n11217,n11157 );
   nand U11359 ( n11214,n11218,n11158 );
   nand U11360 ( n11213,n11154,p1_datao_reg_8_ );
   nand U11361 ( n11212,n11156,p2_ir_reg_8_ );
   nand U11362 ( n11222,p2_ir_reg_9_,n11223 );
   nand U11363 ( n11223,n11191,n11224 );
   nand U11364 ( n11224,n11157,n11225 );
   nand U11365 ( n11221,n11157,n11217,n11226 );
   nand U11366 ( n11220,n11227,n11158 );
   nand U11367 ( n11219,n11154,p1_datao_reg_9_ );
   nand U11368 ( n11231,n11232,n11157 );
   not U11369 ( n11232,n11233 );
   nand U11370 ( n11230,n11158,n11234 );
   nand U11371 ( n11229,n11154,p1_datao_reg_10_ );
   nand U11372 ( n11228,n11156,p2_ir_reg_10_ );
   nand U11373 ( n11238,p2_ir_reg_11_,n11239 );
   nand U11374 ( n11239,n11191,n11240 );
   nand U11375 ( n11240,n11157,n11241 );
   nand U11376 ( n11237,n11157,n11242,n11243 );
   nand U11377 ( n11236,n11244,n11158 );
   nand U11378 ( n11235,n11154,p1_datao_reg_11_ );
   nand U11379 ( n11248,n11249,n11157 );
   not U11380 ( n11249,n11250 );
   nand U11381 ( n11247,n11251,n11158 );
   nand U11382 ( n11246,n11154,p1_datao_reg_12_ );
   nand U11383 ( n11245,n11156,p2_ir_reg_12_ );
   nand U11384 ( n11255,p2_ir_reg_13_,n11256 );
   nand U11385 ( n11256,n11191,n11257 );
   nand U11386 ( n11257,n11157,n11258 );
   nand U11387 ( n11254,n11157,n11259,n11260 );
   nand U11388 ( n11253,n11158,n11261 );
   nand U11389 ( n11252,n11154,p1_datao_reg_13_ );
   nand U11390 ( n11265,n11266,n11157 );
   not U11391 ( n11266,n11267 );
   nand U11392 ( n11264,n11158,n11268 );
   nand U11393 ( n11263,n11154,p1_datao_reg_14_ );
   nand U11394 ( n11262,n11156,p2_ir_reg_14_ );
   nand U11395 ( n11272,p2_ir_reg_15_,n11273 );
   nand U11396 ( n11273,n11191,n11274 );
   nand U11397 ( n11274,n11157,n11275 );
   nand U11398 ( n11271,n11157,n11276,n11277 );
   nand U11399 ( n11270,n11278,n11158 );
   nand U11400 ( n11269,n11154,p1_datao_reg_15_ );
   nand U11401 ( n11282,n11283,n11157 );
   not U11402 ( n11283,n11284 );
   nand U11403 ( n11281,n11285,n11158 );
   nand U11404 ( n11280,p1_datao_reg_16_,n11154 );
   nand U11405 ( n11279,n11156,p2_ir_reg_16_ );
   nand U11406 ( n11289,p2_ir_reg_17_,n11290 );
   nand U11407 ( n11290,n11191,n11291 );
   nand U11408 ( n11291,n11157,n11292 );
   nand U11409 ( n11288,n11157,n11293,n11294 );
   nand U11410 ( n11287,n11295,n11158 );
   nand U11411 ( n11286,p1_datao_reg_17_,n11154 );
   nand U11412 ( n11299,p2_ir_reg_18_,n11300 );
   nand U11413 ( n11300,n11191,n11301 );
   nand U11414 ( n11301,n11157,n11302 );
   nand U11415 ( n11298,n11157,n11303,n11304 );
   nand U11416 ( n11297,n11305,n11158 );
   nand U11417 ( n11296,p1_datao_reg_18_,n11154 );
   nand U11418 ( n11309,n11310,n11311,n11157 );
   nand U11419 ( n11308,n11312,n11158 );
   nand U11420 ( n11307,p1_datao_reg_19_,n11154 );
   nand U11421 ( n11306,n11156,p2_ir_reg_19_ );
   nand U11422 ( n11316,n11317,n11318,n11157 );
   nand U11423 ( n11315,n11319,n11158 );
   nand U11424 ( n11314,p1_datao_reg_20_,n11154 );
   nand U11425 ( n11313,n11156,p2_ir_reg_20_ );
   nand U11426 ( n11323,p2_ir_reg_21_,n11324 );
   nand U11427 ( n11324,n11191,n11325 );
   nand U11428 ( n11325,n11157,n11326 );
   nand U11429 ( n11322,n11157,n11318,n11327 );
   nand U11430 ( n11321,n11328,n11158 );
   nand U11431 ( n11320,p1_datao_reg_21_,n11154 );
   nand U11432 ( n11332,p2_ir_reg_22_,n11333 );
   nand U11433 ( n11333,n11191,n11334 );
   nand U11434 ( n11334,n11157,n11335 );
   nand U11435 ( n11331,n11157,n11336,n11337 );
   nand U11436 ( n11330,n11338,n11158 );
   nand U11437 ( n11329,p1_datao_reg_22_,n11154 );
   nand U11438 ( n11342,n11343,n11344,n11157 );
   nand U11439 ( n11341,n11345,n11158 );
   nand U11440 ( n11340,p1_datao_reg_23_,n11154 );
   nand U11441 ( n11339,n11156,p2_ir_reg_23_ );
   nand U11442 ( n11349,p2_ir_reg_24_,n11350 );
   nand U11443 ( n11350,n11191,n11351 );
   nand U11444 ( n11351,n11352,n11157 );
   nand U11445 ( n11348,n11157,n11343,n11353 );
   nand U11446 ( n11347,n11354,n11158 );
   nand U11447 ( n11346,p1_datao_reg_24_,n11154 );
   nand U11448 ( n11358,p2_ir_reg_25_,n11359 );
   nand U11449 ( n11359,n11191,n11360 );
   nand U11450 ( n11360,n11157,n11361 );
   nand U11451 ( n11357,n11157,n11362,n11363 );
   nand U11452 ( n11356,n11364,n11158 );
   nand U11453 ( n11355,p1_datao_reg_25_,n11154 );
   nand U11454 ( n11368,n11369,n11370,n11157 );
   nand U11455 ( n11367,n11371,n11158 );
   nand U11456 ( n11366,p1_datao_reg_26_,n11154 );
   nand U11457 ( n11365,n11156,p2_ir_reg_26_ );
   nand U11458 ( n11375,p2_ir_reg_27_,n11376 );
   nand U11459 ( n11376,n11191,n11377 );
   nand U11460 ( n11377,n11157,n11378 );
   nand U11461 ( n11374,n11157,n11369,n11379 );
   nand U11462 ( n11373,n11380,n11158 );
   nand U11463 ( n11372,p1_datao_reg_27_,n11154 );
   nand U11464 ( n11384,p2_ir_reg_28_,n11385 );
   nand U11465 ( n11385,n11191,n11386 );
   nand U11466 ( n11386,n11157,n11387 );
   nand U11467 ( n11383,n11157,n11388,n11389 );
   nand U11468 ( n11382,n11390,n11158 );
   nand U11469 ( n11381,p1_datao_reg_28_,n11154 );
   nand U11470 ( n11394,p2_ir_reg_29_,n11395 );
   nand U11471 ( n11395,n11191,n11396 );
   nand U11472 ( n11396,n11397,n11157 );
   nand U11473 ( n11393,n11157,n11398,n11399 );
   not U11474 ( n11399,p2_ir_reg_29_ );
   nand U11475 ( n11392,n11158,n11400 );
   nand U11476 ( n11391,n11154,p1_datao_reg_29_ );
   nand U11477 ( n11404,p2_ir_reg_30_,n11405 );
   nand U11478 ( n11405,n11191,n11406 );
   nand U11479 ( n11406,n11407,n11157 );
   not U11480 ( n11191,n11156 );
   nand U11481 ( n11403,n11157,n11408,n11409 );
   not U11482 ( n11408,n11407 );
   nand U11483 ( n11402,n11410,n11158 );
   nand U11484 ( n11401,n11154,p1_datao_reg_30_ );
   nand U11485 ( n11413,n11154,p1_datao_reg_31_ );
   nand U11486 ( n11412,n11157,n11409,n11407 );
   nor U11487 ( n11407,n11398,p2_ir_reg_29_ );
   not U11488 ( n11409,p2_ir_reg_30_ );
   nor U11489 ( n11441,n11442,n11443,n11444 );
   nor U11490 ( n11444,n11120,n11445 );
   and U11491 ( n11120,n11446,n11447 );
   nand U11492 ( n11447,n11448,n11449 );
   nand U11493 ( n11448,n11450,n11451 );
   nand U11494 ( n11451,n11452,n10663 );
   nand U11495 ( n11446,n11129,n11117 );
   not U11496 ( n11129,n11453 );
   nor U11497 ( n11443,n11454,n11455 );
   nor U11498 ( n11442,n11453,n11456 );
   nand U11499 ( n11440,n11457,p2_reg3_reg_0_ );
   nand U11500 ( n11458,n11459,n11460 );
   nand U11501 ( n11438,n11461,n10660 );
   nor U11502 ( n11469,n11470,n11459 );
   nor U11503 ( n11468,n11471,n11472 );
   and U11504 ( n11467,n11112,n11455 );
   nand U11505 ( n11112,n11473,n11474 );
   nand U11506 ( n11474,n11475,n11449 );
   xor U11507 ( n11475,n11476,n11450 );
   nand U11508 ( n11473,n11477,n10663 );
   nor U11509 ( n11466,n11478,n11455 );
   nand U11510 ( n11464,n11461,n10657 );
   nand U11511 ( n11463,n11479,n11115 );
   xor U11512 ( n11115,n11114,n11125 );
   nand U11513 ( n11462,n11116,n11480 );
   xor U11514 ( n11116,n11481,n11476 );
   nor U11515 ( n11489,n11490,n11459 );
   nor U11516 ( n11488,n11491,n11472 );
   and U11517 ( n11487,n11100,n11455 );
   nand U11518 ( n11100,n11492,n11493 );
   nand U11519 ( n11493,n11494,n11495,n11496 );
   or U11520 ( n11495,n11497,n11498 );
   nand U11521 ( n11494,n11499,n11500 );
   not U11522 ( n11499,n11501 );
   nand U11523 ( n11492,n11477,n10660 );
   nor U11524 ( n11486,n11502,n11455 );
   nand U11525 ( n11484,n11461,n10654 );
   nand U11526 ( n11483,n11103,n11480 );
   and U11527 ( n11103,n11503,n11504 );
   or U11528 ( n11504,n11497,n11505 );
   nand U11529 ( n11503,n11506,n11500,n11505 );
   nor U11530 ( n11505,n11507,n11508 );
   nand U11531 ( n11482,n11479,n11102 );
   and U11532 ( n11102,n11509,n11510 );
   nand U11533 ( n11510,n11104,n11511 );
   nand U11534 ( n11511,n11470,n11452 );
   not U11535 ( n11470,n11114 );
   nor U11536 ( n11519,n11520,n11459 );
   nor U11537 ( n11518,p2_reg3_reg_3_,n11472 );
   and U11538 ( n11517,n11088,n11455 );
   nand U11539 ( n11088,n11521,n11522,n11523 );
   nand U11540 ( n11523,n11477,n10657 );
   nand U11541 ( n11522,n11524,n11525 );
   nand U11542 ( n11525,n11526,n11527 );
   nand U11543 ( n11527,n11528,n11529 );
   nand U11544 ( n11526,n11530,n11529 );
   nand U11545 ( n11521,n11531,n11449,n11532 );
   nor U11546 ( n11516,n11533,n11455 );
   nand U11547 ( n11514,n11461,n10651 );
   nand U11548 ( n11513,n11479,n11091 );
   xor U11549 ( n11091,n11090,n11509 );
   nand U11550 ( n11512,n11092,n11480 );
   xor U11551 ( n11092,n11534,n11532 );
   nor U11552 ( n11534,n11535,n11536 );
   and U11553 ( n11535,n11537,n11507 );
   nor U11554 ( n11545,n11546,n11459 );
   and U11555 ( n11544,n10648,n11461 );
   and U11556 ( n11543,n11076,n11455 );
   nand U11557 ( n11076,n11547,n11548 );
   nand U11558 ( n11548,n11549,n11550,n11449 );
   nand U11559 ( n11550,n11551,n11552 );
   nand U11560 ( n11549,n11553,n11554,n11555 );
   nand U11561 ( n11547,n11477,n10654 );
   nor U11562 ( n11542,n11556,n11455 );
   nand U11563 ( n11540,n11479,n11078 );
   and U11564 ( n11078,n11557,n11558 );
   nand U11565 ( n11558,n11080,n11559 );
   nand U11566 ( n11559,n11560,n11520 );
   nand U11567 ( n11539,n11457,n11561 );
   nand U11568 ( n11538,n11079,n11480 );
   xor U11569 ( n11079,n11551,n11562 );
   nor U11570 ( n11570,n11068,n11459 );
   and U11571 ( n11569,n11571,n11457 );
   nor U11572 ( n11568,n11060,n11445 );
   and U11573 ( n11060,n11572,n11573 );
   nand U11574 ( n11573,n11574,n11449,n11575 );
   nand U11575 ( n11575,n11576,n11577 );
   nand U11576 ( n11574,n11578,n11579 );
   nand U11577 ( n11572,n11477,n10651 );
   nor U11578 ( n11567,n11580,n11455 );
   nand U11579 ( n11565,n11461,n10645 );
   xor U11580 ( n11067,n11581,n11582 );
   nand U11581 ( n11563,n11066,n11480 );
   xor U11582 ( n11066,n11583,n11577 );
   not U11583 ( n11577,n11584 );
   nor U11584 ( n11583,n11585,n11586 );
   nor U11585 ( n11585,n11587,n11562 );
   nor U11586 ( n11595,n11596,n11459 );
   and U11587 ( n11594,n11597,n11457 );
   and U11588 ( n11593,n11053,n11455 );
   nand U11589 ( n11053,n11598,n11599,n11600 );
   nand U11590 ( n11600,n11477,n10648 );
   nand U11591 ( n11599,n11601,n11449,n11602 );
   nand U11592 ( n11598,n11603,n11604,n11449 );
   nand U11593 ( n11604,n11578,n11605 );
   nand U11594 ( n11603,n11606,n11607 );
   nand U11595 ( n11606,n11608,n11609 );
   nor U11596 ( n11592,n11610,n11455 );
   nand U11597 ( n11590,n11461,n10642 );
   nand U11598 ( n11589,n11056,n11480 );
   xor U11599 ( n11056,n11601,n11611 );
   not U11600 ( n11601,n11605 );
   nand U11601 ( n11588,n11479,n11055 );
   and U11602 ( n11055,n11612,n11613 );
   nand U11603 ( n11613,n11614,n11057 );
   nand U11604 ( n11614,n11581,n11068 );
   nor U11605 ( n11622,n11623,n11459 );
   and U11606 ( n11621,n11624,n11457 );
   and U11607 ( n11620,n11040,n11455 );
   nand U11608 ( n11040,n11625,n11626 );
   nand U11609 ( n11626,n11627,n11628,n11496 );
   nand U11610 ( n11496,n11629,n11630,n11631,n11632 );
   nand U11611 ( n11628,n11633,n11634 );
   nand U11612 ( n11627,n11635,n11636 );
   nand U11613 ( n11625,n11477,n10645 );
   nor U11614 ( n11619,n11637,n11455 );
   nand U11615 ( n11617,n11461,n10639 );
   nand U11616 ( n11616,n11044,n11043,n11480 );
   nand U11617 ( n11043,n11638,n11639,n11635 );
   or U11618 ( n11638,n11611,n11640 );
   nand U11619 ( n11044,n11641,n11642,n11643 );
   nand U11620 ( n11641,n11611,n11639 );
   nand U11621 ( n11615,n11479,n11045 );
   xor U11622 ( n11045,n11623,n11644 );
   nor U11623 ( n11652,n11031,n11459 );
   nor U11624 ( n11651,n11653,n11472 );
   nor U11625 ( n11650,n11024,n11445 );
   and U11626 ( n11024,n11654,n11655,n11656,n11657 );
   nor U11627 ( n11657,n11658,n11659,n11660,n11661 );
   nor U11628 ( n11661,n11662,n11629 );
   xor U11629 ( n11662,n11663,n11664 );
   nor U11630 ( n11660,n11665,n11630 );
   nor U11631 ( n11665,n11666,n11667 );
   not U11632 ( n11667,n11668 );
   nor U11633 ( n11666,n11663,n11664 );
   nor U11634 ( n11659,n11669,n11030 );
   nor U11635 ( n11658,n11054,n11670 );
   nand U11636 ( n11656,n11671,n11672 );
   nand U11637 ( n11655,n11673,n11674 );
   nand U11638 ( n11674,n11675,n11668 );
   nand U11639 ( n11668,n11663,n11664 );
   or U11640 ( n11675,n11664,n11663 );
   nand U11641 ( n11673,n11631,n11632 );
   nand U11642 ( n11654,n11671,n11676 );
   and U11643 ( n11649,p2_reg2_reg_8_,n11445 );
   nand U11644 ( n11647,n11461,n10636 );
   or U11645 ( n11646,n11460,n11032 );
   nand U11646 ( n11032,n11677,n11678 );
   nand U11647 ( n11678,n11679,n11680 );
   nand U11648 ( n11680,n11644,n11623 );
   nand U11649 ( n11645,n11681,n11671 );
   not U11650 ( n11671,n11030 );
   xor U11651 ( n11030,n11664,n11682 );
   nor U11652 ( n11690,n11691,n11459 );
   and U11653 ( n11689,n11692,n11457 );
   and U11654 ( n11688,n11016,n11455 );
   nand U11655 ( n11016,n11693,n11694 );
   nand U11656 ( n11694,n11695,n11696,n11449 );
   nand U11657 ( n11696,n11697,n11698,n11699 );
   or U11658 ( n11695,n11700,n11699 );
   nand U11659 ( n11693,n11477,n10639 );
   nor U11660 ( n11687,n11701,n11455 );
   nand U11661 ( n11685,n11461,n10633 );
   nand U11662 ( n11684,n11479,n11019 );
   xor U11663 ( n11019,n11677,n11018 );
   nand U11664 ( n11683,n11020,n11480 );
   nand U11665 ( n11480,n11456,n11702 );
   nand U11666 ( n11702,n11455,n11117 );
   or U11667 ( n11117,n11703,n11704 );
   xor U11668 ( n11020,n11700,n11705 );
   nor U11669 ( n11710,n11007,n11459 );
   and U11670 ( n11709,n11711,n11457 );
   nor U11671 ( n11708,n11000,n11445 );
   and U11672 ( n11000,n11712,n11713,n11714,n11715 );
   nor U11673 ( n11715,n11716,n11717,n11718,n11719 );
   nor U11674 ( n11719,n11632,n11720 );
   nor U11675 ( n11718,n11721,n11006 );
   nor U11676 ( n11717,n11722,n11006 );
   nor U11677 ( n11716,n11669,n11006 );
   nand U11678 ( n11714,n11723,n11724 );
   nand U11679 ( n11713,n11723,n11725 );
   nand U11680 ( n11725,n11629,n11630 );
   not U11681 ( n11723,n11720 );
   nand U11682 ( n11720,n11726,n11727 );
   nand U11683 ( n11727,n11728,n11729,n11730 );
   nand U11684 ( n11726,n11731,n11732 );
   nand U11685 ( n11712,n11477,n10636 );
   nor U11686 ( n11707,n11733,n11455 );
   nand U11687 ( n11008,n11734,n11735 );
   nand U11688 ( n11735,n11736,n11737 );
   nand U11689 ( n11736,n11738,n11691 );
   nand U11690 ( n11006,n11739,n11740 );
   nand U11691 ( n11740,n11741,n11742,n11743 );
   nand U11692 ( n11739,n11744,n11745,n11731 );
   not U11693 ( n11731,n11743 );
   nand U11694 ( n11744,n11705,n11742 );
   not U11695 ( n11705,n11746 );
   nor U11696 ( n11751,n10995,n11459 );
   nor U11697 ( n11750,n11752,n11472 );
   nor U11698 ( n11749,n10989,n11445 );
   and U11699 ( n10989,n11753,n11754 );
   nor U11700 ( n11754,n11755,n11756,n11757,n11758 );
   nor U11701 ( n11758,n11759,n11630 );
   nor U11702 ( n11757,n11669,n10997 );
   nor U11703 ( n11756,n11017,n11670 );
   nor U11704 ( n11755,n11759,n11631 );
   nor U11705 ( n11753,n11760,n11761,n11762,n11763 );
   nor U11706 ( n11763,n11759,n11632 );
   and U11707 ( n11759,n11764,n11765,n11766 );
   not U11708 ( n11766,n11767 );
   nand U11709 ( n11765,n11768,n11730 );
   nand U11710 ( n11764,n11732,n11769 );
   not U11711 ( n11732,n11730 );
   nor U11712 ( n11762,n11721,n10997 );
   nor U11713 ( n11761,n11722,n10997 );
   nor U11714 ( n11760,n11770,n11629 );
   nor U11715 ( n11770,n11767,n11771,n11772 );
   nor U11716 ( n11772,n11773,n11730 );
   and U11717 ( n11771,n11730,n11768 );
   nand U11718 ( n11767,n11774,n11775 );
   nand U11719 ( n11775,n11776,n11769 );
   not U11720 ( n11769,n11773 );
   nand U11721 ( n11773,n11777,n11778 );
   nand U11722 ( n11774,n11779,n11768 );
   nor U11723 ( n11768,n11780,n11776 );
   nor U11724 ( n11748,n11781,n11455 );
   xor U11725 ( n10996,n11782,n11783 );
   xor U11726 ( n10997,n11780,n11784 );
   nor U11727 ( n11792,n10985,n11459 );
   nor U11728 ( n11791,n11793,n11472 );
   nor U11729 ( n11790,n10978,n11445 );
   and U11730 ( n10978,n11794,n11795,n11796,n11797 );
   nor U11731 ( n11797,n11798,n11799,n11800,n11801 );
   nor U11732 ( n11801,n11802,n11670 );
   nor U11733 ( n11800,n11722,n10984 );
   nor U11734 ( n11799,n11629,n11803 );
   nor U11735 ( n11798,n11631,n11803 );
   nor U11736 ( n11796,n11804,n11805 );
   nor U11737 ( n11805,n11669,n10984 );
   nor U11738 ( n11804,n11632,n11803 );
   or U11739 ( n11795,n11803,n11630 );
   xor U11740 ( n11803,n11806,n11807 );
   nand U11741 ( n11794,n11808,n11672 );
   nor U11742 ( n11789,n11809,n11455 );
   nand U11743 ( n11787,n11461,n10624 );
   or U11744 ( n11786,n11460,n10986 );
   nand U11745 ( n10986,n11810,n11811 );
   nand U11746 ( n11811,n11812,n11813 );
   nand U11747 ( n11813,n11783,n10995 );
   nand U11748 ( n11785,n11681,n11808 );
   not U11749 ( n11808,n10984 );
   xor U11750 ( n10984,n11806,n11814 );
   nor U11751 ( n11819,n10973,n11459 );
   nor U11752 ( n11818,n11820,n11472 );
   nor U11753 ( n11817,n10967,n11445 );
   and U11754 ( n10967,n11821,n11822,n11823,n11824 );
   nor U11755 ( n11824,n11825,n11826,n11827,n11828 );
   nor U11756 ( n11828,n11721,n10975 );
   nor U11757 ( n11827,n11722,n10975 );
   nor U11758 ( n11826,n11669,n10975 );
   nor U11759 ( n11825,n11629,n11829 );
   nor U11760 ( n11823,n11830,n11831 );
   nor U11761 ( n11831,n11832,n11670 );
   nor U11762 ( n11830,n11632,n11829 );
   nand U11763 ( n11822,n11833,n11724 );
   nand U11764 ( n11821,n11833,n11528 );
   not U11765 ( n11833,n11829 );
   xor U11766 ( n11829,n11834,n11835 );
   nor U11767 ( n11816,n11836,n11455 );
   xor U11768 ( n10974,n11837,n10973 );
   nand U11769 ( n10975,n11838,n11839 );
   nand U11770 ( n11839,n11840,n11841,n11842 );
   nand U11771 ( n11840,n11843,n11844 );
   nand U11772 ( n11838,n11834,n11844,n11845 );
   nand U11773 ( n11845,n11846,n11814 );
   not U11774 ( n11814,n11843 );
   nor U11775 ( n11843,n11847,n11848 );
   nor U11776 ( n11853,n10963,n11459 );
   nor U11777 ( n11852,n11854,n11472 );
   nor U11778 ( n11851,n10956,n11445 );
   and U11779 ( n10956,n11855,n11856 );
   nor U11780 ( n11856,n11857,n11858,n11859,n11860 );
   nor U11781 ( n11860,n11721,n10962 );
   nor U11782 ( n11859,n11861,n11630 );
   nor U11783 ( n11858,n11631,n11862,n11863 );
   nor U11784 ( n11863,n11864,n11865 );
   nor U11785 ( n11862,n11866,n11867 );
   nor U11786 ( n11857,n11669,n10962 );
   nor U11787 ( n11855,n11868,n11869,n11870,n11871 );
   nor U11788 ( n11871,n11722,n10962 );
   nor U11789 ( n11870,n11872,n11670 );
   nor U11790 ( n11869,n11861,n11632 );
   nor U11791 ( n11868,n11861,n11629 );
   and U11792 ( n11861,n11873,n11874 );
   nand U11793 ( n11874,n11866,n11875 );
   nand U11794 ( n11875,n11876,n11877 );
   nand U11795 ( n11873,n11867,n11878 );
   nor U11796 ( n11850,n11879,n11455 );
   nand U11797 ( n10964,n11880,n11881 );
   nand U11798 ( n11881,n11882,n11883 );
   nand U11799 ( n11882,n11837,n10973 );
   xor U11800 ( n10962,n11884,n11867 );
   nor U11801 ( n11892,n10951,n11459 );
   and U11802 ( n11891,n11893,n11457 );
   nor U11803 ( n11890,n10945,n11445 );
   and U11804 ( n10945,n11894,n11895,n11896,n11897 );
   nor U11805 ( n11897,n11898,n11899,n11900,n11901 );
   nor U11806 ( n11901,n11721,n10953 );
   nor U11807 ( n11900,n11630,n11902 );
   nor U11808 ( n11899,n11631,n11902 );
   nor U11809 ( n11898,n11669,n10953 );
   nor U11810 ( n11896,n11903,n11904 );
   nor U11811 ( n11904,n11632,n11902 );
   nor U11812 ( n11903,n11629,n11902 );
   nand U11813 ( n11902,n11905,n11906 );
   nand U11814 ( n11906,n11907,n11908 );
   nand U11815 ( n11905,n11909,n11910 );
   nand U11816 ( n11895,n11477,n10621 );
   nand U11817 ( n11894,n11911,n11676 );
   nor U11818 ( n11889,n11912,n11455 );
   nand U11819 ( n11887,n11461,n10615 );
   xor U11820 ( n10952,n11913,n11914 );
   nand U11821 ( n11885,n11681,n11911 );
   not U11822 ( n11911,n10953 );
   xor U11823 ( n10953,n11915,n11909 );
   nor U11824 ( n11923,n10941,n11459 );
   nor U11825 ( n11922,n11924,n11472 );
   nor U11826 ( n11921,n10934,n11445 );
   and U11827 ( n10934,n11925,n11926,n11927,n11928 );
   nor U11828 ( n11928,n11929,n11930,n11931,n11932 );
   nor U11829 ( n11932,n10942,n11722 );
   nor U11830 ( n11931,n10942,n11669 );
   not U11831 ( n10942,n11933 );
   nor U11832 ( n11930,n11934,n11632 );
   nor U11833 ( n11929,n11630,n11935,n11936 );
   nor U11834 ( n11936,n11937,n11938 );
   nor U11835 ( n11938,n11939,n11940,n11941 );
   and U11836 ( n11941,n11908,n11910 );
   and U11837 ( n11935,n11939,n11907 );
   nor U11838 ( n11927,n11942,n11943 );
   nor U11839 ( n11943,n11934,n11631 );
   not U11840 ( n11934,n11944 );
   nor U11841 ( n11942,n11945,n11670 );
   nand U11842 ( n11926,n11672,n11933 );
   nand U11843 ( n11925,n11946,n11944 );
   nand U11844 ( n11944,n11947,n11948,n11949,n11950 );
   nand U11845 ( n11950,n11951,n11907 );
   nor U11846 ( n11907,n11910,n11940 );
   nand U11847 ( n11949,n11910,n11937 );
   nor U11848 ( n11910,n11952,n11864 );
   nand U11849 ( n11948,n11940,n11937 );
   and U11850 ( n11937,n11908,n11953,n11954 );
   or U11851 ( n11947,n11908,n11939 );
   nor U11852 ( n11920,n11955,n11455 );
   nand U11853 ( n11918,n11461,n10612 );
   nand U11854 ( n11917,n11681,n11933 );
   xor U11855 ( n11933,n11951,n11956 );
   nand U11856 ( n11916,n11479,n10938 );
   and U11857 ( n10938,n11957,n11958 );
   nand U11858 ( n11958,n11959,n11960 );
   nand U11859 ( n11960,n11914,n10951 );
   nor U11860 ( n11968,n10929,n11459 );
   nor U11861 ( n11967,n11969,n11472 );
   nor U11862 ( n11966,n10923,n11445 );
   and U11863 ( n10923,n11970,n11971,n11972,n11973 );
   nor U11864 ( n11973,n11974,n11975,n11976,n11977 );
   nor U11865 ( n11977,n11978,n11630 );
   nor U11866 ( n11976,n11978,n11631 );
   nor U11867 ( n11975,n11979,n11670 );
   nor U11868 ( n11974,n11978,n11632 );
   nor U11869 ( n11972,n11980,n11981 );
   nor U11870 ( n11981,n11669,n10931 );
   nor U11871 ( n11980,n11978,n11629 );
   xor U11872 ( n11978,n11982,n11983 );
   nand U11873 ( n11971,n11984,n11676 );
   nand U11874 ( n11970,n11984,n11672 );
   nor U11875 ( n11965,n11985,n11455 );
   nand U11876 ( n11963,n11461,n10609 );
   xor U11877 ( n10930,n11986,n11987 );
   nand U11878 ( n11961,n11681,n11984 );
   not U11879 ( n11984,n10931 );
   nand U11880 ( n10931,n11988,n11989 );
   nand U11881 ( n11989,n11990,n11991,n11992 );
   nand U11882 ( n11988,n11993,n11994,n11982 );
   nand U11883 ( n11993,n11995,n11991 );
   nor U11884 ( n12000,n10918,n11459 );
   nor U11885 ( n11999,n12001,n11472 );
   nor U11886 ( n11998,n10912,n11445 );
   and U11887 ( n10912,n12002,n12003,n12004,n12005 );
   nor U11888 ( n12005,n12006,n12007,n12008,n12009 );
   nor U11889 ( n12009,n11722,n10919 );
   nor U11890 ( n12008,n12010,n11670 );
   nor U11891 ( n12007,n11629,n12011 );
   nor U11892 ( n12006,n11721,n10919 );
   nor U11893 ( n12004,n12012,n12013 );
   nor U11894 ( n12013,n11669,n10919 );
   nor U11895 ( n12012,n11632,n12011 );
   not U11896 ( n12011,n12014 );
   nand U11897 ( n12003,n12014,n11528 );
   nand U11898 ( n12002,n12014,n11724 );
   xor U11899 ( n12014,n12015,n12016 );
   nor U11900 ( n11997,n12017,n11455 );
   xor U11901 ( n10919,n12015,n12018 );
   nand U11902 ( n10920,n12019,n12020 );
   nand U11903 ( n12020,n12021,n12022 );
   nand U11904 ( n12022,n11987,n10929 );
   nor U11905 ( n12026,n10907,n11459 );
   nor U11906 ( n12025,n12027,n11472 );
   nor U11907 ( n12024,n10901,n11445 );
   and U11908 ( n10901,n12028,n12029,n12030,n12031 );
   nor U11909 ( n12031,n12032,n12033,n12034,n12035 );
   nor U11910 ( n12035,n11722,n10909 );
   nor U11911 ( n12034,n12036,n11670 );
   nor U11912 ( n12033,n11629,n12037 );
   nor U11913 ( n12032,n11721,n10909 );
   nor U11914 ( n12030,n12038,n12039 );
   nor U11915 ( n12039,n11669,n10909 );
   nor U11916 ( n12038,n11632,n12037 );
   not U11917 ( n12037,n12040 );
   nand U11918 ( n12029,n12040,n11528 );
   nand U11919 ( n12028,n12040,n11724 );
   xor U11920 ( n12040,n12041,n12042 );
   nor U11921 ( n12023,n12043,n11455 );
   xor U11922 ( n10908,n12044,n12045 );
   xor U11923 ( n10909,n12041,n12046 );
   nor U11924 ( n12051,n10897,n11459 );
   nor U11925 ( n12050,n12052,n11472 );
   nor U11926 ( n12049,n10890,n11445 );
   and U11927 ( n10890,n12053,n12054,n12055,n12056 );
   nor U11928 ( n12056,n12057,n12058,n12059,n12060 );
   nor U11929 ( n12060,n11630,n12061 );
   nor U11930 ( n12059,n11631,n12061 );
   nor U11931 ( n12058,n12062,n11670 );
   nor U11932 ( n12057,n11632,n12061 );
   nor U11933 ( n12055,n12063,n12064 );
   nor U11934 ( n12064,n11669,n10896 );
   nor U11935 ( n12063,n11629,n12061 );
   xor U11936 ( n12061,n12065,n12066 );
   nand U11937 ( n12054,n12067,n12068,n11676 );
   nand U11938 ( n12053,n12067,n12068,n11672 );
   and U11939 ( n12048,p2_reg2_reg_20_,n11445 );
   nand U11940 ( n10898,n12069,n12070 );
   nand U11941 ( n12070,n12071,n12072 );
   nand U11942 ( n12072,n12045,n10907 );
   nand U11943 ( n10896,n12067,n12068 );
   nand U11944 ( n12068,n12065,n12073,n12074 );
   nand U11945 ( n12074,n12075,n12076 );
   nand U11946 ( n12067,n12077,n12078,n12079 );
   nand U11947 ( n12077,n12046,n12073 );
   nor U11948 ( n12084,n10885,n11459 );
   and U11949 ( n12083,n12085,n11457 );
   nor U11950 ( n12082,n10879,n11445 );
   and U11951 ( n10879,n12086,n12087 );
   nor U11952 ( n12087,n12088,n12089,n12090,n12091 );
   nor U11953 ( n12091,n11631,n12092 );
   nor U11954 ( n12090,n11722,n10887 );
   nor U11955 ( n12089,n11629,n12092 );
   nor U11956 ( n12088,n12093,n12094,n12095,n11721 );
   nor U11957 ( n12095,n12096,n12097 );
   not U11958 ( n12097,n12098 );
   nor U11959 ( n12096,n12046,n12099 );
   nor U11960 ( n12094,n12100,n12101 );
   nor U11961 ( n12086,n12102,n12103,n12104,n12105 );
   nor U11962 ( n12105,n11669,n10887 );
   nor U11963 ( n12104,n11630,n12092 );
   nor U11964 ( n12103,n12106,n11670 );
   nor U11965 ( n12102,n11632,n12092 );
   nand U11966 ( n12092,n12107,n12108 );
   nand U11967 ( n12108,n12109,n12110 );
   nand U11968 ( n12107,n12111,n12112 );
   and U11969 ( n12081,p2_reg2_reg_21_,n11445 );
   xor U11970 ( n10886,n12113,n12114 );
   nand U11971 ( n10887,n12115,n12116,n12117 );
   nand U11972 ( n12117,n12111,n12118 );
   not U11973 ( n12116,n12093 );
   nor U11974 ( n12093,n12099,n12046,n12101 );
   nand U11975 ( n12115,n12098,n12119 );
   nand U11976 ( n12119,n12079,n12076 );
   not U11977 ( n12076,n12046 );
   nor U11978 ( n12046,n12120,n12121 );
   nor U11979 ( n12098,n12118,n12111 );
   nor U11980 ( n12125,n12126,n12127,n12128,n12129 );
   nor U11981 ( n12129,n10875,n11459 );
   nor U11982 ( n12128,n12130,n11472 );
   nor U11983 ( n12127,n10868,n11445 );
   and U11984 ( n10868,n12131,n12132,n12133,n12134 );
   nor U11985 ( n12134,n12135,n12136,n12137,n12138 );
   nor U11986 ( n12138,n11722,n10874 );
   nor U11987 ( n12137,n12139,n11670 );
   nor U11988 ( n12136,n11632,n12140 );
   nor U11989 ( n12135,n11629,n12140 );
   nor U11990 ( n12133,n12141,n12142 );
   nor U11991 ( n12142,n11631,n12140 );
   nor U11992 ( n12141,n11669,n10874 );
   or U11993 ( n12132,n12140,n11630 );
   nand U11994 ( n12140,n12143,n12144 );
   nand U11995 ( n12144,n12145,n12146,n12147 );
   nand U11996 ( n12143,n12148,n12149 );
   nand U11997 ( n12131,n12150,n11672 );
   and U11998 ( n12126,p2_reg2_reg_22_,n11445 );
   nand U11999 ( n12124,n11461,n10594 );
   or U12000 ( n12123,n11460,n10876 );
   nand U12001 ( n10876,n12151,n12152 );
   nand U12002 ( n12152,n12153,n12154 );
   nand U12003 ( n12154,n12113,n10885 );
   nand U12004 ( n12122,n11681,n12150 );
   not U12005 ( n12150,n10874 );
   xor U12006 ( n10874,n12148,n12155 );
   nor U12007 ( n12160,n10863,n11459 );
   and U12008 ( n12159,n12161,n11457 );
   nor U12009 ( n12158,n10857,n11445 );
   and U12010 ( n10857,n12162,n12163,n12164,n12165 );
   nor U12011 ( n12165,n12166,n12167,n12168,n12169 );
   nor U12012 ( n12169,n10865,n11669 );
   nor U12013 ( n12168,n10865,n11721 );
   nor U12014 ( n12167,n12170,n11670 );
   nor U12015 ( n12166,n12171,n11631 );
   nor U12016 ( n12164,n12172,n12173 );
   nor U12017 ( n12173,n12171,n11629 );
   nor U12018 ( n12172,n12171,n11632 );
   and U12019 ( n12171,n12174,n12175 );
   nand U12020 ( n12174,n12176,n12177 );
   nand U12021 ( n12177,n12146,n12147 );
   nand U12022 ( n12163,n11676,n12178 );
   xor U12023 ( n12178,n12179,n12180 );
   nand U12024 ( n12162,n12181,n12182,n11528 );
   nand U12025 ( n12182,n12147,n12146,n12180 );
   not U12026 ( n12147,n12149 );
   nand U12027 ( n12181,n12175,n12183 );
   not U12028 ( n12183,n12176 );
   nor U12029 ( n12176,n12184,n12185 );
   nand U12030 ( n12175,n12186,n12187 );
   nand U12031 ( n12187,n12149,n12145 );
   nor U12032 ( n12149,n12109,n12188 );
   and U12033 ( n12186,n12185,n12146 );
   and U12034 ( n12157,p2_reg2_reg_23_,n11445 );
   xor U12035 ( n10864,n12189,n12190 );
   xor U12036 ( n10865,n12179,n12185 );
   nor U12037 ( n12194,n12195,n12196,n12197,n12198 );
   nor U12038 ( n12198,n12199,n11459 );
   and U12039 ( n12197,n12200,n11457 );
   and U12040 ( n12196,n10849,n11455 );
   nand U12041 ( n10849,n12201,n12202,n12203,n12204 );
   nand U12042 ( n12204,n10854,n11703 );
   nand U12043 ( n12203,n12205,n11449 );
   xor U12044 ( n12205,n12206,n12207 );
   nand U12045 ( n12202,n11704,n10854 );
   nand U12046 ( n12201,n11477,n10594 );
   and U12047 ( n12195,p2_reg2_reg_24_,n11445 );
   nand U12048 ( n12193,n11461,n10588 );
   nand U12049 ( n12192,n11479,n10852 );
   and U12050 ( n10852,n12208,n12209 );
   nand U12051 ( n12209,n10853,n12210 );
   nand U12052 ( n12210,n12189,n10863 );
   nand U12053 ( n12191,n11681,n10854 );
   xor U12054 ( n10854,n12206,n12211 );
   nor U12055 ( n12216,n10841,n11459 );
   and U12056 ( n12215,n12217,n11457 );
   nor U12057 ( n12214,n10833,n11445 );
   and U12058 ( n10833,n12218,n12219,n12220,n12221 );
   nor U12059 ( n12221,n12222,n12223,n12224,n12225 );
   nor U12060 ( n12225,n10840,n11722 );
   nor U12061 ( n12224,n12226,n11670 );
   nor U12062 ( n12223,n11629,n12227 );
   nor U12063 ( n12222,n10840,n11721 );
   nor U12064 ( n12220,n12228,n12229 );
   nor U12065 ( n12229,n10840,n11669 );
   nor U12066 ( n12228,n11632,n12227 );
   nand U12067 ( n12219,n12230,n11528 );
   nand U12068 ( n12218,n12230,n11724 );
   not U12069 ( n12230,n12227 );
   xor U12070 ( n12227,n12231,n12232 );
   and U12071 ( n12213,p2_reg2_reg_25_,n11445 );
   xor U12072 ( n10840,n12233,n12232 );
   xor U12073 ( n10839,n12234,n12235 );
   nor U12074 ( n12240,n10829,n11459 );
   nor U12075 ( n12239,n12241,n11472 );
   nor U12076 ( n12238,n10822,n11445 );
   and U12077 ( n10822,n12242,n12243,n12244,n12245 );
   nor U12078 ( n12245,n12246,n12247,n12248,n12249 );
   nor U12079 ( n12249,n11629,n12250 );
   nor U12080 ( n12248,n11631,n12250 );
   nor U12081 ( n12247,n10850,n11670 );
   nor U12082 ( n12246,n11632,n12250 );
   nor U12083 ( n12244,n12251,n12252 );
   nor U12084 ( n12252,n11669,n10828 );
   nor U12085 ( n12251,n11630,n12250 );
   nand U12086 ( n12250,n12253,n12254 );
   nand U12087 ( n12254,n12255,n12256 );
   nand U12088 ( n12253,n12257,n12258,n12259 );
   nand U12089 ( n12243,n12260,n12261,n11676 );
   nand U12090 ( n12242,n12260,n12261,n11672 );
   and U12091 ( n12237,p2_reg2_reg_26_,n11445 );
   nand U12092 ( n10830,n12262,n12263 );
   nand U12093 ( n12263,n12264,n12265 );
   nand U12094 ( n12265,n12234,n10841 );
   nand U12095 ( n10828,n12260,n12261 );
   nand U12096 ( n12261,n12266,n12267,n12268 );
   nand U12097 ( n12268,n12233,n12269 );
   not U12098 ( n12233,n12270 );
   nand U12099 ( n12260,n12271,n12272 );
   nand U12100 ( n12272,n12267,n12270 );
   nand U12101 ( n12270,n12273,n12274 );
   nand U12102 ( n12274,n12211,n12275 );
   and U12103 ( n12271,n12255,n12269 );
   not U12104 ( n12255,n12266 );
   nor U12105 ( n12280,n10817,n11459 );
   and U12106 ( n12279,n12281,n11457 );
   nor U12107 ( n12278,n10811,n11445 );
   and U12108 ( n10811,n12282,n12283,n12284,n12285 );
   nor U12109 ( n12285,n12286,n12287 );
   nor U12110 ( n12287,n12288,n11670 );
   nor U12111 ( n12286,n11669,n10819 );
   nand U12112 ( n12284,n12289,n11703 );
   xor U12113 ( n12289,n12290,n12291 );
   nand U12114 ( n12283,n12292,n12293,n11528 );
   nand U12115 ( n12293,n12291,n12294 );
   nand U12116 ( n12292,n12295,n12296 );
   nand U12117 ( n12296,n12258,n12297 );
   nand U12118 ( n12297,n12256,n12257 );
   nand U12119 ( n12282,n12298,n11530 );
   xor U12120 ( n12298,n12291,n12294 );
   and U12121 ( n12277,p2_reg2_reg_27_,n11445 );
   xor U12122 ( n10818,n12299,n12300 );
   xor U12123 ( n10819,n12290,n12295 );
   not U12124 ( n12295,n12291 );
   nor U12125 ( n12290,n12301,n12302 );
   nand U12126 ( n12302,n12303,n12304 );
   nand U12127 ( n12304,n12305,n12306 );
   nor U12128 ( n12310,n12311,n12312,n12313,n12314 );
   nor U12129 ( n12314,n10804,n11459 );
   and U12130 ( n12313,n12315,n11457 );
   nor U12131 ( n12312,n10797,n11445 );
   and U12132 ( n10797,n12316,n12317,n12318,n12319 );
   nor U12133 ( n12319,n12320,n12321,n12322,n12323 );
   nor U12134 ( n12323,n12324,n11670 );
   nor U12135 ( n12322,n11721,n12325 );
   nor U12136 ( n12321,n12326,n11629 );
   nor U12137 ( n12320,n12326,n11631 );
   nor U12138 ( n12318,n12327,n12328 );
   nor U12139 ( n12328,n12326,n11632 );
   not U12140 ( n12326,n12330 );
   nor U12141 ( n12327,n11722,n12325 );
   xor U12142 ( n12325,n12331,n12332 );
   nand U12143 ( n12317,n11528,n12330 );
   xor U12144 ( n12330,n12332,n12333 );
   nand U12145 ( n12316,n10806,n11704 );
   not U12146 ( n11704,n11669 );
   and U12147 ( n12311,p2_reg2_reg_28_,n11445 );
   nand U12148 ( n10807,n12334,n12335 );
   nand U12149 ( n12335,n12336,n12337 );
   nand U12150 ( n12337,n12299,n10817 );
   not U12151 ( n12334,n12338 );
   nand U12152 ( n12308,n11681,n10806 );
   xor U12153 ( n10806,n12339,n12332 );
   not U12154 ( n11681,n11456 );
   nand U12155 ( n12307,n11461,n10576 );
   not U12156 ( n10851,n10808 );
   nor U12157 ( n12346,n10789,n11460 );
   xor U12158 ( n10789,n10791,n12338 );
   and U12159 ( n12345,n12347,n11457 );
   nor U12160 ( n12344,n10793,n11456 );
   nand U12161 ( n11456,n12348,n11455,n12349 );
   nand U12162 ( n12342,n12350,n10791 );
   nand U12163 ( n12341,n11445,p2_reg2_reg_29_ );
   nand U12164 ( n12340,n11455,n10794 );
   nand U12165 ( n10794,n12351,n12352,n12353,n12354 );
   nor U12166 ( n12354,n12355,n12356 );
   and U12167 ( n12356,n10573,n12357 );
   nor U12168 ( n12355,n10793,n11669 );
   xor U12169 ( n10793,n12358,n12359 );
   nand U12170 ( n12359,n12360,n12361 );
   nand U12171 ( n12361,n12339,n12362 );
   and U12172 ( n12339,n12363,n12364 );
   nand U12173 ( n12353,n11477,n10579 );
   nor U12174 ( n11477,n12365,n12366 );
   nand U12175 ( n12352,n12367,n11703 );
   nand U12176 ( n11703,n11721,n11722 );
   nor U12177 ( n11676,n11138,n11137 );
   xor U12178 ( n12367,n12368,n12369 );
   nand U12179 ( n12369,n12360,n12370 );
   nand U12180 ( n12370,n12339,n12362 );
   nand U12181 ( n12331,n12363,n12364 );
   nand U12182 ( n12364,n12301,n12371 );
   nor U12183 ( n12301,n12211,n12372 );
   nand U12184 ( n12372,n12305,n12273 );
   nand U12185 ( n12211,n12373,n12374 );
   nand U12186 ( n12374,n12375,n12179 );
   nand U12187 ( n12179,n12376,n12377 );
   nand U12188 ( n12377,n12155,n12378 );
   and U12189 ( n12155,n12379,n12380,n12381 );
   nand U12190 ( n12381,n12382,n12383 );
   nand U12191 ( n12383,n12100,n12384 );
   nand U12192 ( n12384,n12121,n12079 );
   not U12193 ( n12100,n12118 );
   nand U12194 ( n12118,n12078,n12385 );
   nand U12195 ( n12385,n12386,n12387 );
   nand U12196 ( n12379,n12120,n12382,n12079 );
   not U12197 ( n12079,n12099 );
   nand U12198 ( n12099,n12075,n12387 );
   nor U12199 ( n12120,n12018,n12388 );
   and U12200 ( n12018,n12389,n12390 );
   nand U12201 ( n12390,n12391,n12392 );
   nand U12202 ( n12391,n11991,n11990 );
   nand U12203 ( n11990,n11956,n11994 );
   not U12204 ( n11956,n11995 );
   nand U12205 ( n11995,n12393,n12394 );
   nand U12206 ( n12394,n12395,n10951 );
   or U12207 ( n12395,n11915,n11945 );
   nand U12208 ( n12393,n11945,n11915 );
   nand U12209 ( n11915,n12396,n12397 );
   nand U12210 ( n12397,n10963,n12398 );
   nand U12211 ( n12398,n10621,n11884 );
   or U12212 ( n12396,n11884,n10621 );
   nand U12213 ( n11884,n12399,n12400 );
   nand U12214 ( n12400,n12401,n12402 );
   nand U12215 ( n12401,n11844,n11841,n12403 );
   nand U12216 ( n12403,n11848,n11842 );
   nand U12217 ( n12399,n11847,n11842 );
   and U12218 ( n11842,n12402,n11846 );
   and U12219 ( n11847,n11784,n12404 );
   nand U12220 ( n12404,n11802,n10995 );
   nand U12221 ( n11784,n12405,n12406 );
   nand U12222 ( n12406,n12407,n12408 );
   nand U12223 ( n12407,n11742,n11741 );
   nand U12224 ( n11741,n11745,n11746 );
   nand U12225 ( n11746,n12409,n12410 );
   nand U12226 ( n12409,n11682,n12411 );
   nand U12227 ( n11682,n12412,n12413,n12414 );
   nand U12228 ( n12414,n11640,n11042 );
   nand U12229 ( n12413,n11611,n11639,n12415 );
   nand U12230 ( n12415,n11054,n11623 );
   nand U12231 ( n11611,n12416,n12417,n12418 );
   nand U12232 ( n12418,n11587,n10648 );
   nand U12233 ( n12417,n11562,n12419,n12420 );
   nand U12234 ( n12420,n11077,n11068 );
   not U12235 ( n12419,n11586 );
   nand U12236 ( n11562,n12421,n12422,n12423 );
   nand U12237 ( n12423,n11536,n10654 );
   nand U12238 ( n12422,n12424,n11537,n11507 );
   nor U12239 ( n11507,n11481,n12425 );
   nor U12240 ( n12425,n10660,n11114 );
   nand U12241 ( n12424,n11101,n11520 );
   nand U12242 ( n12421,n12426,n11090 );
   or U12243 ( n12426,n11536,n10654 );
   nand U12244 ( n11536,n12427,n12428 );
   nand U12245 ( n12428,n11508,n11537 );
   not U12246 ( n11508,n12429 );
   nand U12247 ( n12416,n11582,n12430 );
   nand U12248 ( n12430,n11077,n12431 );
   not U12249 ( n12431,n11587 );
   nand U12250 ( n12412,n12432,n10642 );
   nand U12251 ( n12432,n11623,n11642 );
   not U12252 ( n11945,n10618 );
   and U12253 ( n12363,n12433,n12434,n12435 );
   nand U12254 ( n12435,n12436,n12371 );
   nand U12255 ( n12433,n12306,n12371,n12305 );
   and U12256 ( n12305,n12269,n12437 );
   nand U12257 ( n12306,n12267,n12275 );
   nand U12258 ( n12351,n12438,n12439,n11449 );
   nand U12259 ( n11449,n12440,n11630 );
   not U12260 ( n12440,n11530 );
   nand U12261 ( n11530,n12441,n11631 );
   nor U12262 ( n11724,n11130,n12348,n11142 );
   nor U12263 ( n12441,n11946,n12329 );
   not U12264 ( n11946,n11629 );
   nand U12265 ( n12439,n12442,n12443,n12358 );
   nand U12266 ( n12442,n12333,n12444 );
   nand U12267 ( n12438,n12445,n12444,n12368 );
   or U12268 ( n12445,n12333,n12446 );
   nand U12269 ( n12333,n12447,n12448 );
   nand U12270 ( n12448,n12449,n12294 );
   nand U12271 ( n12294,n12257,n12450 );
   nand U12272 ( n12450,n12259,n12258 );
   not U12273 ( n12259,n12256 );
   nand U12274 ( n12256,n12451,n12452 );
   nand U12275 ( n12452,n12453,n12231 );
   nand U12276 ( n12231,n12454,n12455 );
   nand U12277 ( n12455,n12456,n12457 );
   not U12278 ( n12456,n12207 );
   nand U12279 ( n12207,n12458,n12459 );
   nand U12280 ( n12459,n12460,n12461 );
   nand U12281 ( n12461,n12462,n12463 );
   nand U12282 ( n12463,n12188,n12146 );
   nand U12283 ( n12458,n12109,n12464 );
   not U12284 ( n12464,n12465 );
   nor U12285 ( n12109,n12112,n12466 );
   nand U12286 ( n12112,n12467,n12468 );
   nand U12287 ( n12468,n12469,n12066 );
   nand U12288 ( n12066,n12470,n12471 );
   nand U12289 ( n12471,n12472,n12042 );
   nand U12290 ( n12042,n12473,n12474 );
   nand U12291 ( n12474,n12475,n12016 );
   nand U12292 ( n12016,n12476,n12477 );
   nand U12293 ( n12477,n11986,n12478 );
   nand U12294 ( n12478,n10612,n11983 );
   or U12295 ( n12476,n11983,n10612 );
   nand U12296 ( n11983,n12479,n12480 );
   nand U12297 ( n12480,n11953,n12481 );
   nand U12298 ( n12481,n12482,n11954 );
   not U12299 ( n12482,n12483 );
   nand U12300 ( n12479,n11952,n12484 );
   not U12301 ( n11952,n11865 );
   nand U12302 ( n11865,n11866,n11876 );
   not U12303 ( n11866,n11878 );
   nand U12304 ( n11878,n12485,n12486 );
   nand U12305 ( n12486,n12487,n11835 );
   nand U12306 ( n11835,n12488,n12489 );
   nand U12307 ( n12489,n11807,n12490 );
   nand U12308 ( n11807,n12491,n11778 );
   not U12309 ( n11778,n12492 );
   nand U12310 ( n12491,n11777,n12493 );
   nand U12311 ( n12493,n11730,n11729 );
   nand U12312 ( n11730,n12494,n11697 );
   not U12313 ( n11697,n12495 );
   nand U12314 ( n12494,n11698,n11699 );
   nand U12315 ( n11699,n12496,n12497 );
   nand U12316 ( n12497,n12498,n10639 );
   nand U12317 ( n12498,n11663,n11679 );
   or U12318 ( n12496,n11663,n11679 );
   nor U12319 ( n11663,n12499,n11633 );
   nor U12320 ( n11633,n11636,n12500 );
   not U12321 ( n12500,n12501 );
   nand U12322 ( n11636,n12502,n11609 );
   nand U12323 ( n12502,n11608,n11607 );
   not U12324 ( n11607,n11578 );
   nor U12325 ( n11578,n12503,n11576 );
   and U12326 ( n11576,n11553,n12504 );
   nand U12327 ( n12504,n11555,n11554 );
   not U12328 ( n11555,n11552 );
   nand U12329 ( n11552,n12505,n12506 );
   nand U12330 ( n12505,n11531,n12507 );
   not U12331 ( n11531,n11529 );
   nand U12332 ( n12510,n10781,n10782,n11479 );
   nand U12333 ( n10781,n10780,n12512 );
   nand U12334 ( n12512,n12338,n12513 );
   nand U12335 ( n12509,n12350,n10780 );
   nand U12336 ( n12508,n11445,p2_reg2_reg_30_ );
   or U12337 ( n12511,n10769,n11445 );
   nand U12338 ( n10769,n12357,n10570 );
   nand U12339 ( n12357,n12517,n12518 );
   nand U12340 ( n12518,n10808,n12519 );
   nand U12341 ( n12517,n12521,n12522 );
   nand U12342 ( n12516,n11479,n10774 );
   xor U12343 ( n10774,n10782,n10771 );
   nand U12344 ( n10782,n12523,n12513,n12338 );
   nor U12345 ( n12338,n12336,n12300,n12262 );
   not U12346 ( n12262,n12299 );
   nor U12347 ( n12299,n12264,n12235,n12208 );
   not U12348 ( n12208,n12234 );
   nor U12349 ( n12234,n12190,n10853,n12151 );
   not U12350 ( n12151,n12189 );
   nor U12351 ( n12189,n12153,n12114,n12069 );
   not U12352 ( n12069,n12113 );
   nor U12353 ( n12113,n12071,n12044,n12019 );
   not U12354 ( n12019,n12045 );
   nor U12355 ( n12045,n12021,n11986,n11957 );
   not U12356 ( n11957,n11987 );
   nor U12357 ( n11987,n11913,n11959,n11880 );
   not U12358 ( n11880,n11914 );
   nor U12359 ( n11914,n12524,n11883,n11810 );
   not U12360 ( n11810,n11837 );
   nor U12361 ( n11837,n11812,n11782,n11734 );
   not U12362 ( n11734,n11783 );
   nor U12363 ( n11783,n11737,n11018,n11677 );
   not U12364 ( n11677,n11738 );
   nor U12365 ( n11738,n11679,n11042,n11612 );
   not U12366 ( n11612,n11644 );
   nor U12367 ( n11644,n11057,n11582,n11557 );
   not U12368 ( n11557,n11581 );
   nor U12369 ( n11581,n11090,n11080,n11509 );
   not U12370 ( n11509,n11560 );
   nor U12371 ( n11560,n11125,n11104,n11114 );
   nor U12372 ( n11479,n12525,n11445,n10790 );
   nand U12373 ( n12515,n12350,n10771 );
   not U12374 ( n12350,n11459 );
   nand U12375 ( n12514,n11445,p2_reg2_reg_31_ );
   nand U12376 ( n12528,n10763,n11135,n12529,n12530 );
   nor U12377 ( n12530,n10764,n11134 );
   not U12378 ( n11135,n12531 );
   nor U12379 ( n12537,n12538,n12539,n12540 );
   nor U12380 ( n12540,n12541,n12542,n12543 );
   nor U12381 ( n12542,n12544,n12017 );
   xor U12382 ( n12541,n12043,n11130 );
   not U12383 ( n12043,p2_reg2_reg_19_ );
   nor U12384 ( n12539,n12545,n12546,n12544 );
   nor U12385 ( n12544,n12547,n12548 );
   nor U12386 ( n12546,p2_reg2_reg_18_,n12543 );
   nor U12387 ( n12543,n12549,n12550 );
   not U12388 ( n12549,n12548 );
   xor U12389 ( n12545,n11130,p2_reg2_reg_19_ );
   nor U12390 ( n12536,n12551,n12552,n12553 );
   nor U12391 ( n12553,n12554,n12555,n12556 );
   nor U12392 ( n12555,n12557,n12558 );
   xor U12393 ( n12554,p2_reg1_reg_19_,n12525 );
   nor U12394 ( n12552,n12559,n12560,n12557 );
   nor U12395 ( n12557,n12547,n12561 );
   nor U12396 ( n12560,p2_reg1_reg_18_,n12556 );
   nor U12397 ( n12556,n12562,n12550 );
   not U12398 ( n12562,n12561 );
   xor U12399 ( n12559,n11130,p2_reg1_reg_19_ );
   nor U12400 ( n12535,n11130,n12563 );
   nand U12401 ( n12533,n12564,p2_addr_reg_19_ );
   nand U12402 ( n12532,p2_reg3_reg_19_,p2_u3152 );
   nand U12403 ( n12569,n12570,n12563,n12571 );
   nand U12404 ( n12571,n12572,n12573 );
   xor U12405 ( n12573,n12017,n12548 );
   not U12406 ( n12017,p2_reg2_reg_18_ );
   nand U12407 ( n12570,n12574,n12575 );
   xor U12408 ( n12575,n12558,n12561 );
   not U12409 ( n12558,p2_reg1_reg_18_ );
   not U12410 ( n12547,n12550 );
   nand U12411 ( n12567,n12576,n12550 );
   nand U12412 ( n12576,n12577,n12578 );
   nand U12413 ( n12578,n12579,n12574 );
   xor U12414 ( n12579,n12561,p2_reg1_reg_18_ );
   nand U12415 ( n12561,n12580,n12581,n12582 );
   or U12416 ( n12582,n12583,n12584 );
   nand U12417 ( n12581,p2_reg1_reg_17_,n12585 );
   or U12418 ( n12585,n12586,n12587 );
   nand U12419 ( n12580,n12587,n12586 );
   nand U12420 ( n12577,n12588,n12572 );
   xor U12421 ( n12588,n12548,p2_reg2_reg_18_ );
   nand U12422 ( n12548,n12589,n12590,n12591 );
   or U12423 ( n12591,n12592,n12593 );
   nand U12424 ( n12590,p2_reg2_reg_17_,n12594 );
   or U12425 ( n12594,n12586,n12595 );
   nand U12426 ( n12589,n12595,n12586 );
   nand U12427 ( n12566,p2_addr_reg_18_,n12564 );
   nand U12428 ( n12565,p2_reg3_reg_18_,p2_u3152 );
   nor U12429 ( n12601,n12538,n12602,n12603 );
   nor U12430 ( n12603,n12604,n12595,n12605 );
   nor U12431 ( n12605,n12606,n12592 );
   nor U12432 ( n12606,p2_reg2_reg_16_,n12607 );
   xor U12433 ( n12604,n12586,p2_reg2_reg_17_ );
   nor U12434 ( n12602,n12593,n12608,n12609 );
   nor U12435 ( n12609,n11985,n12610 );
   nor U12436 ( n12608,n12595,n12611 );
   nor U12437 ( n12595,n12612,n11955 );
   nand U12438 ( n12593,n12613,n12614 );
   nand U12439 ( n12614,n12612,n11955 );
   nand U12440 ( n12613,n12610,n11985 );
   not U12441 ( n11985,p2_reg2_reg_17_ );
   nor U12442 ( n12600,n12551,n12615,n12616 );
   nor U12443 ( n12616,n12617,n12587,n12618 );
   nor U12444 ( n12618,n12619,n12583 );
   nor U12445 ( n12619,p2_reg1_reg_16_,n12607 );
   xor U12446 ( n12617,n12586,p2_reg1_reg_17_ );
   not U12447 ( n12586,n12610 );
   nor U12448 ( n12615,n12584,n12620,n12621 );
   nor U12449 ( n12621,n12622,n12610 );
   nor U12450 ( n12620,n12587,n12623 );
   nor U12451 ( n12587,n12612,n12624 );
   nand U12452 ( n12584,n12625,n12626 );
   nand U12453 ( n12626,n12612,n12624 );
   nand U12454 ( n12625,n12610,n12622 );
   not U12455 ( n12622,p2_reg1_reg_17_ );
   nor U12456 ( n12599,n12610,n12563 );
   nand U12457 ( n12597,p2_addr_reg_17_,n12564 );
   nand U12458 ( n12596,p2_reg3_reg_17_,p2_u3152 );
   nand U12459 ( n12631,n12632,n12633 );
   nand U12460 ( n12633,n12574,n12634 );
   xor U12461 ( n12634,n12623,p2_reg1_reg_16_ );
   nand U12462 ( n12632,n12572,n12635 );
   xor U12463 ( n12635,n12611,p2_reg2_reg_16_ );
   nand U12464 ( n12629,n12607,n12636 );
   nand U12465 ( n12636,n12637,n12563,n12638 );
   nand U12466 ( n12638,n12639,n12572 );
   xor U12467 ( n12639,n11955,n12611 );
   not U12468 ( n12611,n12592 );
   nand U12469 ( n12592,n12640,n12641 );
   nand U12470 ( n12641,n12642,n11912 );
   or U12471 ( n12642,n12643,n12644 );
   nand U12472 ( n12640,n12643,n12644 );
   not U12473 ( n11955,p2_reg2_reg_16_ );
   nand U12474 ( n12637,n12645,n12574 );
   xor U12475 ( n12645,n12624,n12623 );
   not U12476 ( n12623,n12583 );
   nand U12477 ( n12583,n12646,n12647 );
   nand U12478 ( n12647,n12648,n12649 );
   or U12479 ( n12648,n12644,n12650 );
   nand U12480 ( n12646,n12650,n12644 );
   not U12481 ( n12624,p2_reg1_reg_16_ );
   not U12482 ( n12607,n12612 );
   nand U12483 ( n12628,p2_addr_reg_16_,n12564 );
   nand U12484 ( n12627,p2_reg3_reg_16_,p2_u3152 );
   nand U12485 ( n12656,n12657,n12563,n12658 );
   nand U12486 ( n12658,n12659,n12572 );
   xor U12487 ( n12659,p2_reg2_reg_15_,n12643 );
   nand U12488 ( n12657,n12660,n12574 );
   xor U12489 ( n12660,p2_reg1_reg_15_,n12650 );
   not U12490 ( n12655,n12644 );
   nand U12491 ( n12653,n12661,n12644 );
   nand U12492 ( n12661,n12662,n12663 );
   nand U12493 ( n12663,n12574,n12664 );
   xor U12494 ( n12664,n12650,n12649 );
   not U12495 ( n12649,p2_reg1_reg_15_ );
   nand U12496 ( n12650,n12665,n12666 );
   nand U12497 ( n12666,n12667,n12668 );
   nand U12498 ( n12667,n12669,n12670 );
   or U12499 ( n12665,n12670,n12669 );
   nand U12500 ( n12662,n12572,n12671 );
   xor U12501 ( n12671,n12643,n11912 );
   not U12502 ( n11912,p2_reg2_reg_15_ );
   nand U12503 ( n12643,n12672,n12673 );
   nand U12504 ( n12673,n12674,n11879 );
   nand U12505 ( n12674,n12675,n12670 );
   or U12506 ( n12672,n12670,n12675 );
   nand U12507 ( n12652,p2_addr_reg_15_,n12564 );
   nand U12508 ( n12651,p2_reg3_reg_15_,p2_u3152 );
   nand U12509 ( n12679,n12680,n12681 );
   nand U12510 ( n12681,n12682,n12683 );
   nand U12511 ( n12683,n12574,n12684 );
   xor U12512 ( n12684,n12669,p2_reg1_reg_14_ );
   nand U12513 ( n12682,n12572,n12685 );
   xor U12514 ( n12685,n12675,p2_reg2_reg_14_ );
   nand U12515 ( n12678,n12670,n12686 );
   nand U12516 ( n12686,n12687,n12563,n12688 );
   nand U12517 ( n12688,n12689,n12572 );
   xor U12518 ( n12689,n11879,n12675 );
   nor U12519 ( n12675,n12690,n12691 );
   and U12520 ( n12690,n12692,n12693,n12694 );
   nand U12521 ( n12694,n12695,p2_reg2_reg_13_ );
   not U12522 ( n11879,p2_reg2_reg_14_ );
   nand U12523 ( n12687,n12696,n12574 );
   xor U12524 ( n12696,n12668,n12669 );
   nor U12525 ( n12669,n12697,n12698 );
   and U12526 ( n12697,n12699,n12700,n12701 );
   nand U12527 ( n12701,n12695,p2_reg1_reg_13_ );
   not U12528 ( n12668,p2_reg1_reg_14_ );
   nand U12529 ( n12677,p2_addr_reg_14_,n12564 );
   nand U12530 ( n12676,p2_reg3_reg_14_,p2_u3152 );
   nor U12531 ( n12707,n12538,n12708,n12709 );
   nor U12532 ( n12709,n12710,n12711,n12712 );
   nor U12533 ( n12712,n12713,n12714 );
   xor U12534 ( n12710,n12695,p2_reg2_reg_13_ );
   nor U12535 ( n12708,n12691,n12714,n12715,n12716 );
   nor U12536 ( n12716,n11836,n12717 );
   not U12537 ( n11836,p2_reg2_reg_13_ );
   nor U12538 ( n12715,n12711,n12718 );
   nor U12539 ( n12691,p2_reg2_reg_13_,n12695 );
   nor U12540 ( n12706,n12551,n12719,n12720 );
   nor U12541 ( n12720,n12721,n12722,n12723 );
   nor U12542 ( n12723,n12724,n12725 );
   xor U12543 ( n12721,n12695,p2_reg1_reg_13_ );
   nor U12544 ( n12719,n12698,n12725,n12726,n12727 );
   and U12545 ( n12727,p2_reg1_reg_13_,n12695 );
   nor U12546 ( n12726,n12722,n12728 );
   not U12547 ( n12722,n12700 );
   nor U12548 ( n12698,p2_reg1_reg_13_,n12695 );
   nor U12549 ( n12705,n12717,n12563 );
   nand U12550 ( n12703,p2_addr_reg_13_,n12564 );
   nand U12551 ( n12702,p2_reg3_reg_13_,p2_u3152 );
   nor U12552 ( n12732,n12733,n12734 );
   nor U12553 ( n12733,n12735,n12736 );
   nand U12554 ( n12731,n12737,n12738 );
   nand U12555 ( n12738,n12739,n12563,n12740 );
   nand U12556 ( n12740,p2_reg1_reg_12_,n12728,n12574 );
   nand U12557 ( n12739,p2_reg2_reg_12_,n12718,n12572 );
   nand U12558 ( n12730,n12741,n12699,n12574 );
   nand U12559 ( n12699,n12742,n12728 );
   nand U12560 ( n12741,n12724,n12743 );
   nand U12561 ( n12743,n12700,n12742 );
   not U12562 ( n12742,n12725 );
   nor U12563 ( n12725,n12737,p2_reg1_reg_12_ );
   nand U12564 ( n12700,n12737,p2_reg1_reg_12_ );
   not U12565 ( n12724,n12728 );
   nand U12566 ( n12728,n12744,n12745 );
   nand U12567 ( n12745,n12746,n12747 );
   nand U12568 ( n12747,n12748,n12749 );
   nand U12569 ( n12744,n12750,p2_reg1_reg_11_ );
   nand U12570 ( n12729,n12751,n12692,n12572 );
   nand U12571 ( n12692,n12752,n12718 );
   nand U12572 ( n12751,n12713,n12753 );
   nand U12573 ( n12753,n12693,n12752 );
   not U12574 ( n12752,n12714 );
   nor U12575 ( n12714,n12737,p2_reg2_reg_12_ );
   not U12576 ( n12737,n12754 );
   not U12577 ( n12693,n12711 );
   nor U12578 ( n12711,n12754,n11809 );
   not U12579 ( n11809,p2_reg2_reg_12_ );
   not U12580 ( n12713,n12718 );
   nand U12581 ( n12718,n12755,n12756 );
   nand U12582 ( n12756,n12757,n12758 );
   nand U12583 ( n12758,n11781,n12749 );
   nand U12584 ( n12755,n12750,p2_reg2_reg_11_ );
   nand U12585 ( n12763,n12764,n12563,n12765 );
   nand U12586 ( n12765,n12766,n12572 );
   xor U12587 ( n12766,n11781,n12757 );
   not U12588 ( n11781,p2_reg2_reg_11_ );
   nand U12589 ( n12764,n12767,n12574 );
   xor U12590 ( n12767,n12748,n12746 );
   not U12591 ( n12748,p2_reg1_reg_11_ );
   not U12592 ( n12750,n12749 );
   nand U12593 ( n12761,n12768,n12749 );
   nand U12594 ( n12768,n12769,n12770 );
   nand U12595 ( n12770,n12574,n12771 );
   xor U12596 ( n12771,n12746,p2_reg1_reg_11_ );
   nor U12597 ( n12746,n12772,n12773 );
   and U12598 ( n12772,n12774,n12775,n12776 );
   nand U12599 ( n12776,n12777,p2_reg1_reg_10_ );
   nand U12600 ( n12774,n12778,n12779 );
   nand U12601 ( n12769,n12572,n12780 );
   xor U12602 ( n12780,n12757,p2_reg2_reg_11_ );
   nor U12603 ( n12757,n12781,n12782 );
   and U12604 ( n12781,n12783,n12784,n12785 );
   nand U12605 ( n12785,n12777,p2_reg2_reg_10_ );
   nand U12606 ( n12783,n12786,n12787 );
   nand U12607 ( n12760,p2_addr_reg_11_,n12564 );
   nand U12608 ( n12759,p2_reg3_reg_11_,p2_u3152 );
   nor U12609 ( n12793,n12538,n12794,n12795 );
   nor U12610 ( n12795,n12796,n12797,n12798 );
   nor U12611 ( n12798,n12799,n12800 );
   xor U12612 ( n12796,n12777,p2_reg2_reg_10_ );
   nor U12613 ( n12794,n12782,n12800,n12801,n12802 );
   nor U12614 ( n12802,n11733,n12803 );
   not U12615 ( n11733,p2_reg2_reg_10_ );
   nor U12616 ( n12801,n12797,n12786 );
   nor U12617 ( n12782,n12777,p2_reg2_reg_10_ );
   nor U12618 ( n12792,n12551,n12804,n12805 );
   nor U12619 ( n12805,n12806,n12807,n12808 );
   nor U12620 ( n12808,n12809,n12810 );
   xor U12621 ( n12806,n12777,p2_reg1_reg_10_ );
   nor U12622 ( n12804,n12773,n12810,n12811,n12812 );
   and U12623 ( n12812,p2_reg1_reg_10_,n12777 );
   nor U12624 ( n12811,n12807,n12778 );
   not U12625 ( n12807,n12775 );
   nor U12626 ( n12773,n12777,p2_reg1_reg_10_ );
   nor U12627 ( n12791,n12803,n12563 );
   nand U12628 ( n12789,p2_addr_reg_10_,n12564 );
   nand U12629 ( n12788,p2_reg3_reg_10_,p2_u3152 );
   nor U12630 ( n12816,n12817,n12818 );
   nor U12631 ( n12817,n12735,n12819 );
   nand U12632 ( n12815,n12820,n12821 );
   nand U12633 ( n12821,n12822,n12563,n12823 );
   nand U12634 ( n12823,p2_reg1_reg_9_,n12778,n12574 );
   nand U12635 ( n12822,p2_reg2_reg_9_,n12786,n12572 );
   nand U12636 ( n12814,n12824,n12825,n12574 );
   nand U12637 ( n12825,n12810,n12809 );
   nand U12638 ( n12824,n12826,n12779 );
   not U12639 ( n12779,n12810 );
   nor U12640 ( n12810,p2_reg1_reg_9_,n12820 );
   nand U12641 ( n12826,n12809,n12775 );
   nand U12642 ( n12775,n12820,p2_reg1_reg_9_ );
   not U12643 ( n12809,n12778 );
   nand U12644 ( n12778,n12827,n12828 );
   or U12645 ( n12827,n12829,n12830 );
   nand U12646 ( n12813,n12831,n12832,n12572 );
   nand U12647 ( n12832,n12800,n12799 );
   nand U12648 ( n12831,n12833,n12787 );
   not U12649 ( n12787,n12800 );
   nor U12650 ( n12800,p2_reg2_reg_9_,n12820 );
   not U12651 ( n12820,n12834 );
   nand U12652 ( n12833,n12799,n12784 );
   not U12653 ( n12784,n12797 );
   nor U12654 ( n12797,n12834,n11701 );
   not U12655 ( n11701,p2_reg2_reg_9_ );
   not U12656 ( n12799,n12786 );
   nand U12657 ( n12786,n12835,n12836 );
   or U12658 ( n12835,n12837,n12838 );
   nor U12659 ( n12844,n12538,n12845 );
   xor U12660 ( n12845,n12838,n12846 );
   nor U12661 ( n12846,n12847,n12837 );
   nor U12662 ( n12837,n12848,p2_reg2_reg_8_ );
   not U12663 ( n12847,n12836 );
   nand U12664 ( n12836,n12848,p2_reg2_reg_8_ );
   and U12665 ( n12838,n12849,n12850 );
   nand U12666 ( n12850,p2_reg2_reg_7_,n12851 );
   nand U12667 ( n12851,n12852,n12853 );
   nand U12668 ( n12849,n12854,n12855 );
   nor U12669 ( n12843,n12551,n12856 );
   xor U12670 ( n12856,n12830,n12857 );
   nor U12671 ( n12857,n12858,n12829 );
   nor U12672 ( n12829,n12848,p2_reg1_reg_8_ );
   not U12673 ( n12858,n12828 );
   nand U12674 ( n12828,n12848,p2_reg1_reg_8_ );
   not U12675 ( n12848,n12859 );
   and U12676 ( n12830,n12860,n12861 );
   nand U12677 ( n12861,p2_reg1_reg_7_,n12862 );
   nand U12678 ( n12862,n12863,n12853 );
   nand U12679 ( n12860,n12854,n12864 );
   nor U12680 ( n12842,n12859,n12563 );
   nand U12681 ( n12840,p2_addr_reg_8_,n12564 );
   nand U12682 ( n12839,p2_reg3_reg_8_,p2_u3152 );
   nor U12683 ( n12868,n12869,n12870 );
   nor U12684 ( n12869,n12735,n12871 );
   nand U12685 ( n12867,n12854,n12872 );
   nand U12686 ( n12872,n12873,n12563,n12874 );
   nand U12687 ( n12874,n12875,n12876,n12574 );
   not U12688 ( n12876,p2_reg1_reg_7_ );
   nand U12689 ( n12873,n12877,n11637,n12572 );
   not U12690 ( n11637,p2_reg2_reg_7_ );
   nand U12691 ( n12866,n12878,n12875,n12574 );
   nand U12692 ( n12875,n12879,n12880,n12881 );
   xor U12693 ( n12881,n12854,p2_reg1_reg_7_ );
   nand U12694 ( n12879,n12882,n12883 );
   nand U12695 ( n12878,n12863,n12884 );
   nand U12696 ( n12884,p2_reg1_reg_7_,n12853 );
   not U12697 ( n12863,n12864 );
   nand U12698 ( n12864,n12883,n12885 );
   nand U12699 ( n12865,n12886,n12877,n12572 );
   nand U12700 ( n12877,n12887,n12888,n12889 );
   xor U12701 ( n12889,n12854,p2_reg2_reg_7_ );
   not U12702 ( n12854,n12853 );
   nand U12703 ( n12887,n12890,n12891 );
   nand U12704 ( n12886,n12852,n12892 );
   nand U12705 ( n12892,p2_reg2_reg_7_,n12853 );
   not U12706 ( n12852,n12855 );
   nand U12707 ( n12855,n12891,n12893 );
   nor U12708 ( n12897,n12898,n12899 );
   nor U12709 ( n12898,n12735,n12900 );
   nand U12710 ( n12896,n12901,n12902 );
   nand U12711 ( n12902,n12903,n12563,n12904 );
   nand U12712 ( n12904,p2_reg1_reg_6_,n12905,n12574 );
   nand U12713 ( n12903,p2_reg2_reg_6_,n12906,n12572 );
   nand U12714 ( n12895,n12907,n12885,n12574 );
   nand U12715 ( n12885,n12905,n12880 );
   nand U12716 ( n12907,n12882,n12908 );
   nand U12717 ( n12908,n12883,n12880 );
   or U12718 ( n12880,n12901,p2_reg1_reg_6_ );
   nand U12719 ( n12883,n12901,p2_reg1_reg_6_ );
   not U12720 ( n12882,n12905 );
   nand U12721 ( n12905,n12909,n12910 );
   nand U12722 ( n12910,p2_reg1_reg_5_,n12911 );
   nand U12723 ( n12911,n12912,n12913 );
   nand U12724 ( n12909,n12914,n12915 );
   nand U12725 ( n12894,n12916,n12893,n12572 );
   nand U12726 ( n12893,n12906,n12888 );
   nand U12727 ( n12916,n12890,n12917 );
   nand U12728 ( n12917,n12891,n12888 );
   nand U12729 ( n12888,n12918,n11610 );
   not U12730 ( n11610,p2_reg2_reg_6_ );
   nand U12731 ( n12891,n12901,p2_reg2_reg_6_ );
   not U12732 ( n12890,n12906 );
   nand U12733 ( n12906,n12919,n12920 );
   nand U12734 ( n12920,p2_reg2_reg_5_,n12921 );
   nand U12735 ( n12921,n12922,n12913 );
   nand U12736 ( n12919,n12914,n12923 );
   nor U12737 ( n12927,n12928,n12929 );
   nor U12738 ( n12928,n12735,n12930 );
   nand U12739 ( n12926,n12914,n12931 );
   nand U12740 ( n12931,n12932,n12563,n12933 );
   nand U12741 ( n12933,n12934,n12935,n12574 );
   not U12742 ( n12935,p2_reg1_reg_5_ );
   nand U12743 ( n12932,n12936,n11580,n12572 );
   not U12744 ( n11580,p2_reg2_reg_5_ );
   nand U12745 ( n12925,n12937,n12934,n12574 );
   nand U12746 ( n12934,n12938,n12939,n12940 );
   xor U12747 ( n12940,n12914,p2_reg1_reg_5_ );
   nand U12748 ( n12938,n12941,n12942 );
   nand U12749 ( n12937,n12912,n12943 );
   nand U12750 ( n12943,p2_reg1_reg_5_,n12913 );
   not U12751 ( n12912,n12915 );
   nand U12752 ( n12915,n12942,n12944 );
   nand U12753 ( n12924,n12945,n12936,n12572 );
   nand U12754 ( n12936,n12946,n12947,n12948 );
   xor U12755 ( n12948,n12914,p2_reg2_reg_5_ );
   not U12756 ( n12914,n12913 );
   nand U12757 ( n12946,n12949,n12950 );
   nand U12758 ( n12945,n12922,n12951 );
   nand U12759 ( n12951,p2_reg2_reg_5_,n12913 );
   not U12760 ( n12922,n12923 );
   nand U12761 ( n12923,n12950,n12952 );
   nor U12762 ( n12956,n12957,n12958 );
   nor U12763 ( n12957,n12735,n12959 );
   nand U12764 ( n12955,n12960,n12961 );
   nand U12765 ( n12961,n12962,n12563,n12963 );
   nand U12766 ( n12963,p2_reg1_reg_4_,n12964,n12574 );
   nand U12767 ( n12962,p2_reg2_reg_4_,n12965,n12572 );
   nand U12768 ( n12954,n12966,n12944,n12574 );
   nand U12769 ( n12944,n12964,n12939 );
   nand U12770 ( n12966,n12941,n12967 );
   nand U12771 ( n12967,n12942,n12939 );
   or U12772 ( n12939,n12960,p2_reg1_reg_4_ );
   nand U12773 ( n12942,n12960,p2_reg1_reg_4_ );
   not U12774 ( n12941,n12964 );
   nand U12775 ( n12964,n12968,n12969 );
   nand U12776 ( n12969,n12970,n12971 );
   nand U12777 ( n12971,n12972,n12973 );
   nand U12778 ( n12970,n12974,n12975 );
   nand U12779 ( n12968,n12976,p2_reg1_reg_3_ );
   nand U12780 ( n12953,n12977,n12952,n12572 );
   nand U12781 ( n12952,n12965,n12947 );
   nand U12782 ( n12977,n12949,n12978 );
   nand U12783 ( n12978,n12950,n12947 );
   nand U12784 ( n12947,n12979,n11556 );
   not U12785 ( n11556,p2_reg2_reg_4_ );
   nand U12786 ( n12950,n12960,p2_reg2_reg_4_ );
   not U12787 ( n12960,n12979 );
   not U12788 ( n12949,n12965 );
   nand U12789 ( n12965,n12980,n12981 );
   nand U12790 ( n12981,n12982,n12983 );
   nand U12791 ( n12983,n12972,n11533 );
   nand U12792 ( n12982,n12984,n12985 );
   nand U12793 ( n12980,n12976,p2_reg2_reg_3_ );
   nand U12794 ( n12989,n12972,n12990 );
   nand U12795 ( n12990,n12991,n12992 );
   nand U12796 ( n12992,n12993,n12574 );
   xor U12797 ( n12993,n12994,n12973 );
   not U12798 ( n12973,p2_reg1_reg_3_ );
   nand U12799 ( n12991,n12995,n12572 );
   xor U12800 ( n12995,n12996,n11533 );
   not U12801 ( n11533,p2_reg2_reg_3_ );
   nand U12802 ( n12988,n12976,n12997 );
   nand U12803 ( n12997,n12998,n12563,n12999 );
   nand U12804 ( n12999,n12572,n13000 );
   xor U12805 ( n13000,p2_reg2_reg_3_,n12996 );
   and U12806 ( n12996,n12984,n12985 );
   nand U12807 ( n12985,n13001,n13002 );
   nand U12808 ( n13002,n13003,n11502 );
   and U12809 ( n12984,n13004,n13005 );
   nand U12810 ( n13005,p2_reg2_reg_2_,n13006 );
   nand U12811 ( n13006,n13003,n13007 );
   nand U12812 ( n13004,n13008,n13009 );
   nand U12813 ( n12998,n12574,n13010 );
   xor U12814 ( n13010,p2_reg1_reg_3_,n12994 );
   and U12815 ( n12994,n12974,n12975 );
   nand U12816 ( n12975,n13011,n13012 );
   nand U12817 ( n13012,n13003,n13013 );
   and U12818 ( n12974,n13014,n13015 );
   nand U12819 ( n13015,p2_reg1_reg_2_,n13016 );
   nand U12820 ( n13016,n13003,n13017 );
   nand U12821 ( n13014,n13018,n13009 );
   nand U12822 ( n12987,p2_addr_reg_3_,n12564 );
   nand U12823 ( n12986,p2_reg3_reg_3_,p2_u3152 );
   nor U12824 ( n13024,n12538,n13025,n13026 );
   nor U12825 ( n13026,n13027,n13028 );
   xor U12826 ( n13028,n11502,n13009 );
   not U12827 ( n11502,p2_reg2_reg_2_ );
   nor U12828 ( n13027,n13001,n13008 );
   nor U12829 ( n13025,n13029,n13001,n13008 );
   and U12830 ( n13001,p2_reg2_reg_0_,n13030,p2_ir_reg_0_ );
   xor U12831 ( n13029,n13009,p2_reg2_reg_2_ );
   nor U12832 ( n13023,n12551,n13031,n13032 );
   nor U12833 ( n13032,n13033,n13034 );
   xor U12834 ( n13034,n13013,n13009 );
   not U12835 ( n13013,p2_reg1_reg_2_ );
   nor U12836 ( n13033,n13011,n13018 );
   nor U12837 ( n13031,n13035,n13011,n13018 );
   and U12838 ( n13011,p2_reg1_reg_0_,n13036,p2_ir_reg_0_ );
   xor U12839 ( n13035,n13009,p2_reg1_reg_2_ );
   not U12840 ( n13009,n13003 );
   nor U12841 ( n13022,n13003,n12563 );
   nand U12842 ( n13020,p2_addr_reg_2_,n12564 );
   nand U12843 ( n13019,p2_reg3_reg_2_,p2_u3152 );
   nor U12844 ( n13042,n13043,n12538 );
   xor U12845 ( n13043,n13044,n13045 );
   nand U12846 ( n13045,n13007,n13030 );
   nand U12847 ( n13030,n13046,n11478 );
   not U12848 ( n13007,n13008 );
   nor U12849 ( n13008,n13046,n11478 );
   not U12850 ( n11478,p2_reg2_reg_1_ );
   nor U12851 ( n13044,n11454,n13047 );
   nor U12852 ( n13041,n13048,n12551 );
   xor U12853 ( n13048,n13049,n13050 );
   nand U12854 ( n13050,n13017,n13036 );
   nand U12855 ( n13036,n13046,n13051 );
   not U12856 ( n13017,n13018 );
   nor U12857 ( n13018,n13046,n13051 );
   not U12858 ( n13051,p2_reg1_reg_1_ );
   nor U12859 ( n13049,n13052,n13047 );
   nor U12860 ( n13040,n13046,n12563 );
   nand U12861 ( n13038,p2_addr_reg_1_,n12564 );
   nand U12862 ( n13037,p2_reg3_reg_1_,p2_u3152 );
   nand U12863 ( n13057,n13058,n12563,n13059 );
   nand U12864 ( n13059,n12572,n11454 );
   not U12865 ( n11454,p2_reg2_reg_0_ );
   nand U12866 ( n13058,n12574,n13052 );
   not U12867 ( n13052,p2_reg1_reg_0_ );
   nand U12868 ( n13055,n13061,n13047 );
   nand U12869 ( n13061,n13062,n13063 );
   nand U12870 ( n13063,n12574,p2_reg1_reg_0_ );
   nand U12871 ( n12551,n13064,n13065 );
   nand U12872 ( n13064,n13066,n13067 );
   nand U12873 ( n13066,n12520,n19378 );
   nand U12874 ( n13062,n12572,p2_reg2_reg_0_ );
   nand U12875 ( n12538,n12520,n13060,n13068 );
   nand U12876 ( n13060,n10569,n13067 );
   nand U12877 ( n13067,n13069,n12735 );
   nand U12878 ( n13069,n10764,n13070 );
   nand U12879 ( n13070,n13071,p2_state_reg );
   nand U12880 ( n13054,p2_addr_reg_0_,n12564 );
   not U12881 ( n12564,n12735 );
   nand U12882 ( n12735,n13073,n13072,n13074 );
   nand U12883 ( n13073,n13075,n12366 );
   nand U12884 ( n13053,p2_reg3_reg_0_,p2_u3152 );
   nor U12885 ( n13077,n13078,n13079 );
   nor U12886 ( n13078,p2_u3152,n13080 );
   nor U12887 ( n13076,n13081,n13082,n13079,n13083 );
   nor U12888 ( n13083,n11629,n13084,n13085 );
   nor U12889 ( n13085,n11142,n13086,n13087,n13088 );
   nor U12890 ( n13088,n13089,n13090,n13091 );
   nor U12891 ( n13091,n12446,n13092 );
   nor U12892 ( n13092,n13093,n13094,n13095 );
   nor U12893 ( n13093,n13096,n13097 );
   nor U12894 ( n13096,n13098,n13099 );
   nor U12895 ( n13099,n13100,n13101 );
   nor U12896 ( n13101,n10850,n12235 );
   nor U12897 ( n13100,n13102,n13103 );
   nor U12898 ( n13103,n13104,n13105 );
   nor U12899 ( n13105,n12226,n10853 );
   nor U12900 ( n13104,n13106,n13107 );
   nor U12901 ( n13107,n13108,n13109 );
   nor U12902 ( n13109,n13110,n12465 );
   nand U12903 ( n12465,n12146,n12460 );
   nor U12904 ( n13110,n12188,n12184,n13111,n13112 );
   nor U12905 ( n13112,n12466,n12469 );
   and U12906 ( n13111,n13113,n12467,n13114,n12470 );
   and U12907 ( n13113,n13115,n13116 );
   nand U12908 ( n13116,n13117,n13118 );
   nand U12909 ( n13118,n13119,n13120 );
   nand U12910 ( n13120,n13121,n13122 );
   nand U12911 ( n13122,n12484,n13123 );
   nand U12912 ( n13123,n13124,n11908 );
   nand U12913 ( n13124,n11876,n13125 );
   nand U12914 ( n13125,n12487,n11877,n13126 );
   nand U12915 ( n13126,n13127,n12485,n13128 );
   nand U12916 ( n13127,n13129,n13130,n13131 );
   nand U12917 ( n13129,n13132,n13133 );
   nand U12918 ( n13133,n13134,n11634,n13135 );
   nand U12919 ( n13135,n13136,n11609 );
   nand U12920 ( n13136,n11579,n13137 );
   or U12921 ( n13137,n13138,n12503 );
   not U12922 ( n11877,n11864 );
   nand U12923 ( n13115,n13139,n12472 );
   nor U12924 ( n13108,n13140,n12190 );
   nor U12925 ( n13086,n13141,n13142 );
   nor U12926 ( n13142,n13143,n13144 );
   nor U12927 ( n13144,n10780,n13145 );
   nor U12928 ( n13143,n13090,n13146,n10791 );
   and U12929 ( n13090,n10780,n13145 );
   nor U12930 ( n13084,n11131,n13147 );
   and U12931 ( n13079,p2_b_reg,n13148 );
   nand U12932 ( n13148,n13072,p2_state_reg,n13149,n13150 );
   nand U12933 ( n13150,n13071,n11131 );
   nand U12934 ( n13149,n13080,n13151 );
   nand U12935 ( n13151,n13068,n12520,n13152,n13153 );
   nor U12936 ( n13082,n13154,n13147 );
   nand U12937 ( n13147,n13155,n13156,n13157 );
   nand U12938 ( n13157,n13158,n12523,n13159 );
   nand U12939 ( n13159,n13160,n13145,n13161 );
   nand U12940 ( n13161,n11141,n10573 );
   nand U12941 ( n13145,n10573,n10570 );
   nand U12942 ( n13160,n13162,n13163 );
   not U12943 ( n13156,n13087 );
   nand U12944 ( n13155,n13164,n13165,n13163,n10573 );
   nand U12945 ( n13163,n13166,n12443,n13167 );
   nand U12946 ( n13167,n12513,n10576 );
   not U12947 ( n12443,n12446 );
   nand U12948 ( n13166,n12449,n12444,n13168 );
   nand U12949 ( n13168,n13169,n13170 );
   nand U12950 ( n13170,n12451,n12258,n13171 );
   nand U12951 ( n13171,n12457,n13172,n12453 );
   nand U12952 ( n12453,n10841,n10588 );
   nand U12953 ( n13172,n12454,n12460,n13173 );
   nand U12954 ( n13173,n12462,n13174 );
   nand U12955 ( n13174,n13114,n12146,n13175 );
   nand U12956 ( n13175,n12469,n12110,n13176 );
   nand U12957 ( n13176,n12467,n12470,n13177 );
   nand U12958 ( n13177,n13117,n13178 );
   nand U12959 ( n13178,n13179,n12473,n13119 );
   nand U12960 ( n13119,n11986,n12010 );
   not U12961 ( n12473,n13139 );
   nor U12962 ( n13139,n10918,n10609 );
   nand U12963 ( n13179,n13180,n13181,n13121 );
   and U12964 ( n13121,n11954,n13182 );
   nand U12965 ( n13182,n10929,n10612 );
   nand U12966 ( n11954,n10941,n10615 );
   nand U12967 ( n13181,n12484,n13183,n11876,n12485 );
   nand U12968 ( n12485,n11872,n12524 );
   nand U12969 ( n11876,n13184,n11883 );
   nand U12970 ( n13183,n13185,n12487 );
   nand U12971 ( n12487,n10973,n10624 );
   nand U12972 ( n13185,n13128,n13186 );
   nand U12973 ( n13186,n13130,n13187,n13131 );
   and U12974 ( n13131,n13188,n12490,n11777 );
   and U12975 ( n11777,n11728,n13189 );
   nand U12976 ( n13189,n10995,n10630 );
   not U12977 ( n11728,n11779 );
   nor U12978 ( n11779,n11737,n11017 );
   nand U12979 ( n13188,n11031,n10639,n11729,n11698 );
   nand U12980 ( n13187,n13132,n13190 );
   nand U12981 ( n13190,n11634,n13191 );
   nand U12982 ( n13191,n13192,n11609,n13193 );
   nand U12983 ( n13193,n12503,n13134 );
   nor U12984 ( n12503,n11068,n10648 );
   nand U12985 ( n11609,n13194,n11057 );
   nand U12986 ( n13192,n13138,n11608 );
   and U12987 ( n11608,n13134,n11579 );
   not U12988 ( n11579,n11602 );
   nor U12989 ( n11602,n11582,n11077 );
   nand U12990 ( n13134,n11596,n10645 );
   and U12991 ( n13138,n11553,n13195 );
   nand U12992 ( n13195,n13196,n11554 );
   nand U12993 ( n11554,n11080,n11089 );
   nand U12994 ( n13196,n12507,n13197 );
   nand U12995 ( n13197,n11529,n12506 );
   nand U12996 ( n12506,n11101,n11090 );
   nand U12997 ( n11529,n11501,n11500 );
   nand U12998 ( n11500,n11490,n10657 );
   nand U12999 ( n11501,n11498,n11506 );
   nand U13000 ( n11506,n11104,n11113 );
   and U13001 ( n11498,n13198,n13199 );
   nand U13002 ( n13199,n13200,n11114 );
   nand U13003 ( n13200,n10660,n11450 );
   or U13004 ( n13198,n11450,n10660 );
   nand U13005 ( n12507,n11520,n10654 );
   nand U13006 ( n11553,n11546,n10651 );
   not U13007 ( n11634,n12499 );
   nor U13008 ( n12499,n11042,n11054 );
   and U13009 ( n13132,n13201,n11729,n12501,n11698 );
   nand U13010 ( n11698,n11018,n13202 );
   nand U13011 ( n12501,n11042,n11054 );
   nand U13012 ( n13201,n11679,n11041 );
   nand U13013 ( n13130,n12495,n11729 );
   not U13014 ( n11729,n11776 );
   nor U13015 ( n11776,n10633,n11007 );
   nor U13016 ( n12495,n11018,n13202 );
   and U13017 ( n13128,n12488,n13203 );
   nand U13018 ( n13203,n12492,n12490 );
   nand U13019 ( n12490,n10985,n10627 );
   nor U13020 ( n12492,n10630,n10995 );
   nand U13021 ( n12488,n11832,n11812 );
   and U13022 ( n12484,n11953,n13204 );
   nand U13023 ( n13180,n12483,n11953 );
   nand U13024 ( n11953,n11959,n11979 );
   nand U13025 ( n12483,n11908,n13205 );
   nand U13026 ( n13205,n11864,n13204 );
   not U13027 ( n13204,n11940 );
   nor U13028 ( n11940,n10951,n10618 );
   nor U13029 ( n11864,n11883,n13184 );
   not U13030 ( n13184,n10621 );
   nand U13031 ( n11908,n10951,n10618 );
   and U13032 ( n13117,n12472,n12475 );
   nand U13033 ( n12475,n10918,n10609 );
   nand U13034 ( n12472,n10606,n10907 );
   nand U13035 ( n12470,n12044,n12062 );
   nand U13036 ( n12467,n12071,n12106 );
   not U13037 ( n12110,n12188 );
   nor U13038 ( n12188,n12114,n12139 );
   nand U13039 ( n12469,n10897,n10603 );
   nand U13040 ( n12146,n12170,n12153 );
   not U13041 ( n13114,n12466 );
   nor U13042 ( n12466,n10600,n10885 );
   and U13043 ( n12462,n12145,n13206 );
   nand U13044 ( n13206,n10863,n10594 );
   not U13045 ( n12145,n12184 );
   nor U13046 ( n12184,n12153,n12170 );
   nand U13047 ( n12460,n13140,n12190 );
   not U13048 ( n12454,n13106 );
   nor U13049 ( n13106,n10591,n12199 );
   nand U13050 ( n12457,n12199,n10591 );
   not U13051 ( n12258,n13098 );
   nor U13052 ( n13098,n10829,n10585 );
   not U13053 ( n12451,n13102 );
   nor U13054 ( n13102,n10588,n10841 );
   not U13055 ( n13169,n13097 );
   nand U13056 ( n13097,n12257,n12447 );
   not U13057 ( n12444,n13094 );
   not U13058 ( n12449,n13095 );
   nor U13059 ( n13095,n10582,n10817 );
   nand U13060 ( n13165,n13207,n13153 );
   not U13061 ( n13164,n13089 );
   nand U13062 ( n13089,n13158,n13162 );
   nand U13063 ( n13162,n10791,n13146 );
   not U13064 ( n13158,n13141 );
   nor U13065 ( n13154,n13208,n11528 );
   not U13066 ( n11528,n11630 );
   nor U13067 ( n13208,n12525,n10790 );
   nand U13068 ( n13081,n13210,n13211,n13212,n13213 );
   or U13069 ( n13213,n13214,n12348,n13215 );
   nand U13070 ( n13212,n13209,n11141,n13215 );
   and U13071 ( n13215,n13216,n13217,n13218,n13219 );
   nor U13072 ( n13219,n13220,n13221,n13222,n13223 );
   nand U13073 ( n13223,n11532,n11867,n13224,n11584 );
   xor U13074 ( n11584,n11582,n11077 );
   xor U13075 ( n13224,n12523,n10573 );
   xor U13076 ( n11867,n10621,n10963 );
   not U13077 ( n11532,n11524 );
   xor U13078 ( n11524,n11520,n11101 );
   or U13079 ( n13222,n11635,n11909,n12358,n13141 );
   nor U13080 ( n13141,n10771,n13207 );
   not U13081 ( n13207,n10570 );
   not U13082 ( n12358,n12368 );
   xor U13083 ( n12368,n13146,n10791 );
   not U13084 ( n13146,n10576 );
   xor U13085 ( n11909,n10618,n11913 );
   not U13086 ( n11635,n11643 );
   xor U13087 ( n11643,n11042,n11054 );
   nand U13088 ( n13221,n11476,n11497,n13225,n11605 );
   nand U13089 ( n11605,n11642,n11639 );
   nand U13090 ( n11639,n13194,n11596 );
   not U13091 ( n11642,n11640 );
   nor U13092 ( n11640,n11596,n13194 );
   not U13093 ( n11596,n11057 );
   not U13094 ( n13225,n11551 );
   nor U13095 ( n11551,n11587,n11586 );
   nor U13096 ( n11586,n10651,n11080 );
   nor U13097 ( n11587,n11546,n11089 );
   nand U13098 ( n11497,n11537,n12427 );
   nand U13099 ( n12427,n11104,n10657 );
   nand U13100 ( n11537,n11113,n11490 );
   nand U13101 ( n11476,n12429,n13226 );
   or U13102 ( n13226,n10660,n11114 );
   nand U13103 ( n12429,n11114,n10660 );
   nand U13104 ( n13220,n11664,n11743,n11780,n11806 );
   nand U13105 ( n11806,n11844,n11846 );
   nand U13106 ( n11846,n11832,n10985 );
   not U13107 ( n11832,n10627 );
   nand U13108 ( n11844,n11812,n10627 );
   or U13109 ( n11780,n11848,n13227 );
   nor U13110 ( n13227,n10630,n11782 );
   nor U13111 ( n11848,n10995,n11802 );
   nand U13112 ( n11743,n12408,n12405 );
   nand U13113 ( n12405,n11737,n10633 );
   nand U13114 ( n12408,n11017,n11007 );
   not U13115 ( n11017,n10633 );
   nand U13116 ( n11664,n12410,n12411 );
   nand U13117 ( n12411,n11041,n11031 );
   nand U13118 ( n12410,n11679,n10639 );
   nor U13119 ( n13218,n13228,n13229,n11951,n13087 );
   nor U13120 ( n13087,n10570,n13230 );
   not U13121 ( n11951,n11939 );
   nand U13122 ( n11939,n11994,n11991 );
   nand U13123 ( n11991,n11959,n10615 );
   nand U13124 ( n11994,n11979,n10941 );
   nand U13125 ( n13229,n11453,n11700,n12332 );
   nand U13126 ( n12332,n12360,n12362 );
   nand U13127 ( n11700,n11742,n11745 );
   nand U13128 ( n11745,n13202,n11691 );
   not U13129 ( n13202,n10636 );
   nand U13130 ( n11742,n11018,n10636 );
   nand U13131 ( n11453,n13231,n11481 );
   nand U13132 ( n11481,n11125,n10663 );
   nand U13133 ( n13231,n11452,n13232 );
   nand U13134 ( n13228,n12206,n12232,n12266,n12291 );
   nand U13135 ( n12291,n12434,n12371 );
   nand U13136 ( n12371,n12324,n10817 );
   nand U13137 ( n12266,n12437,n12303 );
   not U13138 ( n12303,n12436 );
   nand U13139 ( n12437,n12288,n10829 );
   nand U13140 ( n12232,n12267,n12269 );
   nand U13141 ( n12269,n10850,n10841 );
   nand U13142 ( n12267,n12235,n10588 );
   nand U13143 ( n12206,n12275,n12273 );
   nand U13144 ( n12273,n12226,n12199 );
   nand U13145 ( n12275,n10853,n10591 );
   nor U13146 ( n13217,n12185,n12148,n12111,n13233 );
   not U13147 ( n13233,n12065 );
   nand U13148 ( n12065,n12078,n12387 );
   nand U13149 ( n12387,n12106,n10897 );
   nand U13150 ( n12078,n12071,n10603 );
   not U13151 ( n12111,n12101 );
   nand U13152 ( n12101,n12380,n12382 );
   nand U13153 ( n12382,n12139,n10885 );
   nand U13154 ( n12380,n12114,n10600 );
   and U13155 ( n12148,n12378,n12376 );
   nand U13156 ( n12376,n12170,n10875 );
   not U13157 ( n12170,n10597 );
   nand U13158 ( n12378,n12153,n10597 );
   not U13159 ( n12185,n12180 );
   nand U13160 ( n12180,n12375,n12373 );
   nand U13161 ( n12373,n13140,n10863 );
   not U13162 ( n13140,n10594 );
   nand U13163 ( n12375,n12190,n10594 );
   nor U13164 ( n13216,n12041,n12015,n11982,n13234 );
   not U13165 ( n13234,n11834 );
   nand U13166 ( n11834,n11841,n12402 );
   nand U13167 ( n12402,n11872,n10973 );
   nand U13168 ( n11841,n12524,n10624 );
   not U13169 ( n11982,n11992 );
   nand U13170 ( n11992,n12392,n12389 );
   nand U13171 ( n12389,n11986,n10612 );
   nand U13172 ( n12392,n12010,n10929 );
   nor U13173 ( n12015,n12121,n12388 );
   nor U13174 ( n12388,n10609,n12021 );
   nor U13175 ( n12121,n10918,n12036 );
   not U13176 ( n12036,n10609 );
   and U13177 ( n12041,n12073,n12075 );
   nand U13178 ( n12075,n12062,n10907 );
   not U13179 ( n12073,n12386 );
   nor U13180 ( n12386,n10907,n12062 );
   nand U13181 ( n13211,n12329,n13235 );
   nor U13182 ( n12329,n11132,n11130,n11142 );
   nand U13183 ( n13210,n13236,n13237,n12348 );
   nand U13184 ( n13237,n13235,n13214 );
   or U13185 ( n13236,n13238,n13152,n13235 );
   nand U13186 ( n13235,n13239,n13240,n13241,n13242 );
   nand U13187 ( n13242,n13243,n13244,n13245,n13246 );
   nor U13188 ( n13246,n13247,n13248,n13249 );
   nor U13189 ( n13249,n13250,n13251 );
   nor U13190 ( n13248,n13252,n13253 );
   nand U13191 ( n13245,n13254,n13255,n13256,n13257 );
   nor U13192 ( n13257,n13258,n13259,n13260,n13261 );
   nor U13193 ( n13261,n13262,n13263,n13264 );
   and U13194 ( n13262,n13265,n12114 );
   nor U13195 ( n13260,n13266,n13267,n13268 );
   not U13196 ( n13267,n13269 );
   not U13197 ( n13259,n13270 );
   nand U13198 ( n13256,n13271,n13272,n13273,n13274 );
   nor U13199 ( n13274,n13275,n13276 );
   nor U13200 ( n13275,n13277,n13278 );
   nand U13201 ( n13273,n13279,n13280 );
   nand U13202 ( n13279,n13281,n13282 );
   nand U13203 ( n13282,n13283,n13284 );
   nand U13204 ( n13281,n13285,n13286 );
   nand U13205 ( n13272,n13287,n13288,n13289 );
   nand U13206 ( n13271,n13287,n13290,n13291,n13292 );
   nand U13207 ( n13292,n13293,n13294 );
   or U13208 ( n13291,n13288,n13289 );
   and U13209 ( n13289,n13295,n13296 );
   nand U13210 ( n13296,n13265,n10615 );
   nand U13211 ( n13295,n13297,n11959 );
   nand U13212 ( n13288,n13298,n13299 );
   nand U13213 ( n13299,n11959,n13265 );
   nand U13214 ( n13298,n13297,n10615 );
   nand U13215 ( n13290,n13300,n13301 );
   or U13216 ( n13301,n13294,n13293 );
   and U13217 ( n13293,n13302,n13303 );
   nand U13218 ( n13303,n11913,n13265 );
   nand U13219 ( n13302,n13297,n10618 );
   nand U13220 ( n13294,n13304,n13305 );
   nand U13221 ( n13305,n13265,n10618 );
   nand U13222 ( n13304,n13297,n11913 );
   nand U13223 ( n13300,n13306,n13307 );
   nand U13224 ( n13307,n13308,n13309 );
   nand U13225 ( n13309,n13310,n13311 );
   nand U13226 ( n13308,n13312,n13313 );
   nand U13227 ( n13313,n13314,n13315 );
   nand U13228 ( n13312,n13316,n13317,n13318,n13319 );
   nand U13229 ( n13319,n13320,n13321,n13322 );
   nand U13230 ( n13318,n13323,n13321,n13324 );
   nand U13231 ( n13324,n13325,n13326 );
   nand U13232 ( n13326,n13327,n13328,n13329 );
   not U13233 ( n13327,n13330 );
   nand U13234 ( n13325,n13331,n13332 );
   nand U13235 ( n13332,n13330,n13333 );
   nand U13236 ( n13333,n13329,n13328 );
   nand U13237 ( n13328,n13334,n13335 );
   and U13238 ( n13329,n13336,n13337,n13338,n13339 );
   nand U13239 ( n13339,n13340,n13341,n13342,n13343 );
   nand U13240 ( n13340,n11679,n13265 );
   nand U13241 ( n13338,n13344,n13345,n13346,n13347 );
   nand U13242 ( n13345,n11042,n13265 );
   nand U13243 ( n13337,n13348,n13349,n13350,n13351 );
   nand U13244 ( n13350,n13352,n13353 );
   nand U13245 ( n13353,n13354,n13355,n13356 );
   nor U13246 ( n13356,n13357,n13358,n13359 );
   and U13247 ( n13359,n13360,n13232 );
   nor U13248 ( n13358,n13232,n11125,n13361 );
   nor U13249 ( n13357,n13297,n11450 );
   nand U13250 ( n11450,n13232,n11125 );
   not U13251 ( n13232,n10663 );
   nand U13252 ( n13355,n13360,n11125 );
   nand U13253 ( n13360,n12366,n13362 );
   nand U13254 ( n13362,n11130,n13153 );
   nand U13255 ( n13354,n13363,n13364 );
   or U13256 ( n13352,n13364,n13363 );
   and U13257 ( n13363,n13365,n13366 );
   nand U13258 ( n13366,n13265,n10660 );
   nand U13259 ( n13365,n13297,n11114 );
   nand U13260 ( n13364,n13367,n13368 );
   nand U13261 ( n13368,n13265,n11114 );
   nand U13262 ( n13367,n13297,n10660 );
   or U13263 ( n13349,n13369,n13370 );
   nand U13264 ( n13336,n13348,n13371 );
   nand U13265 ( n13371,n13372,n13373,n13374,n13375 );
   nand U13266 ( n13375,n13351,n13369,n13370 );
   and U13267 ( n13370,n13376,n13377 );
   nand U13268 ( n13377,n11104,n13265 );
   nand U13269 ( n13376,n13297,n10657 );
   nand U13270 ( n13369,n13378,n13379 );
   nand U13271 ( n13379,n13265,n10657 );
   nand U13272 ( n13378,n13297,n11104 );
   nand U13273 ( n13351,n13380,n13381 );
   or U13274 ( n13374,n13381,n13380 );
   and U13275 ( n13380,n13382,n13383 );
   nand U13276 ( n13383,n13265,n10654 );
   nand U13277 ( n13382,n13297,n11090 );
   nand U13278 ( n13381,n13384,n13385 );
   nand U13279 ( n13385,n13265,n11090 );
   nand U13280 ( n13384,n13297,n10654 );
   or U13281 ( n13373,n13386,n13387 );
   and U13282 ( n13348,n13344,n13388,n13389,n13390 );
   nand U13283 ( n13390,n13391,n13392 );
   nand U13284 ( n13392,n11623,n13346 );
   nand U13285 ( n13346,n13297,n10642 );
   not U13286 ( n13391,n13347 );
   nand U13287 ( n13347,n13393,n13394 );
   nand U13288 ( n13394,n13265,n10642 );
   nand U13289 ( n13393,n13297,n11042 );
   nand U13290 ( n13389,n13372,n13386,n13387 );
   and U13291 ( n13387,n13395,n13396 );
   nand U13292 ( n13396,n13265,n10651 );
   nand U13293 ( n13395,n13297,n11080 );
   nand U13294 ( n13386,n13397,n13398 );
   nand U13295 ( n13398,n11080,n13265 );
   nand U13296 ( n13397,n13297,n10651 );
   and U13297 ( n13372,n13399,n13400 );
   nand U13298 ( n13400,n13401,n13402 );
   nand U13299 ( n13388,n13399,n13403 );
   nand U13300 ( n13403,n13404,n13405 );
   or U13301 ( n13405,n13402,n13401 );
   and U13302 ( n13401,n13406,n13407 );
   nand U13303 ( n13407,n11582,n13265 );
   nand U13304 ( n13406,n13297,n10648 );
   nand U13305 ( n13402,n13408,n13409 );
   nand U13306 ( n13409,n13265,n10648 );
   nand U13307 ( n13408,n13297,n11582 );
   nand U13308 ( n13404,n13410,n13411 );
   or U13309 ( n13399,n13411,n13410 );
   and U13310 ( n13410,n13412,n13413 );
   nand U13311 ( n13413,n13265,n10645 );
   nand U13312 ( n13412,n13297,n11057 );
   nand U13313 ( n13411,n13414,n13415 );
   nand U13314 ( n13415,n13265,n11057 );
   nand U13315 ( n13414,n13297,n10645 );
   and U13316 ( n13344,n13416,n13343 );
   or U13317 ( n13343,n13335,n13334 );
   and U13318 ( n13334,n13417,n13418 );
   nand U13319 ( n13418,n11018,n13265 );
   nand U13320 ( n13417,n13297,n10636 );
   nand U13321 ( n13335,n13419,n13420 );
   nand U13322 ( n13420,n13265,n10636 );
   nand U13323 ( n13419,n13297,n11018 );
   nand U13324 ( n13416,n13421,n13422 );
   nand U13325 ( n13422,n11031,n13341 );
   nand U13326 ( n13341,n13297,n10639 );
   not U13327 ( n13421,n13342 );
   nand U13328 ( n13342,n13423,n13424 );
   nand U13329 ( n13424,n13265,n10639 );
   nand U13330 ( n13423,n13297,n11679 );
   nand U13331 ( n13330,n13425,n13426 );
   nand U13332 ( n13426,n13265,n10633 );
   nand U13333 ( n13425,n13297,n11737 );
   nand U13334 ( n13331,n13427,n13428 );
   nand U13335 ( n13428,n13265,n11737 );
   nand U13336 ( n13427,n13297,n10633 );
   nand U13337 ( n13321,n13429,n13430 );
   or U13338 ( n13323,n13320,n13322 );
   and U13339 ( n13322,n13431,n13432 );
   nand U13340 ( n13432,n13265,n10630 );
   nand U13341 ( n13431,n13297,n11782 );
   nand U13342 ( n13320,n13433,n13434 );
   nand U13343 ( n13434,n11782,n13265 );
   nand U13344 ( n13433,n13297,n10630 );
   or U13345 ( n13317,n13430,n13429 );
   and U13346 ( n13429,n13435,n13436 );
   nand U13347 ( n13436,n11812,n13265 );
   nand U13348 ( n13435,n13297,n10627 );
   nand U13349 ( n13430,n13437,n13438 );
   nand U13350 ( n13438,n13265,n10627 );
   nand U13351 ( n13437,n13297,n11812 );
   or U13352 ( n13316,n13315,n13314 );
   and U13353 ( n13314,n13439,n13440 );
   nand U13354 ( n13440,n13265,n12524 );
   nand U13355 ( n13439,n13297,n10624 );
   nand U13356 ( n13315,n13441,n13442 );
   nand U13357 ( n13442,n13265,n10624 );
   nand U13358 ( n13441,n13297,n12524 );
   or U13359 ( n13306,n13311,n13310 );
   and U13360 ( n13310,n13443,n13444 );
   nand U13361 ( n13444,n13265,n10621 );
   nand U13362 ( n13443,n13297,n11883 );
   nand U13363 ( n13311,n13445,n13446 );
   nand U13364 ( n13446,n13265,n11883 );
   nand U13365 ( n13445,n13297,n10621 );
   and U13366 ( n13287,n13280,n13447 );
   or U13367 ( n13447,n13284,n13283 );
   and U13368 ( n13283,n13448,n13449 );
   nand U13369 ( n13449,n13265,n10612 );
   nand U13370 ( n13448,n13297,n11986 );
   nand U13371 ( n13284,n13450,n13451 );
   nand U13372 ( n13451,n11986,n13265 );
   nand U13373 ( n13450,n13297,n10612 );
   or U13374 ( n13280,n13286,n13285 );
   and U13375 ( n13285,n13452,n13453 );
   nand U13376 ( n13453,n13265,n10609 );
   nand U13377 ( n13452,n13297,n12021 );
   nand U13378 ( n13286,n13454,n13455 );
   nand U13379 ( n13455,n12021,n13265 );
   nand U13380 ( n13454,n13297,n10609 );
   nand U13381 ( n13255,n13456,n13278,n13277 );
   and U13382 ( n13277,n13457,n13458 );
   nand U13383 ( n13458,n12044,n13265 );
   nand U13384 ( n13457,n13297,n10606 );
   nand U13385 ( n13278,n13459,n13460 );
   nand U13386 ( n13460,n13265,n10606 );
   nand U13387 ( n13459,n13297,n12044 );
   not U13388 ( n13456,n13276 );
   nand U13389 ( n13276,n13269,n13461 );
   nand U13390 ( n13461,n13268,n13266 );
   nand U13391 ( n13266,n13462,n13463 );
   nand U13392 ( n13463,n12071,n13265 );
   nand U13393 ( n13462,n13297,n10603 );
   and U13394 ( n13268,n13464,n13465 );
   nand U13395 ( n13465,n13265,n10603 );
   nand U13396 ( n13464,n13297,n12071 );
   nand U13397 ( n13269,n13263,n13466 );
   or U13398 ( n13466,n12114,n13264 );
   nor U13399 ( n13264,n13361,n12139 );
   and U13400 ( n13263,n13467,n13468 );
   nand U13401 ( n13468,n13265,n10600 );
   nand U13402 ( n13467,n13297,n12114 );
   nand U13403 ( n13254,n13469,n13470 );
   nand U13404 ( n13243,n13270,n13471,n13472 );
   nand U13405 ( n13472,n13473,n13474 );
   or U13406 ( n13474,n13470,n13469 );
   and U13407 ( n13469,n13475,n13476 );
   nand U13408 ( n13476,n12153,n13265 );
   nand U13409 ( n13475,n13297,n10597 );
   nand U13410 ( n13470,n13477,n13478 );
   nand U13411 ( n13478,n13265,n10597 );
   nand U13412 ( n13477,n13297,n12153 );
   nand U13413 ( n13473,n13479,n13480 );
   not U13414 ( n13471,n13258 );
   nor U13415 ( n13258,n13480,n13479 );
   and U13416 ( n13479,n13481,n13482 );
   nand U13417 ( n13482,n13265,n10594 );
   nand U13418 ( n13481,n13297,n12190 );
   nand U13419 ( n13480,n13483,n13484 );
   nand U13420 ( n13484,n12190,n13265 );
   nand U13421 ( n13483,n13297,n10594 );
   nand U13422 ( n13270,n13252,n13253 );
   nand U13423 ( n13253,n13485,n13486 );
   nand U13424 ( n13486,n13265,n10591 );
   nand U13425 ( n13485,n13297,n10853 );
   and U13426 ( n13252,n13487,n13488 );
   nand U13427 ( n13488,n10853,n13265 );
   nand U13428 ( n13487,n13297,n10591 );
   nand U13429 ( n13241,n13489,n13490 );
   nand U13430 ( n13490,n13491,n13492 );
   nand U13431 ( n13492,n13251,n13244,n13250 );
   and U13432 ( n13250,n13493,n13494 );
   nand U13433 ( n13494,n12235,n13265 );
   nand U13434 ( n13493,n13297,n10588 );
   nand U13435 ( n13244,n13495,n13496 );
   nand U13436 ( n13251,n13497,n13498 );
   nand U13437 ( n13498,n13265,n10588 );
   nand U13438 ( n13497,n13297,n12235 );
   or U13439 ( n13491,n13496,n13495 );
   and U13440 ( n13495,n13499,n13500 );
   nand U13441 ( n13500,n13265,n10585 );
   nand U13442 ( n13499,n13297,n12264 );
   nand U13443 ( n13496,n13501,n13502 );
   nand U13444 ( n13502,n12264,n13265 );
   nand U13445 ( n13501,n13297,n10585 );
   not U13446 ( n13489,n13247 );
   nand U13447 ( n13247,n13503,n13504,n13505,n13506 );
   or U13448 ( n13504,n13507,n13508 );
   nand U13449 ( n13240,n13509,n13506 );
   nand U13450 ( n13506,n13510,n13511 );
   nand U13451 ( n13509,n13512,n13513,n13514 );
   nand U13452 ( n13514,n13515,n13516 );
   nand U13453 ( n13513,n13517,n13518,n13519 );
   nand U13454 ( n13512,n13503,n13520 );
   nand U13455 ( n13520,n13521,n13522 );
   nand U13456 ( n13522,n13505,n13507,n13508 );
   and U13457 ( n13508,n13523,n13524 );
   nand U13458 ( n13524,n12300,n13265 );
   nand U13459 ( n13523,n13297,n10582 );
   nand U13460 ( n13507,n13525,n13526 );
   nand U13461 ( n13526,n10582,n13265 );
   nand U13462 ( n13525,n13297,n12300 );
   nand U13463 ( n13505,n13527,n13528 );
   or U13464 ( n13521,n13528,n13527 );
   and U13465 ( n13527,n13529,n13530 );
   nand U13466 ( n13530,n10579,n13265 );
   nand U13467 ( n13529,n13297,n12336 );
   nand U13468 ( n13528,n13531,n13532 );
   nand U13469 ( n13532,n12336,n13265 );
   nand U13470 ( n13531,n13297,n10579 );
   and U13471 ( n13503,n13518,n13533 );
   or U13472 ( n13533,n13517,n13519 );
   and U13473 ( n13519,n13534,n13535 );
   nand U13474 ( n13535,n10791,n13265 );
   nand U13475 ( n13534,n13297,n10576 );
   nand U13476 ( n13517,n13536,n13537 );
   nand U13477 ( n13537,n13265,n10576 );
   nand U13478 ( n13536,n13297,n10791 );
   not U13479 ( n10791,n12513 );
   nand U13480 ( n12513,n13538,n13539,n13075 );
   nand U13481 ( n13539,n11416,n13540 );
   or U13482 ( n13538,n11416,n11400 );
   or U13483 ( n13518,n13516,n13515 );
   and U13484 ( n13515,n13541,n13542 );
   nand U13485 ( n13542,n10780,n13265 );
   nand U13486 ( n13541,n13297,n10573 );
   nand U13487 ( n13516,n13543,n13544 );
   nand U13488 ( n13544,n10573,n13265 );
   nand U13489 ( n10573,n13545,n13546,n13547 );
   nand U13490 ( n13547,p2_reg2_reg_30_,n13548 );
   nand U13491 ( n13546,p2_reg0_reg_30_,n13549 );
   nand U13492 ( n13545,p2_reg1_reg_30_,n13550 );
   nand U13493 ( n13543,n13297,n10780 );
   not U13494 ( n10780,n12523 );
   nand U13495 ( n12523,n13551,n13552,n13075 );
   or U13496 ( n13552,n11414,p1_datao_reg_30_ );
   nand U13497 ( n13551,n13553,n11414 );
   or U13498 ( n13239,n13511,n13510 );
   and U13499 ( n13510,n13554,n13555 );
   nand U13500 ( n13555,n10771,n13265 );
   nand U13501 ( n13554,n13297,n10570 );
   nand U13502 ( n13511,n13556,n13557 );
   nand U13503 ( n13557,n13265,n10570 );
   nand U13504 ( n10570,n13558,n13559,n13560 );
   nand U13505 ( n13560,p2_reg2_reg_31_,n13548 );
   nand U13506 ( n13559,p2_reg0_reg_31_,n13549 );
   nand U13507 ( n13558,p2_reg1_reg_31_,n13550 );
   not U13508 ( n12366,n12522 );
   nand U13509 ( n13556,n13297,n10771 );
   not U13510 ( n10771,n13230 );
   nand U13511 ( n13230,n13561,n13562,n13075 );
   or U13512 ( n13562,n11414,p1_datao_reg_31_ );
   nand U13513 ( n13561,n11414,n13563 );
   nor U13514 ( n13567,n13568,n13569,n13570 );
   nor U13515 ( n13570,n11979,n13571 );
   not U13516 ( n11979,n10615 );
   nor U13517 ( n13569,n13572,n10951 );
   nor U13518 ( n13568,p2_state_reg,n13573 );
   nand U13519 ( n13566,n13574,n10621 );
   or U13520 ( n13565,n13575,n13576 );
   xor U13521 ( n13575,n13577,n13578 );
   xor U13522 ( n13577,n13579,n13580 );
   nand U13523 ( n13564,n11893,n13581 );
   nor U13524 ( n13585,n13586,n13587,n13588 );
   nor U13525 ( n13588,n12324,n13571 );
   nor U13526 ( n13587,n10850,n13589 );
   nor U13527 ( n13586,p2_state_reg,n13590 );
   nand U13528 ( n13584,n12264,n13591 );
   nand U13529 ( n13583,n13592,n13593,n13594 );
   nand U13530 ( n13593,n13595,n13596,n13597 );
   nand U13531 ( n13597,n13598,n13599 );
   nand U13532 ( n13595,n13600,n13601 );
   nand U13533 ( n13592,n13598,n13602,n13603 );
   nand U13534 ( n13582,n13604,n13605 );
   nor U13535 ( n13609,n12899,n13610,n13611 );
   nor U13536 ( n13611,n11077,n13589 );
   nor U13537 ( n13610,n11054,n13571 );
   nor U13538 ( n12899,p2_state_reg,n13612 );
   not U13539 ( n13612,p2_reg3_reg_6_ );
   nand U13540 ( n13608,n11597,n13581 );
   nand U13541 ( n13607,n13613,n13614,n13594 );
   or U13542 ( n13614,n13615,n13616 );
   xor U13543 ( n13615,n13617,n13618 );
   nand U13544 ( n13613,n13619,n13620,n13616 );
   nand U13545 ( n13606,n13591,n11057 );
   nor U13546 ( n13624,n13625,n13626,n13627 );
   nor U13547 ( n13627,n12062,n13571 );
   nor U13548 ( n13626,n12010,n13589 );
   nor U13549 ( n13625,p2_state_reg,n13628 );
   nand U13550 ( n13623,n12021,n13591 );
   or U13551 ( n13622,n13629,n13576 );
   xor U13552 ( n13629,n13630,n13631 );
   xor U13553 ( n13630,n13632,n13633 );
   nand U13554 ( n13621,n13634,n13581 );
   nand U13555 ( n13638,n11104,n13591 );
   nor U13556 ( n13637,n13639,n13640 );
   nor U13557 ( n13640,n13641,n11491 );
   not U13558 ( n11491,p2_reg3_reg_2_ );
   nor U13559 ( n13639,n13576,n13642,n13643 );
   and U13560 ( n13643,n13644,n13645,n13646 );
   nor U13561 ( n13642,n13644,n13647 );
   xor U13562 ( n13647,n13648,n13649 );
   nand U13563 ( n13636,n13650,n10654 );
   nand U13564 ( n13635,n13574,n10660 );
   nor U13565 ( n13654,n13655,n13656,n13657 );
   nor U13566 ( n13657,n13658,n11752 );
   not U13567 ( n11752,n13659 );
   nor U13568 ( n13656,n13572,n10995 );
   and U13569 ( n13655,p2_u3152,p2_reg3_reg_11_ );
   nand U13570 ( n13653,n13650,n10627 );
   nand U13571 ( n13652,n13594,n13660 );
   nand U13572 ( n13660,n13661,n13662,n13663 );
   nand U13573 ( n13663,n13664,n13665 );
   nand U13574 ( n13662,n13666,n13667,n13668 );
   not U13575 ( n13668,n13669 );
   nand U13576 ( n13661,n13670,n13669 );
   xor U13577 ( n13670,n13666,n13667 );
   nand U13578 ( n13651,n13574,n10633 );
   nor U13579 ( n13674,n13675,n13676,n13677 );
   nor U13580 ( n13677,n12139,n13589 );
   nor U13581 ( n13676,n13572,n10875 );
   nor U13582 ( n13675,p2_state_reg,n13678 );
   nand U13583 ( n13673,n13650,n10594 );
   or U13584 ( n13672,n13679,n13576 );
   xor U13585 ( n13679,n13680,n13681 );
   xor U13586 ( n13680,n13682,n13683 );
   nand U13587 ( n13671,n13684,n13605 );
   nor U13588 ( n13688,n13689,n13690,n13691 );
   nor U13589 ( n13691,n10973,n13572 );
   nor U13590 ( n13690,n13658,n11820 );
   not U13591 ( n11820,n13692 );
   and U13592 ( n13689,p2_u3152,p2_reg3_reg_13_ );
   nand U13593 ( n13687,n13574,n10627 );
   nand U13594 ( n13694,n13695,n13696 );
   nand U13595 ( n13696,n13697,n13698 );
   nand U13596 ( n13693,n13699,n13700,n13697,n13698 );
   nand U13597 ( n13699,n13701,n13702 );
   nand U13598 ( n13685,n13650,n10621 );
   nor U13599 ( n13706,n13707,n13708,n13709 );
   nor U13600 ( n13709,n12139,n13571 );
   not U13601 ( n12139,n10600 );
   nor U13602 ( n13708,n12062,n13589 );
   not U13603 ( n12062,n10606 );
   nor U13604 ( n13707,p2_state_reg,n13710 );
   nand U13605 ( n13705,n12071,n13591 );
   nand U13606 ( n13704,n13711,n13594 );
   xor U13607 ( n13711,n13712,n13713 );
   nand U13608 ( n13713,n13714,n13715 );
   nand U13609 ( n13703,n13716,n13605 );
   nand U13610 ( n13720,n13594,n13721 );
   xor U13611 ( n13721,n13722,n13723 );
   nand U13612 ( n13723,n13724,n13725 );
   nand U13613 ( n13725,n13726,n10663 );
   nand U13614 ( n13724,n13727,n13728 );
   nand U13615 ( n13719,p2_reg3_reg_0_,n13729 );
   not U13616 ( n13729,n13641 );
   nand U13617 ( n13718,n13591,n11125 );
   nand U13618 ( n13717,n13650,n10660 );
   nor U13619 ( n13733,n12818,n13734,n13735 );
   nor U13620 ( n13735,n11041,n13589 );
   nor U13621 ( n13734,n13572,n11691 );
   nor U13622 ( n12818,p2_state_reg,n13736 );
   nand U13623 ( n13732,n11692,n13581 );
   xor U13624 ( n13737,n13738,n13739 );
   xor U13625 ( n13738,n13740,n13741 );
   nand U13626 ( n13730,n13650,n10633 );
   nor U13627 ( n13745,n12958,n13746,n13747 );
   nor U13628 ( n13747,n11101,n13589 );
   not U13629 ( n11101,n10654 );
   nor U13630 ( n13746,n11077,n13571 );
   not U13631 ( n11077,n10648 );
   nor U13632 ( n12958,p2_state_reg,n13748 );
   nand U13633 ( n13744,n11080,n13591 );
   or U13634 ( n13743,n13749,n13576 );
   xor U13635 ( n13749,n13750,n13751 );
   xor U13636 ( n13750,n13752,n13753 );
   nand U13637 ( n13742,n11561,n13581 );
   nor U13638 ( n13757,n13758,n13759,n13760 );
   nor U13639 ( n13760,n10850,n13571 );
   not U13640 ( n10850,n10588 );
   nor U13641 ( n13759,n13572,n12199 );
   nor U13642 ( n13758,p2_state_reg,n13761 );
   nand U13643 ( n13756,n13574,n10594 );
   nand U13644 ( n13755,n13594,n13762 );
   xor U13645 ( n13762,n13763,n13764 );
   nand U13646 ( n13763,n13765,n13766 );
   nand U13647 ( n13754,n12200,n13605 );
   nor U13648 ( n13770,n13771,n13772,n13773 );
   nor U13649 ( n13773,n13572,n10929 );
   nor U13650 ( n13772,n13658,n11969 );
   not U13651 ( n11969,n13774 );
   and U13652 ( n13771,p2_u3152,p2_reg3_reg_17_ );
   nand U13653 ( n13769,n13574,n10615 );
   nand U13654 ( n13776,n13777,n13778 );
   nand U13655 ( n13778,n13779,n13780 );
   nand U13656 ( n13775,n13781,n13782,n13779,n13780 );
   nand U13657 ( n13781,n13783,n13784 );
   nand U13658 ( n13767,n13650,n10609 );
   nor U13659 ( n13788,n12929,n13789,n13790 );
   nor U13660 ( n13790,n11089,n13589 );
   not U13661 ( n11089,n10651 );
   nor U13662 ( n13789,n13194,n13571 );
   nor U13663 ( n12929,p2_state_reg,n13791 );
   nand U13664 ( n13787,n11571,n13581 );
   or U13665 ( n13786,n13792,n13576 );
   xor U13666 ( n13792,n13793,n13794 );
   xor U13667 ( n13793,n13795,n13796 );
   nand U13668 ( n13785,n11582,n13591 );
   nor U13669 ( n13800,n13801,n13802,n13803 );
   nor U13670 ( n13803,n12010,n13571 );
   not U13671 ( n12010,n10612 );
   nor U13672 ( n13802,n13658,n11924 );
   not U13673 ( n11924,n13804 );
   nor U13674 ( n13801,p2_state_reg,n13805 );
   nand U13675 ( n13799,n11959,n13591 );
   or U13676 ( n13807,n13808,n13809 );
   xor U13677 ( n13808,n13810,n13811 );
   nand U13678 ( n13806,n13782,n13784,n13809 );
   nand U13679 ( n13797,n13574,n10618 );
   nor U13680 ( n13815,n13816,n13817,n13818 );
   nor U13681 ( n13818,n12288,n13571 );
   nor U13682 ( n13817,n13572,n10841 );
   and U13683 ( n13816,p2_u3152,p2_reg3_reg_25_ );
   nand U13684 ( n13814,n13574,n10591 );
   nand U13685 ( n13813,n13819,n13820,n13594 );
   nand U13686 ( n13820,n13600,n13596,n13601 );
   or U13687 ( n13819,n13821,n13601 );
   xor U13688 ( n13821,n13822,n13823 );
   nand U13689 ( n13812,n12217,n13605 );
   nor U13690 ( n13827,n12734,n13828,n13829 );
   nor U13691 ( n13829,n11872,n13571 );
   nor U13692 ( n13828,n11802,n13589 );
   nor U13693 ( n12734,p2_state_reg,n13830 );
   nand U13694 ( n13826,n11812,n13591 );
   nand U13695 ( n13825,n13831,n13594 );
   xor U13696 ( n13831,n13701,n13832 );
   nand U13697 ( n13832,n13700,n13702 );
   nand U13698 ( n13824,n13833,n13581 );
   nor U13699 ( n13837,n13838,n13839,n13840 );
   nor U13700 ( n13840,n13572,n10885 );
   nor U13701 ( n13839,n12106,n13589 );
   not U13702 ( n12106,n10603 );
   nor U13703 ( n13838,p2_state_reg,n13841 );
   nand U13704 ( n13836,n13650,n10597 );
   nand U13705 ( n13835,n13842,n13843,n13594 );
   nand U13706 ( n13843,n13844,n13845 );
   nand U13707 ( n13845,n13846,n13847 );
   nand U13708 ( n13842,n13848,n13714,n13846,n13847 );
   nand U13709 ( n13848,n13712,n13715 );
   nand U13710 ( n13834,n12085,n13605 );
   nand U13711 ( n13852,n13591,n11114 );
   nor U13712 ( n13851,n13853,n13854 );
   nor U13713 ( n13854,n13641,n11471 );
   not U13714 ( n11471,p2_reg3_reg_1_ );
   nor U13715 ( n13641,n13581,p2_u3152 );
   nor U13716 ( n13853,n13855,n13576 );
   xor U13717 ( n13855,n13856,n13857 );
   xor U13718 ( n13856,n13858,n13859 );
   nand U13719 ( n13850,n13650,n10657 );
   nand U13720 ( n13849,n13574,n10663 );
   nor U13721 ( n13863,n13864,n13865,n13866 );
   nor U13722 ( n13866,n11054,n13589 );
   not U13723 ( n11054,n10642 );
   nor U13724 ( n13865,n13658,n11653 );
   nor U13725 ( n13864,p2_state_reg,n13867 );
   nand U13726 ( n13862,n11679,n13591 );
   xor U13727 ( n13868,n13869,n13870 );
   xor U13728 ( n13869,n13871,n13872 );
   nand U13729 ( n13860,n13650,n10636 );
   nor U13730 ( n13876,n13877,n13878,n13879 );
   nor U13731 ( n13879,n12324,n13589 );
   not U13732 ( n12324,n10582 );
   and U13733 ( n13878,n13605,n12315 );
   nor U13734 ( n13877,p2_state_reg,n13880 );
   nand U13735 ( n13875,n12336,n13591 );
   nand U13736 ( n13882,n13883,n13884 );
   nand U13737 ( n13883,n13885,n13886 );
   nand U13738 ( n13886,n13887,n13888 );
   nand U13739 ( n13881,n13889,n13890 );
   nand U13740 ( n13890,n13888,n13891 );
   nand U13741 ( n13891,n13885,n13892 );
   not U13742 ( n13889,n13884 );
   nand U13743 ( n13884,n13893,n13894,n13895,n13896 );
   or U13744 ( n13896,n12360,n13726 );
   nand U13745 ( n12360,n13897,n10804 );
   nand U13746 ( n13895,n13094,n13726 );
   nor U13747 ( n13094,n10579,n10804 );
   nand U13748 ( n13894,n12446,n13898 );
   nor U13749 ( n12446,n13897,n12336 );
   not U13750 ( n13897,n10579 );
   or U13751 ( n13893,n12362,n13898 );
   nand U13752 ( n12362,n12336,n10579 );
   not U13753 ( n12336,n10804 );
   nand U13754 ( n10804,n13899,n13900,n13075 );
   nand U13755 ( n13900,n11416,n13901 );
   or U13756 ( n13899,n11390,n11416 );
   nand U13757 ( n13873,n13650,n10576 );
   nand U13758 ( n10576,n13902,n13903,n13904,n13905 );
   nand U13759 ( n13905,n13906,n12347 );
   nor U13760 ( n12347,n13907,n13908,n13880 );
   nand U13761 ( n13904,p2_reg0_reg_29_,n13549 );
   nand U13762 ( n13903,p2_reg1_reg_29_,n13550 );
   nand U13763 ( n13902,p2_reg2_reg_29_,n13548 );
   nor U13764 ( n13912,n13913,n13914,n13915 );
   nor U13765 ( n13915,n13658,n12027 );
   not U13766 ( n12027,n13916 );
   nor U13767 ( n13914,n13572,n10907 );
   and U13768 ( n13913,p2_u3152,p2_reg3_reg_19_ );
   nand U13769 ( n13911,n13650,n10603 );
   nand U13770 ( n13917,n13918,n13919,n13920 );
   nand U13771 ( n13920,n13921,n13922 );
   nand U13772 ( n13919,n13923,n13924,n13925 );
   not U13773 ( n13925,n13926 );
   nand U13774 ( n13918,n13927,n13926 );
   xor U13775 ( n13927,n13923,n13924 );
   nand U13776 ( n13909,n13574,n10609 );
   nor U13777 ( n13931,n13932,n13933,n13934 );
   nor U13778 ( n13934,p2_reg3_reg_3_,n13658 );
   not U13779 ( n13658,n13581 );
   nor U13780 ( n13933,p2_state_reg,n13935 );
   nor U13781 ( n13932,n11113,n13589 );
   not U13782 ( n11113,n10657 );
   nand U13783 ( n13930,n13650,n10651 );
   nand U13784 ( n13929,n13936,n13937,n13594 );
   nand U13785 ( n13937,n13938,n13646,n13939,n13940 );
   nand U13786 ( n13938,n13645,n13941 );
   nand U13787 ( n13936,n13942,n13943 );
   nand U13788 ( n13943,n13939,n13940 );
   nand U13789 ( n13928,n13591,n11090 );
   nor U13790 ( n13947,n13948,n13949,n13950 );
   nor U13791 ( n13950,n11802,n13571 );
   not U13792 ( n11802,n10630 );
   nor U13793 ( n13949,n11007,n13572 );
   nor U13794 ( n13948,p2_state_reg,n13951 );
   nand U13795 ( n13946,n13574,n10636 );
   or U13796 ( n13945,n13576,n13952 );
   xor U13797 ( n13952,n13953,n13954 );
   xor U13798 ( n13954,n13955,n13956 );
   nand U13799 ( n13944,n11711,n13581 );
   nor U13800 ( n13960,n13961,n13962,n13963 );
   nor U13801 ( n13963,n12226,n13571 );
   not U13802 ( n12226,n10591 );
   nor U13803 ( n13962,n13572,n10863 );
   nor U13804 ( n13961,p2_state_reg,n13964 );
   nand U13805 ( n13959,n13574,n10597 );
   or U13806 ( n13958,n13965,n13576 );
   xor U13807 ( n13965,n13966,n13967 );
   xor U13808 ( n13966,n13968,n13969 );
   nand U13809 ( n13957,n12161,n13605 );
   nor U13810 ( n13973,n13974,n13975,n13976 );
   nor U13811 ( n13976,n11872,n13589 );
   not U13812 ( n11872,n10624 );
   nor U13813 ( n13975,n10963,n13572 );
   nor U13814 ( n13974,p2_state_reg,n13977 );
   nand U13815 ( n13972,n13978,n13581 );
   xor U13816 ( n13979,n13980,n13981 );
   xor U13817 ( n13981,n13982,n13983 );
   nand U13818 ( n13970,n13650,n10618 );
   nor U13819 ( n13987,n13988,n13989,n13990 );
   nor U13820 ( n13990,n12288,n13589 );
   nor U13821 ( n13989,n13572,n10817 );
   nor U13822 ( n13988,p2_state_reg,n13907 );
   not U13823 ( n13907,p2_reg3_reg_27_ );
   nand U13824 ( n13986,n13650,n10579 );
   nand U13825 ( n10579,n13991,n13992,n13993,n13994 );
   nand U13826 ( n13994,n13906,n12315 );
   xor U13827 ( n12315,n13880,n13995 );
   nand U13828 ( n13995,p2_reg3_reg_27_,n13996 );
   not U13829 ( n13880,p2_reg3_reg_28_ );
   nand U13830 ( n13993,p2_reg0_reg_28_,n13549 );
   nand U13831 ( n13992,p2_reg1_reg_28_,n13550 );
   nand U13832 ( n13991,p2_reg2_reg_28_,n13548 );
   nand U13833 ( n13985,n13997,n13594 );
   xor U13834 ( n13997,n13892,n13998 );
   nand U13835 ( n13998,n13885,n13888 );
   nand U13836 ( n13888,n13999,n14000 );
   nand U13837 ( n14000,n14001,n10582 );
   xor U13838 ( n13999,n13726,n12300 );
   and U13839 ( n13885,n14002,n14003 );
   or U13840 ( n14003,n12434,n13728 );
   nand U13841 ( n12434,n12300,n10582 );
   not U13842 ( n12300,n10817 );
   or U13843 ( n14002,n12447,n13898 );
   nand U13844 ( n12447,n10817,n10582 );
   nand U13845 ( n10582,n14004,n14005,n14006,n14007 );
   nand U13846 ( n14007,n13906,n12281 );
   nand U13847 ( n14006,p2_reg0_reg_27_,n13549 );
   nand U13848 ( n14005,p2_reg1_reg_27_,n13550 );
   nand U13849 ( n14004,p2_reg2_reg_27_,n13548 );
   nand U13850 ( n10817,n14008,n14009,n13075 );
   nand U13851 ( n14009,n11416,n14010 );
   or U13852 ( n14008,n11380,n11416 );
   not U13853 ( n13892,n13887 );
   nand U13854 ( n13887,n13598,n14011 );
   nand U13855 ( n14011,n13603,n13602 );
   nand U13856 ( n13602,n14012,n13596 );
   or U13857 ( n13596,n13823,n13822 );
   not U13858 ( n14012,n13601 );
   nand U13859 ( n13601,n13765,n14013 );
   nand U13860 ( n14013,n14014,n13766 );
   nand U13861 ( n13766,n14015,n14016 );
   nand U13862 ( n14016,n14001,n10591 );
   xor U13863 ( n14015,n13726,n10853 );
   not U13864 ( n14014,n13764 );
   nand U13865 ( n13764,n14017,n14018 );
   nand U13866 ( n14018,n13967,n14019 );
   or U13867 ( n14019,n13969,n13968 );
   xor U13868 ( n13967,n13726,n12190 );
   not U13869 ( n12190,n10863 );
   nand U13870 ( n10863,n14020,n14021,n13075 );
   nand U13871 ( n14021,n11416,n14022 );
   or U13872 ( n14020,n11345,n11416 );
   nand U13873 ( n14017,n13968,n13969 );
   nand U13874 ( n13969,n14023,n14024 );
   nand U13875 ( n14024,n14025,n13683 );
   nand U13876 ( n13683,n14026,n13847 );
   nand U13877 ( n13847,n14027,n14028 );
   nand U13878 ( n14028,n14001,n10600 );
   xor U13879 ( n14027,n13726,n12114 );
   nand U13880 ( n14026,n13844,n13846 );
   nand U13881 ( n13846,n14001,n10600,n14029 );
   xor U13882 ( n14029,n13728,n12114 );
   not U13883 ( n12114,n10885 );
   nand U13884 ( n10885,n14030,n14031,n13075 );
   nand U13885 ( n14031,n11416,n14032 );
   or U13886 ( n14030,n11328,n11416 );
   nand U13887 ( n10600,n14033,n14034,n14035,n14036 );
   nand U13888 ( n14036,n13906,n12085 );
   xor U13889 ( n12085,n13841,n14037 );
   nand U13890 ( n14035,p2_reg0_reg_21_,n13549 );
   nand U13891 ( n14034,p2_reg1_reg_21_,n13550 );
   nand U13892 ( n14033,p2_reg2_reg_21_,n13548 );
   and U13893 ( n13844,n13715,n14038 );
   nand U13894 ( n14038,n14039,n13714 );
   nand U13895 ( n13714,n14040,n14041 );
   nand U13896 ( n14041,n14001,n10603 );
   not U13897 ( n14039,n13712 );
   nor U13898 ( n13712,n13921,n14042 );
   and U13899 ( n14042,n13922,n14043 );
   nand U13900 ( n14043,n13926,n13924 );
   not U13901 ( n13922,n13923 );
   nand U13902 ( n13923,n14044,n14045 );
   nand U13903 ( n14045,n14046,n13633 );
   nand U13904 ( n13633,n14047,n13780 );
   nand U13905 ( n13780,n14048,n14049 );
   nand U13906 ( n14049,n14001,n10612 );
   xor U13907 ( n14048,n13726,n11986 );
   nand U13908 ( n14047,n13777,n13779 );
   nand U13909 ( n13779,n14001,n10612,n14050 );
   xor U13910 ( n14050,n13728,n11986 );
   not U13911 ( n11986,n10929 );
   nand U13912 ( n10929,n14051,n14052,n14053 );
   nand U13913 ( n14053,n12521,n12610 );
   nand U13914 ( n12610,n14054,n14055,n11303 );
   nand U13915 ( n14055,n11294,n14056 );
   not U13916 ( n11294,p2_ir_reg_17_ );
   nand U13917 ( n14054,p2_ir_reg_17_,n11293,p2_ir_reg_31_ );
   nand U13918 ( n14052,n14057,n14058 );
   nand U13919 ( n14051,n14059,n14060 );
   nand U13920 ( n10612,n14061,n14062,n14063,n14064 );
   nand U13921 ( n14064,n13906,n13774 );
   xor U13922 ( n13774,p2_reg3_reg_17_,n14065 );
   nand U13923 ( n14063,p2_reg0_reg_17_,n13549 );
   nand U13924 ( n14062,p2_reg1_reg_17_,n13550 );
   nand U13925 ( n14061,p2_reg2_reg_17_,n13548 );
   and U13926 ( n13777,n13784,n14066 );
   nand U13927 ( n14066,n13809,n13782 );
   nand U13928 ( n13782,n13810,n13811 );
   not U13929 ( n13809,n13783 );
   nand U13930 ( n13783,n14067,n14068 );
   nand U13931 ( n14068,n13578,n14069 );
   or U13932 ( n14069,n13579,n13580 );
   xor U13933 ( n13578,n13726,n11913 );
   not U13934 ( n11913,n10951 );
   nand U13935 ( n10951,n14070,n14071,n14072 );
   nand U13936 ( n14072,n12521,n12644 );
   nand U13937 ( n12644,n14073,n14074,n14075 );
   nand U13938 ( n14074,n11277,n14056 );
   nand U13939 ( n14073,p2_ir_reg_15_,n11276,p2_ir_reg_31_ );
   nand U13940 ( n14071,n14057,n14076 );
   nand U13941 ( n14070,n14059,n14077 );
   not U13942 ( n14077,p1_datao_reg_15_ );
   nand U13943 ( n14067,n13579,n13580 );
   nand U13944 ( n13580,n14078,n14079 );
   nand U13945 ( n14079,n14080,n13983 );
   nand U13946 ( n13983,n14081,n13698 );
   nand U13947 ( n13698,n14082,n14083 );
   nand U13948 ( n14083,n14001,n10624 );
   xor U13949 ( n14082,n13728,n10973 );
   nand U13950 ( n14081,n13695,n13697 );
   nand U13951 ( n13697,n14001,n10624,n14084 );
   xor U13952 ( n14084,n13726,n10973 );
   not U13953 ( n10973,n12524 );
   nand U13954 ( n12524,n14085,n14086,n14087 );
   nand U13955 ( n14087,n12695,n12521 );
   not U13956 ( n12695,n12717 );
   nand U13957 ( n12717,n14088,n14089,n14090 );
   nand U13958 ( n14089,n11260,n14056 );
   nand U13959 ( n14088,p2_ir_reg_13_,n11259,p2_ir_reg_31_ );
   nand U13960 ( n14086,n14057,n11261 );
   nand U13961 ( n14085,p1_datao_reg_13_,n14059 );
   nand U13962 ( n10624,n14091,n14092,n14093,n14094 );
   nand U13963 ( n14094,n13906,n13692 );
   xor U13964 ( n13692,p2_reg3_reg_13_,n14095 );
   nand U13965 ( n14093,p2_reg0_reg_13_,n13549 );
   nand U13966 ( n14092,p2_reg1_reg_13_,n13550 );
   nand U13967 ( n14091,p2_reg2_reg_13_,n13548 );
   and U13968 ( n13695,n13702,n14096 );
   nand U13969 ( n14096,n14097,n13700 );
   nand U13970 ( n13700,n14098,n14099 );
   nand U13971 ( n14099,n14001,n10627 );
   not U13972 ( n14097,n13701 );
   nor U13973 ( n13701,n13664,n14100 );
   and U13974 ( n14100,n13665,n14101 );
   nand U13975 ( n14101,n13669,n13667 );
   not U13976 ( n13665,n13666 );
   nand U13977 ( n13666,n14102,n14103 );
   nand U13978 ( n14103,n13953,n14104 );
   or U13979 ( n14104,n13956,n13955 );
   xor U13980 ( n13953,n13728,n11007 );
   not U13981 ( n11007,n11737 );
   nand U13982 ( n11737,n14105,n14106,n14107 );
   nand U13983 ( n14107,n12777,n12521 );
   not U13984 ( n12777,n12803 );
   nand U13985 ( n12803,n14108,n14109 );
   or U13986 ( n14109,p2_ir_reg_10_,p2_ir_reg_31_ );
   nand U13987 ( n14108,p2_ir_reg_31_,n11233 );
   nand U13988 ( n11233,n11242,n14110 );
   nand U13989 ( n14110,p2_ir_reg_10_,n14111 );
   nand U13990 ( n14106,n14057,n11234 );
   nand U13991 ( n14105,p1_datao_reg_10_,n14059 );
   nand U13992 ( n14102,n13955,n13956 );
   nand U13993 ( n13956,n14112,n14113 );
   nand U13994 ( n14113,n13739,n14114 );
   or U13995 ( n14114,n13741,n13740 );
   xor U13996 ( n13739,n11018,n13726 );
   not U13997 ( n11018,n11691 );
   nand U13998 ( n11691,n14115,n14116,n14117 );
   nand U13999 ( n14117,n12521,n12834 );
   nand U14000 ( n12834,n14118,n14119,n14111 );
   nand U14001 ( n14119,n14056,n11226 );
   nand U14002 ( n14118,p2_ir_reg_31_,n11217,p2_ir_reg_9_ );
   nand U14003 ( n14116,n14057,n14120 );
   not U14004 ( n14120,n11227 );
   nand U14005 ( n14115,n14059,n14121 );
   nand U14006 ( n14112,n13740,n13741 );
   nand U14007 ( n13741,n14122,n14123 );
   nand U14008 ( n14123,n14124,n13872 );
   nand U14009 ( n13872,n14125,n14126 );
   nand U14010 ( n14125,n14127,n14128 );
   or U14011 ( n14124,n13871,n13870 );
   nand U14012 ( n14122,n13870,n13871 );
   nand U14013 ( n13871,n14001,n10639 );
   xor U14014 ( n13870,n11679,n13726 );
   not U14015 ( n11679,n11031 );
   nand U14016 ( n11031,n14129,n14130,n14131 );
   nand U14017 ( n14131,n12521,n12859 );
   nand U14018 ( n12859,n14132,n14133 );
   or U14019 ( n14133,p2_ir_reg_31_,p2_ir_reg_8_ );
   nand U14020 ( n14132,p2_ir_reg_31_,n14134 );
   nand U14021 ( n14134,n11217,n11216 );
   nand U14022 ( n11216,p2_ir_reg_8_,n14135 );
   not U14023 ( n11217,n11225 );
   nand U14024 ( n14130,n14057,n14136 );
   not U14025 ( n14136,n11218 );
   nand U14026 ( n14129,n14059,n14137 );
   nand U14027 ( n13740,n14001,n10636 );
   nand U14028 ( n10636,n14138,n14139,n14140,n14141 );
   nand U14029 ( n14141,n13906,n11692 );
   xor U14030 ( n11692,p2_reg3_reg_9_,n14142 );
   nand U14031 ( n14140,p2_reg0_reg_9_,n13549 );
   nand U14032 ( n14139,p2_reg1_reg_9_,n13550 );
   nand U14033 ( n14138,p2_reg2_reg_9_,n13548 );
   nand U14034 ( n13955,n14001,n10633 );
   nand U14035 ( n10633,n14143,n14144,n14145,n14146 );
   nand U14036 ( n14146,n11711,n13906 );
   nor U14037 ( n11711,n14147,n14148 );
   and U14038 ( n14147,n13951,n14149 );
   nand U14039 ( n14149,p2_reg3_reg_9_,n14142 );
   nand U14040 ( n14145,p2_reg0_reg_10_,n13549 );
   nand U14041 ( n14144,p2_reg1_reg_10_,n13550 );
   nand U14042 ( n14143,p2_reg2_reg_10_,n13548 );
   nor U14043 ( n13664,n13667,n13669 );
   xor U14044 ( n13669,n13726,n11782 );
   not U14045 ( n11782,n10995 );
   nand U14046 ( n10995,n14150,n14151,n14152 );
   nand U14047 ( n14152,n12521,n12749 );
   nand U14048 ( n12749,n14153,n14154,n14155 );
   nand U14049 ( n14154,n11243,n14056 );
   nand U14050 ( n14153,p2_ir_reg_11_,n11242,p2_ir_reg_31_ );
   not U14051 ( n11242,n11241 );
   nand U14052 ( n14151,n14057,n14156 );
   not U14053 ( n14156,n11244 );
   nand U14054 ( n14150,n14059,n14157 );
   not U14055 ( n14157,p1_datao_reg_11_ );
   nand U14056 ( n13667,n14001,n10630 );
   nand U14057 ( n10630,n14158,n14159,n14160,n14161 );
   nand U14058 ( n14161,n13906,n13659 );
   xor U14059 ( n13659,p2_reg3_reg_11_,n14148 );
   nand U14060 ( n14160,p2_reg0_reg_11_,n13549 );
   nand U14061 ( n14159,p2_reg1_reg_11_,n13550 );
   nand U14062 ( n14158,p2_reg2_reg_11_,n13548 );
   nand U14063 ( n13702,n14001,n10627,n14162 );
   not U14064 ( n14162,n14098 );
   xor U14065 ( n14098,n13726,n11812 );
   not U14066 ( n11812,n10985 );
   nand U14067 ( n10985,n14163,n14164,n14165 );
   nand U14068 ( n14165,n12521,n12754 );
   nand U14069 ( n12754,n14166,n14167 );
   or U14070 ( n14167,p2_ir_reg_12_,p2_ir_reg_31_ );
   nand U14071 ( n14166,p2_ir_reg_31_,n11250 );
   nand U14072 ( n11250,n11259,n14168 );
   nand U14073 ( n14168,p2_ir_reg_12_,n14155 );
   not U14074 ( n11259,n11258 );
   nand U14075 ( n14164,n14057,n14169 );
   not U14076 ( n14169,n11251 );
   nand U14077 ( n14163,n14059,n14170 );
   nand U14078 ( n10627,n14171,n14172,n14173,n14174 );
   nand U14079 ( n14174,n13833,n13906 );
   not U14080 ( n13833,n11793 );
   nand U14081 ( n11793,n14175,n14176 );
   nand U14082 ( n14175,n13830,n14177 );
   nand U14083 ( n14177,p2_reg3_reg_11_,n14148 );
   not U14084 ( n13830,p2_reg3_reg_12_ );
   nand U14085 ( n14173,p2_reg0_reg_12_,n13549 );
   nand U14086 ( n14172,p2_reg1_reg_12_,n13550 );
   nand U14087 ( n14171,p2_reg2_reg_12_,n13548 );
   nand U14088 ( n14080,n14178,n13980 );
   or U14089 ( n14078,n13980,n14178 );
   not U14090 ( n14178,n13982 );
   nand U14091 ( n13982,n14001,n10621 );
   nand U14092 ( n10621,n14179,n14180,n14181,n14182 );
   nand U14093 ( n14182,n13978,n13906 );
   not U14094 ( n13978,n11854 );
   nand U14095 ( n11854,n14183,n14184 );
   nand U14096 ( n14183,n13977,n14185 );
   nand U14097 ( n14185,p2_reg3_reg_13_,n14095 );
   not U14098 ( n13977,p2_reg3_reg_14_ );
   nand U14099 ( n14181,p2_reg0_reg_14_,n13549 );
   nand U14100 ( n14180,p2_reg1_reg_14_,n13550 );
   nand U14101 ( n14179,p2_reg2_reg_14_,n13548 );
   xor U14102 ( n13980,n13726,n10963 );
   not U14103 ( n10963,n11883 );
   nand U14104 ( n11883,n14186,n14187,n14188 );
   nand U14105 ( n14188,n12670,n12521 );
   not U14106 ( n12670,n12680 );
   nand U14107 ( n12680,n14189,n14190 );
   or U14108 ( n14190,p2_ir_reg_14_,p2_ir_reg_31_ );
   nand U14109 ( n14189,p2_ir_reg_31_,n11267 );
   nand U14110 ( n11267,n11276,n14191 );
   nand U14111 ( n14191,p2_ir_reg_14_,n14090 );
   not U14112 ( n11276,n11275 );
   nand U14113 ( n14187,n14057,n11268 );
   nand U14114 ( n14186,p1_datao_reg_14_,n14059 );
   nand U14115 ( n13579,n14001,n10618 );
   nand U14116 ( n10618,n14192,n14193,n14194,n14195 );
   nand U14117 ( n14195,n13906,n11893 );
   xor U14118 ( n11893,n13573,n14184 );
   nand U14119 ( n14194,p2_reg0_reg_15_,n13549 );
   nand U14120 ( n14193,p2_reg1_reg_15_,n13550 );
   nand U14121 ( n14192,p2_reg2_reg_15_,n13548 );
   or U14122 ( n13784,n13811,n13810 );
   xor U14123 ( n13810,n13726,n11959 );
   not U14124 ( n11959,n10941 );
   nand U14125 ( n10941,n14196,n14197,n14198 );
   nand U14126 ( n14198,n12521,n12612 );
   nand U14127 ( n12612,n14199,n14200 );
   or U14128 ( n14200,p2_ir_reg_16_,p2_ir_reg_31_ );
   nand U14129 ( n14199,p2_ir_reg_31_,n11284 );
   nand U14130 ( n11284,n11293,n14201 );
   nand U14131 ( n14201,p2_ir_reg_16_,n14075 );
   nand U14132 ( n14197,n14057,n14202 );
   nand U14133 ( n14196,n14059,n14203 );
   nand U14134 ( n13811,n14001,n10615 );
   nand U14135 ( n10615,n14204,n14205,n14206,n14207 );
   nand U14136 ( n14207,n13804,n13906 );
   nor U14137 ( n13804,n14208,n14065 );
   and U14138 ( n14208,n13805,n14209 );
   or U14139 ( n14209,n13573,n14184 );
   nand U14140 ( n14206,p2_reg0_reg_16_,n13549 );
   nand U14141 ( n14205,p2_reg1_reg_16_,n13550 );
   nand U14142 ( n14204,p2_reg2_reg_16_,n13548 );
   or U14143 ( n14046,n13632,n13631 );
   nand U14144 ( n14044,n13631,n13632 );
   nand U14145 ( n13632,n14001,n10609 );
   nand U14146 ( n10609,n14210,n14211,n14212,n14213 );
   nand U14147 ( n14213,n13634,n13906 );
   not U14148 ( n13634,n12001 );
   nand U14149 ( n12001,n14214,n14215 );
   nand U14150 ( n14214,n13628,n14216 );
   nand U14151 ( n14216,p2_reg3_reg_17_,n14065 );
   not U14152 ( n13628,p2_reg3_reg_18_ );
   nand U14153 ( n14212,p2_reg0_reg_18_,n13549 );
   nand U14154 ( n14211,p2_reg1_reg_18_,n13550 );
   nand U14155 ( n14210,p2_reg2_reg_18_,n13548 );
   xor U14156 ( n13631,n13726,n12021 );
   not U14157 ( n12021,n10918 );
   nand U14158 ( n10918,n14217,n14218,n14219 );
   nand U14159 ( n14219,n12521,n12550 );
   nand U14160 ( n12550,n14220,n14221,n14222 );
   nand U14161 ( n14221,n11304,n14056 );
   nand U14162 ( n14220,p2_ir_reg_18_,n11303,p2_ir_reg_31_ );
   not U14163 ( n11303,n11302 );
   nand U14164 ( n14218,n14057,n14223 );
   not U14165 ( n14223,n11305 );
   nand U14166 ( n14217,n14059,n14224 );
   nor U14167 ( n13921,n13924,n13926 );
   xor U14168 ( n13926,n13726,n12044 );
   not U14169 ( n12044,n10907 );
   nand U14170 ( n10907,n14225,n14226,n14227 );
   nand U14171 ( n14227,n12521,n11130 );
   nand U14172 ( n14226,n14057,n14228 );
   not U14173 ( n14228,n11312 );
   nand U14174 ( n14225,n14059,n14229 );
   nand U14175 ( n13924,n14001,n10606 );
   nand U14176 ( n10606,n14230,n14231,n14232,n14233 );
   nand U14177 ( n14233,n13906,n13916 );
   xor U14178 ( n13916,p2_reg3_reg_19_,n14234 );
   nand U14179 ( n14232,p2_reg0_reg_19_,n13549 );
   nand U14180 ( n14231,p2_reg1_reg_19_,n13550 );
   nand U14181 ( n14230,p2_reg2_reg_19_,n13548 );
   nand U14182 ( n13715,n14001,n10603,n14235 );
   not U14183 ( n14235,n14040 );
   xor U14184 ( n14040,n13726,n12071 );
   not U14185 ( n12071,n10897 );
   nand U14186 ( n10897,n14236,n14237,n13075 );
   nand U14187 ( n14237,n11416,n14238 );
   or U14188 ( n14236,n11319,n11416 );
   nand U14189 ( n10603,n14239,n14240,n14241,n14242 );
   nand U14190 ( n14242,n13716,n13906 );
   not U14191 ( n13716,n12052 );
   nand U14192 ( n12052,n14243,n14037 );
   nand U14193 ( n14243,n13710,n14244 );
   nand U14194 ( n14244,p2_reg3_reg_19_,n14234 );
   not U14195 ( n13710,p2_reg3_reg_20_ );
   nand U14196 ( n14241,p2_reg0_reg_20_,n13549 );
   nand U14197 ( n14240,p2_reg1_reg_20_,n13550 );
   nand U14198 ( n14239,p2_reg2_reg_20_,n13548 );
   or U14199 ( n14025,n13682,n13681 );
   nand U14200 ( n14023,n13681,n13682 );
   nand U14201 ( n13682,n14001,n10597 );
   nand U14202 ( n10597,n14245,n14246,n14247,n14248 );
   nand U14203 ( n14248,n13684,n13906 );
   not U14204 ( n13684,n12130 );
   nand U14205 ( n12130,n14249,n14250 );
   nand U14206 ( n14249,n13678,n14251 );
   or U14207 ( n14251,n13841,n14037 );
   nand U14208 ( n14247,p2_reg0_reg_22_,n13549 );
   nand U14209 ( n14246,p2_reg1_reg_22_,n13550 );
   nand U14210 ( n14245,p2_reg2_reg_22_,n13548 );
   xor U14211 ( n13681,n13726,n12153 );
   not U14212 ( n12153,n10875 );
   nand U14213 ( n10875,n14252,n14253,n13075 );
   nand U14214 ( n14253,n11416,n14254 );
   or U14215 ( n14252,n11338,n11416 );
   nand U14216 ( n13968,n14001,n10594 );
   nand U14217 ( n10594,n14255,n14256,n14257,n14258 );
   nand U14218 ( n14258,n13906,n12161 );
   xor U14219 ( n12161,p2_reg3_reg_23_,n14259 );
   nand U14220 ( n14257,p2_reg0_reg_23_,n13549 );
   nand U14221 ( n14256,p2_reg1_reg_23_,n13550 );
   nand U14222 ( n14255,p2_reg2_reg_23_,n13548 );
   nand U14223 ( n13765,n14001,n10591,n14260 );
   xor U14224 ( n14260,n13728,n10853 );
   not U14225 ( n10853,n12199 );
   nand U14226 ( n12199,n14261,n14262,n13075 );
   nand U14227 ( n14262,n11416,n14263 );
   or U14228 ( n14261,n11354,n11416 );
   nand U14229 ( n10591,n14264,n14265,n14266,n14267 );
   nand U14230 ( n14267,n12200,n13906 );
   nor U14231 ( n12200,n14268,n14269 );
   and U14232 ( n14268,n13761,n14270 );
   nand U14233 ( n14270,p2_reg3_reg_23_,n14259 );
   nand U14234 ( n14266,p2_reg0_reg_24_,n13549 );
   nand U14235 ( n14265,p2_reg1_reg_24_,n13550 );
   nand U14236 ( n14264,p2_reg2_reg_24_,n13548 );
   and U14237 ( n13603,n13600,n13599 );
   nand U14238 ( n13599,n14271,n14272 );
   nand U14239 ( n14272,n14001,n10585 );
   xor U14240 ( n14271,n13726,n12264 );
   not U14241 ( n12264,n10829 );
   nand U14242 ( n13600,n13822,n13823 );
   nand U14243 ( n13823,n14001,n10588 );
   nand U14244 ( n10588,n14273,n14274,n14275,n14276 );
   nand U14245 ( n14276,n13906,n12217 );
   xor U14246 ( n12217,p2_reg3_reg_25_,n14269 );
   nand U14247 ( n14275,p2_reg0_reg_25_,n13549 );
   nand U14248 ( n14274,p2_reg1_reg_25_,n13550 );
   nand U14249 ( n14273,p2_reg2_reg_25_,n13548 );
   xor U14250 ( n13822,n13726,n12235 );
   not U14251 ( n12235,n10841 );
   nand U14252 ( n10841,n14277,n14278,n13075 );
   nand U14253 ( n14278,n11416,n14279 );
   or U14254 ( n14277,n11364,n11416 );
   and U14255 ( n13598,n14280,n14281 );
   nand U14256 ( n14281,n12436,n13726 );
   nor U14257 ( n12436,n10829,n12288 );
   not U14258 ( n12288,n10585 );
   or U14259 ( n14280,n12257,n13898 );
   nand U14260 ( n13898,n13728,n14001 );
   nand U14261 ( n12257,n10829,n10585 );
   nand U14262 ( n10585,n14282,n14283,n14284,n14285 );
   nand U14263 ( n14285,n13604,n13906 );
   not U14264 ( n13604,n12241 );
   nand U14265 ( n12241,n13908,n14286 );
   nand U14266 ( n14286,n14287,n13590 );
   not U14267 ( n13908,n13996 );
   nand U14268 ( n14284,p2_reg0_reg_26_,n13549 );
   nand U14269 ( n14283,p2_reg1_reg_26_,n13550 );
   nand U14270 ( n14282,p2_reg2_reg_26_,n13548 );
   nand U14271 ( n10829,n14288,n14289,n13075 );
   nand U14272 ( n14289,n11416,n14290 );
   or U14273 ( n14288,n11371,n11416 );
   nand U14274 ( n13984,n12281,n13605 );
   nand U14275 ( n13605,n14291,n14292 );
   nand U14276 ( n14292,n14293,n14294 );
   nand U14277 ( n14294,n14295,n14296 );
   nand U14278 ( n14295,n12526,p2_state_reg );
   xor U14279 ( n12281,p2_reg3_reg_27_,n13996 );
   nor U14280 ( n13996,n13590,n14287 );
   nand U14281 ( n14287,p2_reg3_reg_25_,n14269 );
   nor U14282 ( n14269,n13964,n14250,n13761 );
   not U14283 ( n13761,p2_reg3_reg_24_ );
   not U14284 ( n14250,n14259 );
   nor U14285 ( n14259,n13841,n14037,n13678 );
   not U14286 ( n13678,p2_reg3_reg_22_ );
   nand U14287 ( n14037,p2_reg3_reg_19_,n14234,p2_reg3_reg_20_ );
   not U14288 ( n14234,n14215 );
   nand U14289 ( n14215,p2_reg3_reg_17_,n14065,p2_reg3_reg_18_ );
   nor U14290 ( n14065,n13573,n14184,n13805 );
   not U14291 ( n13805,p2_reg3_reg_16_ );
   nand U14292 ( n14184,p2_reg3_reg_13_,n14095,p2_reg3_reg_14_ );
   not U14293 ( n14095,n14176 );
   nand U14294 ( n14176,p2_reg3_reg_11_,n14148,p2_reg3_reg_12_ );
   nor U14295 ( n14148,n13951,n14297,n13736 );
   not U14296 ( n13736,p2_reg3_reg_9_ );
   not U14297 ( n13951,p2_reg3_reg_10_ );
   not U14298 ( n13573,p2_reg3_reg_15_ );
   not U14299 ( n13841,p2_reg3_reg_21_ );
   not U14300 ( n13964,p2_reg3_reg_23_ );
   not U14301 ( n13590,p2_reg3_reg_26_ );
   nor U14302 ( n14301,n12870,n14302,n14303 );
   nor U14303 ( n14303,n13194,n13589 );
   nor U14304 ( n13574,n14293,n12365,n14296 );
   not U14305 ( n13194,n10645 );
   nor U14306 ( n14302,n11041,n13571 );
   not U14307 ( n13571,n13650 );
   nor U14308 ( n13650,n14293,n12520,n14296 );
   not U14309 ( n11041,n10639 );
   nand U14310 ( n10639,n14304,n14305,n14306,n14307 );
   nand U14311 ( n14307,n14308,n13906 );
   not U14312 ( n14308,n11653 );
   nand U14313 ( n11653,n14309,n14297 );
   not U14314 ( n14297,n14142 );
   nor U14315 ( n14142,n14310,n14311,n13867 );
   nand U14316 ( n14309,n13867,n14312 );
   or U14317 ( n14312,n14310,n14311 );
   not U14318 ( n13867,p2_reg3_reg_8_ );
   nand U14319 ( n14306,p2_reg0_reg_8_,n13549 );
   nand U14320 ( n14305,p2_reg1_reg_8_,n13550 );
   nand U14321 ( n14304,p2_reg2_reg_8_,n13548 );
   nor U14322 ( n12870,p2_state_reg,n14310 );
   nand U14323 ( n14300,n11624,n13581 );
   nand U14324 ( n13581,n14291,n14313 );
   nand U14325 ( n14313,n14314,n14293 );
   nand U14326 ( n14314,n14296,n14315 );
   nand U14327 ( n14315,n11436,n12526 );
   nand U14328 ( n14296,n11436,n13153,n13152 );
   nand U14329 ( n14291,n14316,p2_state_reg );
   nand U14330 ( n14316,n13080,n14317,n12529,n13072 );
   nand U14331 ( n13072,n14318,n13080 );
   nand U14332 ( n12529,n12522,n11137 );
   nand U14333 ( n14317,n14319,n14293 );
   not U14334 ( n14293,n14320 );
   not U14335 ( n13080,n13071 );
   nand U14336 ( n14299,n14321,n14322,n13594 );
   not U14337 ( n13594,n13576 );
   nand U14338 ( n13576,n11436,n14319,n14320 );
   nand U14339 ( n14319,n13361,n11721,n14323,n14324 );
   nor U14340 ( n14324,n14325,n14326 );
   nor U14341 ( n14326,n11142,n13214 );
   nor U14342 ( n14325,n13153,n11669 );
   nand U14343 ( n14323,n11130,n14327 );
   nand U14344 ( n14327,n10790,n11138 );
   not U14345 ( n11138,n13238 );
   nor U14346 ( n13238,n11141,n11131 );
   nor U14347 ( n11672,n14328,n13153 );
   nand U14348 ( n13361,n12349,n11142 );
   nor U14349 ( n12349,n11141,n11130 );
   not U14350 ( n11130,n12525 );
   nand U14351 ( n14322,n14127,n14329 );
   nand U14352 ( n14329,n14128,n14126 );
   and U14353 ( n14127,n13620,n14330 );
   nand U14354 ( n14330,n13616,n13619 );
   not U14355 ( n13616,n14331 );
   nand U14356 ( n14321,n14332,n13619,n14128,n14126 );
   nand U14357 ( n14126,n14333,n14334 );
   nand U14358 ( n14334,n14001,n10642 );
   xor U14359 ( n14333,n11623,n13728 );
   nand U14360 ( n14128,n14001,n10642,n14335 );
   xor U14361 ( n14335,n11623,n13726 );
   nand U14362 ( n10642,n14336,n14337,n14338,n14339 );
   nand U14363 ( n14339,n13906,n11624 );
   xor U14364 ( n11624,n14310,n14311 );
   nand U14365 ( n14311,p2_reg3_reg_6_,n14340 );
   not U14366 ( n14310,p2_reg3_reg_7_ );
   nand U14367 ( n14338,p2_reg0_reg_7_,n13549 );
   nand U14368 ( n14337,p2_reg1_reg_7_,n13550 );
   nand U14369 ( n14336,p2_reg2_reg_7_,n13548 );
   nand U14370 ( n13619,n13617,n13618 );
   nand U14371 ( n14332,n13620,n14331 );
   nand U14372 ( n14331,n14341,n14342 );
   nand U14373 ( n14342,n13794,n14343 );
   or U14374 ( n14343,n13796,n13795 );
   xor U14375 ( n13794,n11582,n13726 );
   not U14376 ( n11582,n11068 );
   nand U14377 ( n11068,n14344,n14345,n14346 );
   nand U14378 ( n14346,n12521,n12913 );
   nand U14379 ( n12913,n14347,n14348,n14349 );
   nand U14380 ( n14348,n14056,n11194 );
   nand U14381 ( n14347,p2_ir_reg_31_,n11184,p2_ir_reg_5_ );
   nand U14382 ( n14345,n14057,n14350 );
   not U14383 ( n14350,n11195 );
   nand U14384 ( n14344,n14059,n14351 );
   nand U14385 ( n14341,n13795,n13796 );
   nand U14386 ( n13796,n14352,n14353 );
   nand U14387 ( n14353,n14354,n13753 );
   nand U14388 ( n13753,n14355,n13940 );
   nand U14389 ( n13940,n14356,n14357 );
   nand U14390 ( n14355,n13942,n13939 );
   or U14391 ( n13939,n14357,n14356 );
   xor U14392 ( n14356,n11520,n13728 );
   not U14393 ( n11520,n11090 );
   nand U14394 ( n11090,n14358,n14359,n14360 );
   nand U14395 ( n14360,n12976,n12521 );
   not U14396 ( n12976,n12972 );
   nand U14397 ( n12972,n14361,n14362 );
   or U14398 ( n14362,p2_ir_reg_31_,p2_ir_reg_3_ );
   or U14399 ( n14361,n11177,n14056 );
   xor U14400 ( n11177,p2_ir_reg_3_,n14363 );
   nand U14401 ( n14359,n14057,n11178 );
   nand U14402 ( n14358,p1_datao_reg_3_,n14059 );
   nand U14403 ( n14357,n10654,n14001 );
   nand U14404 ( n10654,n14364,n14365,n14366,n14367 );
   nand U14405 ( n14367,p2_reg0_reg_3_,n13549 );
   nand U14406 ( n14366,p2_reg1_reg_3_,n13550 );
   nand U14407 ( n14365,p2_reg2_reg_3_,n13548 );
   nand U14408 ( n14364,n13906,n13935 );
   and U14409 ( n13942,n13645,n14368 );
   nand U14410 ( n14368,n13644,n13646 );
   nand U14411 ( n13646,n13648,n13649 );
   not U14412 ( n13644,n13941 );
   nand U14413 ( n13941,n14369,n14370 );
   nand U14414 ( n14370,n13857,n14371 );
   or U14415 ( n14371,n13859,n13858 );
   xor U14416 ( n13857,n11114,n13726 );
   nand U14417 ( n11114,n14372,n14373,n14374 );
   or U14418 ( n14374,n13046,n13075 );
   nand U14419 ( n13046,n14375,n14376 );
   nand U14420 ( n14376,n14377,n14056 );
   or U14421 ( n14375,n11164,n14056 );
   xor U14422 ( n11164,p2_ir_reg_0_,p2_ir_reg_1_ );
   nand U14423 ( n14373,n11165,n14057 );
   nand U14424 ( n14372,p1_datao_reg_1_,n14059 );
   nand U14425 ( n14369,n13858,n13859 );
   nand U14426 ( n13859,n14378,n14379 );
   nand U14427 ( n14379,n13726,n14380 );
   nand U14428 ( n14380,n14381,n13722 );
   or U14429 ( n14378,n13722,n14381 );
   not U14430 ( n14381,n13727 );
   nand U14431 ( n13727,n14001,n10663 );
   nand U14432 ( n10663,n14382,n14383,n14384,n14385 );
   nand U14433 ( n14385,p2_reg0_reg_0_,n13549 );
   nand U14434 ( n14384,p2_reg1_reg_0_,n13550 );
   nand U14435 ( n14383,p2_reg2_reg_0_,n13548 );
   nand U14436 ( n14382,p2_reg3_reg_0_,n13906 );
   xor U14437 ( n13722,n11452,n13726 );
   not U14438 ( n11452,n11125 );
   nand U14439 ( n11125,n14386,n14387,n14388 );
   nand U14440 ( n14388,p2_ir_reg_0_,n12521 );
   nand U14441 ( n14387,n11159,n14057 );
   nand U14442 ( n14386,n14059,p1_datao_reg_0_ );
   nand U14443 ( n13858,n14001,n10660 );
   nand U14444 ( n10660,n14389,n14390,n14391,n14392 );
   nand U14445 ( n14392,p2_reg0_reg_1_,n13549 );
   nand U14446 ( n14391,p2_reg1_reg_1_,n13550 );
   nand U14447 ( n14390,p2_reg2_reg_1_,n13548 );
   nand U14448 ( n14389,p2_reg3_reg_1_,n13906 );
   or U14449 ( n13645,n13649,n13648 );
   xor U14450 ( n13648,n11104,n13726 );
   not U14451 ( n11104,n11490 );
   nand U14452 ( n11490,n14393,n14394,n14395 );
   nand U14453 ( n14395,n12521,n13003 );
   nand U14454 ( n13003,n14396,n14397 );
   or U14455 ( n14397,p2_ir_reg_2_,p2_ir_reg_31_ );
   nand U14456 ( n14396,p2_ir_reg_31_,n11171 );
   nand U14457 ( n11171,n14363,n14398 );
   nand U14458 ( n14398,p2_ir_reg_2_,n14399 );
   nand U14459 ( n14399,n14377,n13047 );
   not U14460 ( n13047,p2_ir_reg_0_ );
   not U14461 ( n14377,p2_ir_reg_1_ );
   nand U14462 ( n14394,n14057,n14400 );
   not U14463 ( n14400,n11172 );
   nand U14464 ( n14393,n14059,n14401 );
   not U14465 ( n14401,p1_datao_reg_2_ );
   nand U14466 ( n13649,n14001,n10657 );
   nand U14467 ( n10657,n14402,n14403,n14404,n14405 );
   nand U14468 ( n14405,p2_reg0_reg_2_,n13549 );
   nand U14469 ( n14404,p2_reg1_reg_2_,n13550 );
   nand U14470 ( n14403,p2_reg2_reg_2_,n13548 );
   nand U14471 ( n14402,p2_reg3_reg_2_,n13906 );
   or U14472 ( n14354,n13752,n13751 );
   nand U14473 ( n14352,n13751,n13752 );
   nand U14474 ( n13752,n14001,n10651 );
   nand U14475 ( n10651,n14406,n14407,n14408,n14409 );
   nand U14476 ( n14409,n11561,n13906 );
   and U14477 ( n11561,n14410,n14411 );
   nand U14478 ( n14410,n13748,n13935 );
   not U14479 ( n13935,p2_reg3_reg_3_ );
   not U14480 ( n13748,p2_reg3_reg_4_ );
   nand U14481 ( n14408,p2_reg0_reg_4_,n13549 );
   nand U14482 ( n14407,p2_reg1_reg_4_,n13550 );
   nand U14483 ( n14406,p2_reg2_reg_4_,n13548 );
   xor U14484 ( n13751,n11080,n13726 );
   not U14485 ( n11080,n11546 );
   nand U14486 ( n11546,n14412,n14413,n14414 );
   nand U14487 ( n14414,n12521,n12979 );
   nand U14488 ( n12979,n14415,n14416 );
   or U14489 ( n14416,p2_ir_reg_31_,p2_ir_reg_4_ );
   nand U14490 ( n14415,p2_ir_reg_31_,n14417 );
   nand U14491 ( n14417,n11184,n11183 );
   nand U14492 ( n11183,p2_ir_reg_4_,n14418 );
   not U14493 ( n11184,n11193 );
   nand U14494 ( n14413,n14057,n14419 );
   not U14495 ( n14419,n11185 );
   nand U14496 ( n14412,n14059,n14420 );
   not U14497 ( n14420,p1_datao_reg_4_ );
   nand U14498 ( n13795,n14001,n10648 );
   nand U14499 ( n10648,n14421,n14422,n14423,n14424 );
   nand U14500 ( n14424,n13906,n11571 );
   xor U14501 ( n11571,n13791,n14411 );
   nand U14502 ( n14423,p2_reg0_reg_5_,n13549 );
   nand U14503 ( n14422,p2_reg1_reg_5_,n13550 );
   nand U14504 ( n14421,p2_reg2_reg_5_,n13548 );
   or U14505 ( n13620,n13618,n13617 );
   xor U14506 ( n13617,n11057,n13726 );
   nand U14507 ( n14425,n14426,n11142 );
   nand U14508 ( n14426,n12348,n13153 );
   nand U14509 ( n11057,n14427,n14428,n14429 );
   nand U14510 ( n14429,n12901,n12521 );
   not U14511 ( n12901,n12918 );
   nand U14512 ( n12918,n14430,n14431 );
   or U14513 ( n14431,p2_ir_reg_31_,p2_ir_reg_6_ );
   nand U14514 ( n14430,p2_ir_reg_31_,n14432 );
   nand U14515 ( n14432,n11200,n11201 );
   nand U14516 ( n11200,p2_ir_reg_6_,n14349 );
   nand U14517 ( n14428,n14057,n11202 );
   nand U14518 ( n14427,p1_datao_reg_6_,n14059 );
   nand U14519 ( n13618,n10645,n14001 );
   not U14520 ( n14328,n13152 );
   nor U14521 ( n13152,n11137,n11142 );
   not U14522 ( n11137,n14433 );
   nor U14523 ( n14433,n11132,n12525 );
   nand U14524 ( n10645,n14434,n14435,n14436,n14437 );
   nand U14525 ( n14437,p2_reg0_reg_6_,n13549 );
   nand U14526 ( n14436,p2_reg1_reg_6_,n13550 );
   nand U14527 ( n14435,p2_reg2_reg_6_,n13548 );
   not U14528 ( n14440,n14439 );
   nand U14529 ( n14434,n13906,n11597 );
   xor U14530 ( n11597,n14340,p2_reg3_reg_6_ );
   nor U14531 ( n14340,n13791,n14411 );
   nand U14532 ( n14411,p2_reg3_reg_4_,p2_reg3_reg_3_ );
   not U14533 ( n13791,p2_reg3_reg_5_ );
   xor U14534 ( n14438,p2_ir_reg_31_,p2_ir_reg_30_ );
   xor U14535 ( n14439,p2_ir_reg_31_,p2_ir_reg_29_ );
   nand U14536 ( n14298,n11042,n13591 );
   nand U14537 ( n13591,n12527,n14441 );
   nand U14538 ( n14441,n11436,n12526,n14320 );
   nor U14539 ( n14320,n10763,n12531,n11134 );
   nand U14540 ( n11134,n11147,n14442 );
   or U14541 ( n14442,n11437,p2_d_reg_1_ );
   nand U14542 ( n11147,n14443,n14444 );
   nor U14543 ( n12531,n11437,n14445 );
   and U14544 ( n14445,n14446,n14447,n14448,n14449 );
   nor U14545 ( n14449,n14450,n14451,n14452,n14453 );
   nand U14546 ( n14453,n11430,n11431,n11429 );
   not U14547 ( n11429,p2_d_reg_25_ );
   not U14548 ( n11431,p2_d_reg_27_ );
   not U14549 ( n11430,p2_d_reg_26_ );
   nand U14550 ( n14452,n11432,n11433,n11417,n11434 );
   not U14551 ( n11434,p2_d_reg_30_ );
   not U14552 ( n11417,p2_d_reg_2_ );
   not U14553 ( n11433,p2_d_reg_29_ );
   not U14554 ( n11432,p2_d_reg_28_ );
   nand U14555 ( n14451,n11435,n11418,n11419,n11420 );
   not U14556 ( n11420,p2_d_reg_5_ );
   not U14557 ( n11419,p2_d_reg_4_ );
   not U14558 ( n11418,p2_d_reg_3_ );
   not U14559 ( n11435,p2_d_reg_31_ );
   nand U14560 ( n14450,n11421,n11422,n11423,n11424 );
   not U14561 ( n11424,p2_d_reg_9_ );
   not U14562 ( n11423,p2_d_reg_8_ );
   not U14563 ( n11422,p2_d_reg_7_ );
   not U14564 ( n11421,p2_d_reg_6_ );
   nor U14565 ( n14448,n14454,p2_d_reg_10_,p2_d_reg_12_,p2_d_reg_11_ );
   nand U14566 ( n14454,n11425,n11426,n11427,n11428 );
   not U14567 ( n11428,p2_d_reg_16_ );
   not U14568 ( n11427,p2_d_reg_15_ );
   not U14569 ( n11426,p2_d_reg_14_ );
   not U14570 ( n11425,p2_d_reg_13_ );
   nor U14571 ( n14447,p2_d_reg_24_,p2_d_reg_23_,p2_d_reg_22_,p2_d_reg_21_ );
   nor U14572 ( n14446,p2_d_reg_20_,p2_d_reg_19_,p2_d_reg_18_,p2_d_reg_17_ );
   nand U14573 ( n10763,n11150,n14455 );
   or U14574 ( n14455,n11437,p2_d_reg_0_ );
   nand U14575 ( n11437,n14456,n14457 );
   nand U14576 ( n14457,n14458,n14444 );
   xor U14577 ( n14458,n12519,n14459 );
   not U14578 ( n12519,p2_b_reg );
   nand U14579 ( n11150,n14443,n14459 );
   nand U14580 ( n12526,n11128,n14460 );
   nand U14581 ( n14460,n11127,n11132 );
   nor U14582 ( n11127,n13214,n11131 );
   nand U14583 ( n13214,n12525,n11141 );
   nand U14584 ( n11128,n11142,n11141,n13209 );
   nor U14585 ( n13209,n12525,n12348 );
   not U14586 ( n12348,n11132 );
   nand U14587 ( n12527,n11436,n12525,n10773 );
   nor U14588 ( n10773,n11131,n13153,n11132 );
   nand U14589 ( n11132,n14461,n14462 );
   nand U14590 ( n14462,p2_ir_reg_20_,n14056 );
   nand U14591 ( n14461,n11317,n11318,p2_ir_reg_31_ );
   nand U14592 ( n11317,p2_ir_reg_20_,n11311 );
   not U14593 ( n13153,n11141 );
   not U14594 ( n11131,n11142 );
   nand U14595 ( n12525,n14463,n14464 );
   nand U14596 ( n14464,p2_ir_reg_19_,n14056 );
   nand U14597 ( n14463,n11310,n11311,p2_ir_reg_31_ );
   nand U14598 ( n11310,p2_ir_reg_19_,n14222 );
   nor U14599 ( n11436,n14318,p2_u3152,n13071 );
   not U14600 ( n11042,n11623 );
   nand U14601 ( n11623,n14465,n14466,n14467 );
   nand U14602 ( n14467,n12521,n12853 );
   nand U14603 ( n12853,n14468,n14469,n14135 );
   nand U14604 ( n14469,n14056,n11210 );
   nand U14605 ( n14468,p2_ir_reg_31_,n11201,p2_ir_reg_7_ );
   not U14606 ( n11201,n11209 );
   nand U14607 ( n14466,n14057,n14470 );
   not U14608 ( n14470,n11211 );
   nand U14609 ( n14465,n14059,n14471 );
   not U14610 ( n14471,p1_datao_reg_7_ );
   nor U14611 ( n12522,n11142,n11141 );
   nand U14612 ( n11141,n14473,n14474,n11336 );
   nand U14613 ( n14474,n11327,n14056 );
   nand U14614 ( n14473,p2_ir_reg_21_,n11318,p2_ir_reg_31_ );
   nand U14615 ( n11142,n14475,n14476,n14477 );
   nand U14616 ( n14476,n11337,n14056 );
   nand U14617 ( n14475,p2_ir_reg_22_,n11336,p2_ir_reg_31_ );
   not U14618 ( n11336,n11335 );
   nor U14619 ( n14318,n14443,n14459,n14444 );
   nand U14620 ( n14444,n14478,n14479,n14480 );
   nand U14621 ( n14479,n11363,n14056 );
   nand U14622 ( n14478,p2_ir_reg_25_,n11362,p2_ir_reg_31_ );
   xor U14623 ( n14459,n14481,n11353 );
   not U14624 ( n11353,p2_ir_reg_24_ );
   nor U14625 ( n14481,n11352,n14056 );
   not U14626 ( n14443,n14456 );
   nand U14627 ( n14456,n14482,n14483 );
   nand U14628 ( n14483,p2_ir_reg_26_,n14056 );
   nand U14629 ( n14482,n11369,n11370,p2_ir_reg_31_ );
   nand U14630 ( n11370,p2_ir_reg_26_,n14480 );
   and U14631 ( n13074,n14484,p2_state_reg );
   nand U14632 ( n14484,n13071,n13075 );
   not U14633 ( n13075,n12521 );
   not U14634 ( n13068,n13065 );
   nand U14635 ( n13065,n14485,n14486,n11388 );
   nand U14636 ( n14486,n11379,n14056 );
   not U14637 ( n11379,p2_ir_reg_27_ );
   nand U14638 ( n14485,p2_ir_reg_27_,n11369,p2_ir_reg_31_ );
   not U14639 ( n12520,n12365 );
   nand U14640 ( n12365,n14487,n14488,n11398 );
   not U14641 ( n11398,n11397 );
   nor U14642 ( n11397,n11388,p2_ir_reg_28_ );
   nand U14643 ( n14488,n11389,n14056 );
   not U14644 ( n11389,p2_ir_reg_28_ );
   nand U14645 ( n14487,p2_ir_reg_28_,n11388,p2_ir_reg_31_ );
   not U14646 ( n11388,n11387 );
   nor U14647 ( n11387,n11369,p2_ir_reg_27_ );
   not U14648 ( n11369,n11378 );
   nor U14649 ( n11378,n14480,p2_ir_reg_26_ );
   nand U14650 ( n14480,n11361,n11363 );
   not U14651 ( n11363,p2_ir_reg_25_ );
   not U14652 ( n11361,n11362 );
   nand U14653 ( n11362,n14489,n11327,n14490,n14491 );
   nor U14654 ( n14491,p2_ir_reg_19_,p2_ir_reg_18_,p2_ir_reg_17_,n11293 );
   nor U14655 ( n14490,p2_ir_reg_22_,p2_ir_reg_24_,p2_ir_reg_23_ );
   not U14656 ( n11327,p2_ir_reg_21_ );
   not U14657 ( n14489,p2_ir_reg_20_ );
   nand U14658 ( n13071,n14492,n14493 );
   nand U14659 ( n14493,p2_ir_reg_23_,n14056 );
   not U14660 ( n14056,p2_ir_reg_31_ );
   nand U14661 ( n14492,n11343,n11344,p2_ir_reg_31_ );
   nand U14662 ( n11344,p2_ir_reg_23_,n14477 );
   not U14663 ( n11343,n11352 );
   nor U14664 ( n11352,n14477,p2_ir_reg_23_ );
   nand U14665 ( n14477,n11335,n11337 );
   not U14666 ( n11337,p2_ir_reg_22_ );
   nor U14667 ( n11335,n11318,p2_ir_reg_21_ );
   not U14668 ( n11318,n11326 );
   nor U14669 ( n11326,n11311,p2_ir_reg_20_ );
   or U14670 ( n11311,n14222,p2_ir_reg_19_ );
   nand U14671 ( n14222,n11302,n11304 );
   not U14672 ( n11304,p2_ir_reg_18_ );
   nor U14673 ( n11302,n11293,p2_ir_reg_17_ );
   not U14674 ( n11293,n11292 );
   nor U14675 ( n11292,n14075,p2_ir_reg_16_ );
   nand U14676 ( n14075,n11275,n11277 );
   not U14677 ( n11277,p2_ir_reg_15_ );
   nor U14678 ( n11275,n14090,p2_ir_reg_14_ );
   nand U14679 ( n14090,n11258,n11260 );
   not U14680 ( n11260,p2_ir_reg_13_ );
   nor U14681 ( n11258,n14155,p2_ir_reg_12_ );
   nand U14682 ( n14155,n11241,n11243 );
   not U14683 ( n11243,p2_ir_reg_11_ );
   nor U14684 ( n11241,n14111,p2_ir_reg_10_ );
   nand U14685 ( n14111,n11225,n11226 );
   not U14686 ( n11226,p2_ir_reg_9_ );
   nor U14687 ( n11225,n14135,p2_ir_reg_8_ );
   nand U14688 ( n14135,n11209,n11210 );
   not U14689 ( n11210,p2_ir_reg_7_ );
   nor U14690 ( n11209,n14349,p2_ir_reg_6_ );
   nand U14691 ( n14349,n11193,n11194 );
   not U14692 ( n11194,p2_ir_reg_5_ );
   nor U14693 ( n11193,n14418,p2_ir_reg_4_ );
   or U14694 ( n14418,n14363,p2_ir_reg_3_ );
   or U14695 ( n14363,p2_ir_reg_1_,p2_ir_reg_2_,p2_ir_reg_0_ );
   nand U14696 ( n14494,p1_u4006,n14497 );
   nand U14697 ( n14498,p1_u4006,n14500 );
   nand U14698 ( n14501,p1_u4006,n14503 );
   nand U14699 ( n14504,p1_u4006,n14506 );
   nand U14700 ( n14507,p1_u4006,n14509 );
   nand U14701 ( n14510,p1_u4006,n14512 );
   nand U14702 ( n14513,p1_u4006,n14515 );
   nand U14703 ( n14516,p1_u4006,n14518 );
   nand U14704 ( n14519,p1_u4006,n14521 );
   nand U14705 ( n14522,p1_u4006,n14524 );
   nand U14706 ( n14525,p1_u4006,n14527 );
   nand U14707 ( n14528,p1_u4006,n14530 );
   nand U14708 ( n14531,p1_u4006,n14533 );
   nand U14709 ( n14534,p1_u4006,n14536 );
   nand U14710 ( n14537,p1_u4006,n14539 );
   nand U14711 ( n14540,p1_u4006,n14542 );
   nand U14712 ( n14543,p1_u4006,n14545 );
   nand U14713 ( n14546,p1_u4006,n14548 );
   nand U14714 ( n14549,p1_u4006,n14551 );
   nand U14715 ( n14552,p1_u4006,n14554 );
   nand U14716 ( n14555,p1_u4006,n14557 );
   nand U14717 ( n14558,p1_u4006,n14560 );
   nand U14718 ( n14561,p1_u4006,n14563 );
   nand U14719 ( n14564,p1_u4006,n14566 );
   nand U14720 ( n14567,p1_u4006,n14569 );
   nand U14721 ( n14570,p1_u4006,n14572 );
   nand U14722 ( n14573,p1_u4006,n14575 );
   nand U14723 ( n14576,p1_u4006,n14578 );
   nand U14724 ( n14579,p1_u4006,n14581 );
   nand U14725 ( n14582,p1_u4006,n14584 );
   nand U14726 ( n14585,p1_u4006,n14587 );
   nand U14727 ( n14588,p1_u4006,n14590 );
   nand U14728 ( n14591,p1_reg1_reg_31_,n14595 );
   nand U14729 ( n14597,p1_reg1_reg_30_,n14595 );
   nand U14730 ( n14596,n14593,n14598 );
   nand U14731 ( n14600,p1_reg1_reg_29_,n14595 );
   nand U14732 ( n14599,n14593,n14601 );
   nand U14733 ( n14603,p1_reg1_reg_28_,n14595 );
   nand U14734 ( n14602,n14593,n14604 );
   nand U14735 ( n14606,p1_reg1_reg_27_,n14595 );
   nand U14736 ( n14605,n14593,n14607 );
   nand U14737 ( n14609,p1_reg1_reg_26_,n14595 );
   nand U14738 ( n14608,n14593,n14610 );
   nand U14739 ( n14612,p1_reg1_reg_25_,n14595 );
   nand U14740 ( n14611,n14593,n14613 );
   nand U14741 ( n14615,p1_reg1_reg_24_,n14595 );
   nand U14742 ( n14614,n14593,n14616 );
   nand U14743 ( n14618,p1_reg1_reg_23_,n14595 );
   nand U14744 ( n14617,n14593,n14619 );
   nand U14745 ( n14621,p1_reg1_reg_22_,n14595 );
   nand U14746 ( n14620,n14593,n14622 );
   nand U14747 ( n14624,p1_reg1_reg_21_,n14595 );
   nand U14748 ( n14623,n14593,n14625 );
   nand U14749 ( n14627,p1_reg1_reg_20_,n14595 );
   nand U14750 ( n14626,n14593,n14628 );
   nand U14751 ( n14630,p1_reg1_reg_19_,n14595 );
   nand U14752 ( n14629,n14593,n14631 );
   nand U14753 ( n14633,p1_reg1_reg_18_,n14595 );
   nand U14754 ( n14632,n14593,n14634 );
   nand U14755 ( n14636,p1_reg1_reg_17_,n14595 );
   nand U14756 ( n14635,n14593,n14637 );
   nand U14757 ( n14639,p1_reg1_reg_16_,n14595 );
   nand U14758 ( n14638,n14593,n14640 );
   nand U14759 ( n14642,p1_reg1_reg_15_,n14595 );
   nand U14760 ( n14641,n14593,n14643 );
   nand U14761 ( n14645,p1_reg1_reg_14_,n14595 );
   nand U14762 ( n14644,n14593,n14646 );
   nand U14763 ( n14648,p1_reg1_reg_13_,n14595 );
   nand U14764 ( n14647,n14593,n14649 );
   nand U14765 ( n14651,p1_reg1_reg_12_,n14595 );
   nand U14766 ( n14650,n14593,n14652 );
   nand U14767 ( n14654,p1_reg1_reg_11_,n14595 );
   nand U14768 ( n14653,n14593,n14655 );
   nand U14769 ( n14657,p1_reg1_reg_10_,n14595 );
   nand U14770 ( n14656,n14593,n14658 );
   nand U14771 ( n14660,p1_reg1_reg_9_,n14595 );
   nand U14772 ( n14659,n14593,n14661 );
   nand U14773 ( n14663,p1_reg1_reg_8_,n14595 );
   nand U14774 ( n14662,n14593,n14664 );
   nand U14775 ( n14666,p1_reg1_reg_7_,n14595 );
   nand U14776 ( n14665,n14593,n14667 );
   nand U14777 ( n14669,p1_reg1_reg_6_,n14595 );
   nand U14778 ( n14668,n14593,n14670 );
   nand U14779 ( n14672,p1_reg1_reg_5_,n14595 );
   nand U14780 ( n14671,n14593,n14673 );
   nand U14781 ( n14675,p1_reg1_reg_4_,n14595 );
   nand U14782 ( n14674,n14593,n14676 );
   nand U14783 ( n14678,p1_reg1_reg_3_,n14595 );
   nand U14784 ( n14677,n14593,n14679 );
   nand U14785 ( n14681,p1_reg1_reg_2_,n14595 );
   nand U14786 ( n14680,n14593,n14682 );
   nand U14787 ( n14684,p1_reg1_reg_1_,n14595 );
   nand U14788 ( n14683,n14593,n14685 );
   nand U14789 ( n14687,p1_reg1_reg_0_,n14595 );
   nand U14790 ( n14686,n14593,n14688 );
   nand U14791 ( n14594,n14694,n14695,n14696 );
   nand U14792 ( n14696,n14697,n14698 );
   nand U14793 ( n14694,n14699,n14700 );
   nand U14794 ( n14691,p1_reg0_reg_31_,n14701 );
   nand U14795 ( n14598,n14704,n14695,n14705 );
   nand U14796 ( n14705,n14706,n14698 );
   not U14797 ( n14695,n14707 );
   nand U14798 ( n14704,n14708,n14709,n14699 );
   nand U14799 ( n14702,p1_reg0_reg_30_,n14701 );
   nand U14800 ( n14601,n14712,n14713,n14714,n14715 );
   nand U14801 ( n14715,n14699,n14716 );
   nand U14802 ( n14714,n14717,n14718 );
   nand U14803 ( n14713,n14719,n14698 );
   not U14804 ( n14712,n14720 );
   nand U14805 ( n14710,p1_reg0_reg_29_,n14701 );
   nand U14806 ( n14604,n14723,n14724,n14725 );
   nor U14807 ( n14725,n14726,n14727,n14728 );
   nor U14808 ( n14728,n14729,n14730 );
   and U14809 ( n14727,n14699,n14731 );
   nor U14810 ( n14726,n14732,n14733 );
   nand U14811 ( n14724,n14734,n14698 );
   nand U14812 ( n14721,p1_reg0_reg_28_,n14701 );
   nand U14813 ( n14607,n14737,n14738,n14739 );
   nor U14814 ( n14739,n14740,n14741,n14742 );
   nor U14815 ( n14742,n14729,n14743 );
   and U14816 ( n14741,n14744,n14699 );
   nor U14817 ( n14740,n14745,n14733 );
   nand U14818 ( n14738,n14746,n14698 );
   nand U14819 ( n14735,p1_reg0_reg_27_,n14701 );
   nand U14820 ( n14610,n14749,n14750,n14751 );
   nor U14821 ( n14751,n14752,n14753,n14754 );
   nor U14822 ( n14754,n14729,n14755 );
   nor U14823 ( n14753,n14756,n14757 );
   nor U14824 ( n14752,n14758,n14733 );
   nand U14825 ( n14750,n14759,n14698 );
   nand U14826 ( n14747,p1_reg0_reg_26_,n14701 );
   nand U14827 ( n14613,n14762,n14763,n14764,n14765 );
   nand U14828 ( n14765,n14766,n14512 );
   nor U14829 ( n14764,n14767,n14768 );
   nor U14830 ( n14768,n14769,n14729 );
   and U14831 ( n14767,n14770,n14699 );
   nand U14832 ( n14763,n14771,n14698 );
   nand U14833 ( n14760,p1_reg0_reg_25_,n14701 );
   nand U14834 ( n14616,n14774,n14775,n14776,n14777 );
   nand U14835 ( n14777,n14766,n14515 );
   nor U14836 ( n14776,n14778,n14779 );
   nor U14837 ( n14779,n14780,n14729 );
   nor U14838 ( n14778,n14756,n14781 );
   nand U14839 ( n14775,n14782,n14698 );
   nand U14840 ( n14772,p1_reg0_reg_24_,n14701 );
   nand U14841 ( n14619,n14785,n14786,n14787 );
   nor U14842 ( n14787,n14788,n14789,n14790 );
   nor U14843 ( n14790,n14791,n14729 );
   and U14844 ( n14789,n14792,n14699 );
   nor U14845 ( n14788,n14793,n14733 );
   nand U14846 ( n14786,n14794,n14698 );
   nand U14847 ( n14783,p1_reg0_reg_23_,n14701 );
   nand U14848 ( n14622,n14797,n14798,n14799,n14800 );
   nor U14849 ( n14800,n14801,n14802 );
   nor U14850 ( n14801,n14803,n14804 );
   nand U14851 ( n14799,n14766,n14521 );
   nand U14852 ( n14798,n14805,n14806 );
   nand U14853 ( n14797,n14807,n14699 );
   nand U14854 ( n14795,p1_reg0_reg_22_,n14701 );
   nand U14855 ( n14625,n14810,n14811,n14812 );
   nor U14856 ( n14812,n14813,n14814,n14815 );
   nor U14857 ( n14815,n14729,n14816 );
   and U14858 ( n14814,n14817,n14699 );
   nor U14859 ( n14813,n14818,n14733 );
   nand U14860 ( n14811,n14819,n14698 );
   nand U14861 ( n14808,p1_reg0_reg_21_,n14701 );
   nand U14862 ( n14628,n14822,n14823,n14824,n14825 );
   nor U14863 ( n14825,n14826,n14827 );
   nor U14864 ( n14826,n14803,n14828 );
   nand U14865 ( n14824,n14766,n14527 );
   nand U14866 ( n14823,n14829,n14699 );
   nand U14867 ( n14822,n14830,n14717 );
   nand U14868 ( n14820,p1_reg0_reg_20_,n14701 );
   nand U14869 ( n14631,n14833,n14834,n14835,n14836 );
   nor U14870 ( n14836,n14837,n14838 );
   nor U14871 ( n14837,n14803,n14839 );
   nand U14872 ( n14835,n14766,n14530 );
   nand U14873 ( n14834,n14699,n14840 );
   nand U14874 ( n14833,n14841,n14717 );
   nand U14875 ( n14831,p1_reg0_reg_19_,n14701 );
   nand U14876 ( n14634,n14844,n14845,n14846,n14847 );
   nor U14877 ( n14847,n14848,n14849 );
   nor U14878 ( n14848,n14803,n14850 );
   nand U14879 ( n14846,n14766,n14533 );
   nand U14880 ( n14845,n14851,n14806 );
   nand U14881 ( n14844,n14852,n14699 );
   nand U14882 ( n14842,p1_reg0_reg_18_,n14701 );
   nand U14883 ( n14637,n14855,n14856,n14857 );
   nor U14884 ( n14857,n14858,n14859,n14860 );
   nor U14885 ( n14860,n14729,n14861 );
   and U14886 ( n14859,n14862,n14699 );
   nor U14887 ( n14858,n14863,n14733 );
   nand U14888 ( n14856,n14864,n14698 );
   nand U14889 ( n14853,p1_reg0_reg_17_,n14701 );
   nand U14890 ( n14640,n14867,n14868,n14869,n14870 );
   nand U14891 ( n14870,n14766,n14539 );
   nor U14892 ( n14869,n14871,n14872 );
   nor U14893 ( n14872,n14873,n14729 );
   nor U14894 ( n14871,n14756,n14874 );
   nand U14895 ( n14868,n14875,n14698 );
   nand U14896 ( n14865,p1_reg0_reg_16_,n14701 );
   nand U14897 ( n14643,n14878,n14879,n14880,n14881 );
   nor U14898 ( n14881,n14882,n14883 );
   nor U14899 ( n14882,n14803,n14884 );
   nand U14900 ( n14880,n14766,n14542 );
   nand U14901 ( n14879,n14699,n14885 );
   nand U14902 ( n14878,n14886,n14806 );
   nand U14903 ( n14876,p1_reg0_reg_15_,n14701 );
   nand U14904 ( n14646,n14889,n14890,n14891,n14892 );
   nor U14905 ( n14892,n14893,n14894 );
   nor U14906 ( n14893,n14803,n14895 );
   nand U14907 ( n14891,n14766,n14545 );
   nand U14908 ( n14890,n14896,n14806 );
   nand U14909 ( n14889,n14897,n14699 );
   nand U14910 ( n14887,p1_reg0_reg_14_,n14701 );
   nand U14911 ( n14649,n14900,n14901,n14902 );
   nor U14912 ( n14902,n14903,n14904,n14905 );
   nor U14913 ( n14905,n14729,n14906 );
   and U14914 ( n14904,n14907,n14699 );
   nor U14915 ( n14903,n14908,n14733 );
   nand U14916 ( n14901,n14909,n14698 );
   nand U14917 ( n14898,p1_reg0_reg_13_,n14701 );
   nand U14918 ( n14652,n14912,n14913,n14914,n14915 );
   nor U14919 ( n14915,n14916,n14917 );
   nor U14920 ( n14916,n14803,n14918 );
   nand U14921 ( n14914,n14766,n14551 );
   nand U14922 ( n14913,n14919,n14806 );
   nand U14923 ( n14912,n14920,n14699 );
   nand U14924 ( n14910,p1_reg0_reg_12_,n14701 );
   nand U14925 ( n14655,n14923,n14924,n14925 );
   nor U14926 ( n14925,n14926,n14927,n14928 );
   nor U14927 ( n14928,n14729,n14929 );
   and U14928 ( n14927,n14930,n14699 );
   nor U14929 ( n14926,n14931,n14733 );
   nand U14930 ( n14924,n14932,n14698 );
   nand U14931 ( n14921,p1_reg0_reg_11_,n14701 );
   nand U14932 ( n14658,n14935,n14936,n14937,n14938 );
   nor U14933 ( n14938,n14939,n14940 );
   nor U14934 ( n14939,n14803,n14941 );
   nand U14935 ( n14937,n14766,n14557 );
   nand U14936 ( n14936,n14942,n14699 );
   nand U14937 ( n14935,n14943,n14717 );
   nand U14938 ( n14933,p1_reg0_reg_10_,n14701 );
   nand U14939 ( n14661,n14946,n14947,n14948,n14949 );
   nor U14940 ( n14949,n14950,n14951 );
   nor U14941 ( n14950,n14803,n14952 );
   nand U14942 ( n14948,n14766,n14560 );
   nand U14943 ( n14947,n14699,n14953 );
   nand U14944 ( n14946,n14954,n14806 );
   nand U14945 ( n14944,p1_reg0_reg_9_,n14701 );
   nand U14946 ( n14664,n14957,n14958,n14959 );
   nor U14947 ( n14959,n14960,n14961,n14962 );
   nor U14948 ( n14962,n14729,n14963 );
   nor U14949 ( n14961,n14756,n14964 );
   nor U14950 ( n14960,n14965,n14733 );
   nand U14951 ( n14958,n14966,n14698 );
   nand U14952 ( n14955,p1_reg0_reg_8_,n14701 );
   nand U14953 ( n14667,n14969,n14970,n14971 );
   nor U14954 ( n14971,n14972,n14973,n14974 );
   nor U14955 ( n14974,n14729,n14975 );
   and U14956 ( n14973,n14976,n14699 );
   nor U14957 ( n14972,n14977,n14733 );
   nand U14958 ( n14970,n14978,n14698 );
   nand U14959 ( n14967,p1_reg0_reg_7_,n14701 );
   nand U14960 ( n14670,n14981,n14982,n14983 );
   nor U14961 ( n14983,n14984,n14985,n14986 );
   nor U14962 ( n14986,n14729,n14987 );
   nor U14963 ( n14985,n14756,n14988 );
   nor U14964 ( n14984,n14989,n14733 );
   nand U14965 ( n14982,n14990,n14698 );
   nand U14966 ( n14979,p1_reg0_reg_6_,n14701 );
   nand U14967 ( n14673,n14993,n14994,n14995 );
   nor U14968 ( n14995,n14996,n14997,n14998 );
   nor U14969 ( n14998,n14999,n14729 );
   and U14970 ( n14997,n15000,n14699 );
   nor U14971 ( n14996,n15001,n14733 );
   nand U14972 ( n14994,n15002,n14698 );
   nand U14973 ( n14991,p1_reg0_reg_5_,n14701 );
   nand U14974 ( n14676,n15005,n15006,n15007,n15008 );
   nor U14975 ( n15008,n15009,n15010 );
   nor U14976 ( n15009,n14803,n15011 );
   nand U14977 ( n15007,n14766,n14575 );
   nand U14978 ( n15006,n15012,n14806 );
   nand U14979 ( n15005,n15013,n14699 );
   nand U14980 ( n15003,p1_reg0_reg_4_,n14701 );
   nand U14981 ( n14679,n15016,n15017,n15018,n15019 );
   nor U14982 ( n15019,n15020,n15021 );
   nor U14983 ( n15020,n14803,n15022 );
   nand U14984 ( n15018,n14766,n14578 );
   nand U14985 ( n15017,n14699,n15023 );
   nand U14986 ( n15016,n15024,n14806 );
   nand U14987 ( n15014,p1_reg0_reg_3_,n14701 );
   nand U14988 ( n14682,n15027,n15028,n15029,n15030 );
   nand U14989 ( n15030,n14766,n14581 );
   nor U14990 ( n15029,n15031,n15032 );
   nor U14991 ( n15032,n14756,n15033 );
   nor U14992 ( n15031,n15034,n15035 );
   nand U14993 ( n15028,n15036,n14698 );
   nand U14994 ( n15025,p1_reg0_reg_2_,n14701 );
   nand U14995 ( n14685,n15039,n15040,n15041,n15042 );
   nor U14996 ( n15042,n15043,n15044 );
   nor U14997 ( n15043,n14803,n15045 );
   nand U14998 ( n15041,n14766,n14584 );
   nand U14999 ( n15040,n14699,n15046 );
   nand U15000 ( n15039,n15047,n14806 );
   not U15001 ( n14806,n15034 );
   nor U15002 ( n15034,n15048,n14717 );
   nand U15003 ( n15037,p1_reg0_reg_1_,n14701 );
   nand U15004 ( n14688,n15051,n15052,n15053,n15054 );
   nand U15005 ( n15054,n15055,n15056 );
   nand U15006 ( n15055,n14803,n14756 );
   nand U15007 ( n15053,n14766,n14587 );
   nand U15008 ( n15052,n15057,n14717 );
   not U15009 ( n15051,n15058 );
   nand U15010 ( n15049,p1_reg0_reg_0_,n14701 );
   and U15011 ( n14690,n15060,n15061,n15062 );
   nor U15012 ( n15062,n15063,n15064,n15065 );
   nor U15013 ( n15063,n15066,n14756 );
   nand U15014 ( n15067,n15070,n15071 );
   nand U15015 ( n15072,n15070,n15074 );
   and U15016 ( n15081,n14716,n15082 );
   xor U15017 ( n14716,n15083,n15084 );
   and U15018 ( n15080,n15085,n15086 );
   and U15019 ( n15079,n14718,n15087 );
   nand U15020 ( n15077,n15088,n14719 );
   nand U15021 ( n15076,p1_reg2_reg_29_,n15089 );
   nand U15022 ( n15075,n15090,n14720 );
   nand U15023 ( n14720,n15091,n15092,n15093,n15094 );
   nand U15024 ( n15094,n15095,n15096 );
   nand U15025 ( n15096,n15097,n15098,n15099 );
   not U15026 ( n15099,n15100 );
   nand U15027 ( n15098,n15101,n15102,n15103 );
   or U15028 ( n15097,n15101,n15104,n15103 );
   nor U15029 ( n15093,n15105,n15106 );
   nor U15030 ( n15106,n15107,n15108 );
   nor U15031 ( n15105,n15109,n15110 );
   nor U15032 ( n15110,n15100,n15111,n15112 );
   nor U15033 ( n15112,n15103,n15104,n15113 );
   and U15034 ( n15111,n15103,n15102,n15113 );
   nand U15035 ( n15100,n15114,n15115 );
   nand U15036 ( n15115,n15104,n15103 );
   or U15037 ( n15114,n15102,n15103 );
   nand U15038 ( n15092,n14718,n15048 );
   xor U15039 ( n14718,n15116,n15117 );
   nand U15040 ( n15117,n15118,n15119 );
   nand U15041 ( n15119,n14745,n15120 );
   nand U15042 ( n15120,n14734,n15121 );
   or U15043 ( n15118,n15121,n14734 );
   nand U15044 ( n15091,n15122,n14506 );
   nand U15045 ( n15125,n15126,n11159 );
   or U15046 ( n15127,n15128,n15129 );
   nand U15047 ( n15123,n15130,p2_datao_reg_0_ );
   nand U15048 ( n15134,n15129,n15135 );
   nand U15049 ( n15133,n15130,p2_datao_reg_1_ );
   nand U15050 ( n15132,n15128,p1_ir_reg_1_ );
   nand U15051 ( n15131,n15126,n11165 );
   nand U15052 ( n15139,n15140,n15141,n15129 );
   nand U15053 ( n15138,n15130,p2_datao_reg_2_ );
   nand U15054 ( n15137,n15128,p1_ir_reg_2_ );
   nand U15055 ( n15136,n15126,n11172 );
   nand U15056 ( n15145,n15146,n15129 );
   nand U15057 ( n15144,n15130,p2_datao_reg_3_ );
   nand U15058 ( n15143,n15128,p1_ir_reg_3_ );
   nand U15059 ( n15142,n15126,n11178 );
   nand U15060 ( n15150,n15151,n15152,n15129 );
   nand U15061 ( n15149,n15130,p2_datao_reg_4_ );
   nand U15062 ( n15148,n15128,p1_ir_reg_4_ );
   nand U15063 ( n15147,n15126,n11185 );
   nand U15064 ( n15156,p1_ir_reg_5_,n15157 );
   nand U15065 ( n15157,n15158,n15159 );
   nand U15066 ( n15159,n15129,n15160 );
   nand U15067 ( n15155,n15129,n15152,n15161 );
   nand U15068 ( n15154,n15130,p2_datao_reg_5_ );
   nand U15069 ( n15153,n15126,n11195 );
   nand U15070 ( n15165,n15166,n15167,n15129 );
   nand U15071 ( n15164,n15130,p2_datao_reg_6_ );
   nand U15072 ( n15163,n15128,p1_ir_reg_6_ );
   nand U15073 ( n15162,n15126,n11202 );
   nand U15074 ( n15171,p1_ir_reg_7_,n15172 );
   nand U15075 ( n15172,n15158,n15173 );
   nand U15076 ( n15173,n15129,n15174 );
   nand U15077 ( n15170,n15129,n15167,n15175 );
   nand U15078 ( n15169,n15130,p2_datao_reg_7_ );
   nand U15079 ( n15168,n15126,n11211 );
   nand U15080 ( n15179,n15180,n15181,n15129 );
   nand U15081 ( n15178,n15130,p2_datao_reg_8_ );
   nand U15082 ( n15177,n15128,p1_ir_reg_8_ );
   nand U15083 ( n15176,n15126,n11218 );
   nand U15084 ( n15185,n15186,n15129 );
   nand U15085 ( n15184,n15130,p2_datao_reg_9_ );
   nand U15086 ( n15183,n15128,p1_ir_reg_9_ );
   nand U15087 ( n15182,n15126,n11227 );
   nand U15088 ( n15190,n15191,n15129 );
   not U15089 ( n15191,n15192 );
   nand U15090 ( n15189,n15130,p2_datao_reg_10_ );
   nand U15091 ( n15188,n15128,p1_ir_reg_10_ );
   nand U15092 ( n15187,n15126,n11234 );
   nand U15093 ( n15196,n15197,n15129 );
   nand U15094 ( n15195,n15130,p2_datao_reg_11_ );
   nand U15095 ( n15194,n15128,p1_ir_reg_11_ );
   nand U15096 ( n15193,n15126,n11244 );
   nand U15097 ( n15201,n15202,n15203,n15129 );
   nand U15098 ( n15200,n15130,p2_datao_reg_12_ );
   nand U15099 ( n15199,n15128,p1_ir_reg_12_ );
   nand U15100 ( n15198,n15126,n11251 );
   nand U15101 ( n15207,p1_ir_reg_13_,n15208 );
   nand U15102 ( n15208,n15158,n15209 );
   nand U15103 ( n15209,n15129,n15210 );
   nand U15104 ( n15206,n15129,n15203,n15211 );
   nand U15105 ( n15205,n15130,p2_datao_reg_13_ );
   nand U15106 ( n15204,n15126,n11261 );
   nand U15107 ( n15215,n15216,n15129 );
   not U15108 ( n15216,n15217 );
   nand U15109 ( n15214,n15130,p2_datao_reg_14_ );
   nand U15110 ( n15213,n15128,p1_ir_reg_14_ );
   nand U15111 ( n15212,n15126,n11268 );
   nand U15112 ( n15221,p1_ir_reg_15_,n15222 );
   nand U15113 ( n15222,n15158,n15223 );
   nand U15114 ( n15223,n15129,n15224 );
   nand U15115 ( n15220,n15129,n15225,n15226 );
   nand U15116 ( n15219,n15130,p2_datao_reg_15_ );
   nand U15117 ( n15218,n15126,n11278 );
   nand U15118 ( n15230,n15231,n15232,n15129 );
   nand U15119 ( n15229,n15130,p2_datao_reg_16_ );
   nand U15120 ( n15228,n15128,p1_ir_reg_16_ );
   nand U15121 ( n15227,n15126,n11285 );
   nand U15122 ( n15236,p1_ir_reg_17_,n15237 );
   nand U15123 ( n15237,n15158,n15238 );
   nand U15124 ( n15238,n15129,n15239 );
   nand U15125 ( n15235,n15129,n15232,n15240 );
   nand U15126 ( n15234,n15130,p2_datao_reg_17_ );
   nand U15127 ( n15233,n15126,n11295 );
   nand U15128 ( n15244,p1_ir_reg_18_,n15245 );
   nand U15129 ( n15245,n15158,n15246 );
   nand U15130 ( n15246,n15129,n15247 );
   nand U15131 ( n15243,n15129,n15248,n15249 );
   nand U15132 ( n15242,n15130,p2_datao_reg_18_ );
   nand U15133 ( n15241,n15126,n11305 );
   nand U15134 ( n15253,n15254,n15255,n15129 );
   nand U15135 ( n15252,n15130,p2_datao_reg_19_ );
   nand U15136 ( n15251,n15128,p1_ir_reg_19_ );
   nand U15137 ( n15250,n15126,n11312 );
   nand U15138 ( n15259,n15260,n15261,n15129 );
   nand U15139 ( n15258,n15130,p2_datao_reg_20_ );
   nand U15140 ( n15257,n15128,p1_ir_reg_20_ );
   nand U15141 ( n15256,n15126,n11319 );
   nand U15142 ( n15265,p1_ir_reg_21_,n15266 );
   nand U15143 ( n15266,n15158,n15267 );
   nand U15144 ( n15267,n15129,n15268 );
   nand U15145 ( n15264,n15129,n15261,n15269 );
   nand U15146 ( n15263,n15130,p2_datao_reg_21_ );
   nand U15147 ( n15262,n15126,n11328 );
   nand U15148 ( n15273,n15274,n15275,n15129 );
   nand U15149 ( n15272,n15130,p2_datao_reg_22_ );
   nand U15150 ( n15271,n15128,p1_ir_reg_22_ );
   nand U15151 ( n15270,n15126,n11338 );
   nand U15152 ( n15279,p1_ir_reg_23_,n15280 );
   nand U15153 ( n15280,n15158,n15281 );
   nand U15154 ( n15281,n15129,n15282 );
   nand U15155 ( n15278,n15129,n15275,n15283 );
   nand U15156 ( n15277,n15130,p2_datao_reg_23_ );
   nand U15157 ( n15276,n15126,n11345 );
   nand U15158 ( n15287,n15288,n15289,n15129 );
   nand U15159 ( n15286,n15130,p2_datao_reg_24_ );
   nand U15160 ( n15285,n15128,p1_ir_reg_24_ );
   nand U15161 ( n15284,n15126,n11354 );
   nand U15162 ( n15293,p1_ir_reg_25_,n15294 );
   nand U15163 ( n15294,n15158,n15295 );
   nand U15164 ( n15295,n15129,n15296 );
   nand U15165 ( n15292,n15129,n15289,n15297 );
   nand U15166 ( n15291,n15130,p2_datao_reg_25_ );
   nand U15167 ( n15290,n15126,n11364 );
   nand U15168 ( n15301,n15302,n15303,n15129 );
   nand U15169 ( n15300,n15130,p2_datao_reg_26_ );
   nand U15170 ( n15299,n15128,p1_ir_reg_26_ );
   nand U15171 ( n15298,n15126,n11371 );
   nand U15172 ( n15307,p1_ir_reg_27_,n15308 );
   nand U15173 ( n15308,n15158,n15309 );
   nand U15174 ( n15309,n15129,n15310 );
   nand U15175 ( n15306,n15129,n15303,n15311 );
   nand U15176 ( n15305,n15130,p2_datao_reg_27_ );
   nand U15177 ( n15304,n15126,n11380 );
   nand U15178 ( n15315,n15316,n15317,n15129 );
   nand U15179 ( n15314,n15130,p2_datao_reg_28_ );
   nand U15180 ( n15313,n15128,p1_ir_reg_28_ );
   nand U15181 ( n15312,n15126,n11390 );
   nand U15182 ( n15321,p1_ir_reg_29_,n15322 );
   nand U15183 ( n15322,n15158,n15323 );
   nand U15184 ( n15323,n15324,n15129 );
   nand U15185 ( n15320,n15129,n15317,n15325 );
   not U15186 ( n15325,p1_ir_reg_29_ );
   nand U15187 ( n15319,n15130,p2_datao_reg_29_ );
   nand U15188 ( n15318,n15126,n11400 );
   nand U15189 ( n15329,p1_ir_reg_30_,n15330 );
   nand U15190 ( n15330,n15158,n15331 );
   nand U15191 ( n15331,n15332,n15129 );
   not U15192 ( n15158,n15128 );
   nand U15193 ( n15328,n15129,n15333,n15334 );
   not U15194 ( n15333,n15332 );
   nand U15195 ( n15327,n15130,p2_datao_reg_30_ );
   nand U15196 ( n15326,n15126,n11410 );
   nand U15197 ( n15337,n15126,n11415 );
   nand U15198 ( n15336,n15129,n15334,n15332 );
   nor U15199 ( n15332,n15317,p1_ir_reg_29_ );
   not U15200 ( n15334,p1_ir_reg_30_ );
   nand U15201 ( n15335,n15130,p2_datao_reg_31_ );
   nor U15202 ( n15355,n15356,n15357 );
   nor U15203 ( n15354,n15358,n15359 );
   nor U15204 ( n15359,n15082,n15088 );
   nor U15205 ( n15353,n15360,n15361 );
   nand U15206 ( n15351,n15086,p1_reg3_reg_0_ );
   nand U15207 ( n15349,n15090,n15058 );
   nand U15208 ( n15058,n15362,n15363 );
   nand U15209 ( n15363,n15364,n15365 );
   nand U15210 ( n15364,n15366,n15367 );
   nand U15211 ( n15362,n15057,n15048 );
   not U15212 ( n15057,n15360 );
   nor U15213 ( n15375,n15045,n15376 );
   nor U15214 ( n15374,n15377,n15378 );
   and U15215 ( n15373,n15044,n15090 );
   nand U15216 ( n15044,n15379,n15380 );
   nand U15217 ( n15380,n15381,n15365 );
   xor U15218 ( n15381,n15382,n15366 );
   nand U15219 ( n15379,n15122,n14590 );
   nor U15220 ( n15372,n15090,n15383 );
   nand U15221 ( n15370,n15384,n14584 );
   nand U15222 ( n15369,n15082,n15046 );
   xor U15223 ( n15046,n15056,n15385 );
   nand U15224 ( n15368,n15047,n15386 );
   xor U15225 ( n15047,n15387,n15382 );
   nor U15226 ( n15395,n15396,n15376 );
   nor U15227 ( n15394,n15397,n15378 );
   nor U15228 ( n15393,n15027,n15089 );
   and U15229 ( n15027,n15398,n15399 );
   nand U15230 ( n15399,n15400,n15401,n15402 );
   nand U15231 ( n15402,n15403,n15404,n15405 );
   nand U15232 ( n15401,n15406,n15407 );
   nand U15233 ( n15400,n15408,n15409 );
   not U15234 ( n15408,n15410 );
   nand U15235 ( n15398,n15122,n14587 );
   nor U15236 ( n15392,n15090,n15411 );
   nand U15237 ( n15390,n15384,n14581 );
   nand U15238 ( n15389,n15412,n15386 );
   not U15239 ( n15412,n15035 );
   nand U15240 ( n15035,n15413,n15414 );
   or U15241 ( n15414,n15410,n15415 );
   nand U15242 ( n15413,n15416,n15407,n15415 );
   nor U15243 ( n15415,n15417,n15418 );
   not U15244 ( n15416,n15419 );
   nand U15245 ( n15388,n15082,n15420 );
   not U15246 ( n15420,n15033 );
   nand U15247 ( n15033,n15421,n15422 );
   nand U15248 ( n15422,n15423,n15036 );
   nand U15249 ( n15423,n15045,n15358 );
   nor U15250 ( n15431,n15022,n15376 );
   nor U15251 ( n15430,p1_reg3_reg_3_,n15378 );
   and U15252 ( n15429,n15021,n15090 );
   nand U15253 ( n15021,n15432,n15433,n15434 );
   nand U15254 ( n15434,n15122,n14584 );
   nand U15255 ( n15433,n15435,n15436 );
   nand U15256 ( n15435,n15405,n15404 );
   nand U15257 ( n15432,n15437,n15436 );
   nand U15258 ( n15436,n15438,n15439 );
   or U15259 ( n15439,n15440,n15441 );
   nand U15260 ( n15438,n15440,n15441 );
   nor U15261 ( n15428,n15090,n15442 );
   nand U15262 ( n15426,n15384,n14578 );
   nand U15263 ( n15425,n15082,n15023 );
   xor U15264 ( n15023,n15421,n15443 );
   nand U15265 ( n15424,n15024,n15386 );
   xor U15266 ( n15024,n15440,n15444 );
   nand U15267 ( n15444,n15445,n15446 );
   nand U15268 ( n15446,n15417,n15447 );
   nor U15269 ( n15455,n15011,n15376 );
   nor U15270 ( n15454,n15456,n15357 );
   not U15271 ( n15357,n15384 );
   and U15272 ( n15453,n15010,n15090 );
   nand U15273 ( n15010,n15457,n15458 );
   nand U15274 ( n15458,n15459,n15460,n15365 );
   nand U15275 ( n15460,n15461,n15462,n15463 );
   or U15276 ( n15459,n15464,n15463 );
   nand U15277 ( n15457,n15122,n14581 );
   and U15278 ( n15452,n15089,p1_reg2_reg_4_ );
   nand U15279 ( n15450,n15082,n15013 );
   and U15280 ( n15013,n15465,n15466 );
   nand U15281 ( n15466,n15467,n15468 );
   nand U15282 ( n15467,n15469,n15022 );
   nand U15283 ( n15449,n15086,n15470 );
   nand U15284 ( n15448,n15012,n15386 );
   xor U15285 ( n15012,n15471,n15472 );
   nor U15286 ( n15480,n15481,n15376 );
   and U15287 ( n15479,n15482,n15086 );
   nor U15288 ( n15478,n14993,n15089 );
   and U15289 ( n14993,n15483,n15484,n15485,n15486 );
   nor U15290 ( n15486,n15487,n15488,n15489,n15490 );
   nor U15291 ( n15490,n14999,n15491 );
   nor U15292 ( n15489,n14999,n15492 );
   nor U15293 ( n15488,n15493,n15494 );
   nor U15294 ( n15487,n15495,n15494 );
   nor U15295 ( n15485,n15496,n15497 );
   nor U15296 ( n15497,n15403,n15494 );
   nor U15297 ( n15496,n14999,n15498 );
   not U15298 ( n14999,n15499 );
   or U15299 ( n15484,n15494,n15404 );
   nand U15300 ( n15494,n15500,n15501 );
   nand U15301 ( n15501,n15502,n15503,n15504 );
   nand U15302 ( n15500,n15505,n15506 );
   nand U15303 ( n15483,n15122,n14578 );
   nor U15304 ( n15477,n15090,n15507 );
   nand U15305 ( n15475,n15384,n14572 );
   nand U15306 ( n15474,n15082,n15000 );
   xor U15307 ( n15000,n15481,n15508 );
   nand U15308 ( n15473,n15087,n15499 );
   xor U15309 ( n15499,n15509,n15505 );
   nor U15310 ( n15509,n15510,n15511 );
   nor U15311 ( n15510,n15512,n15472 );
   nor U15312 ( n15520,n15521,n15376 );
   nor U15313 ( n15519,n15522,n15378 );
   nor U15314 ( n15518,n14981,n15089 );
   and U15315 ( n14981,n15523,n15524 );
   nor U15316 ( n15524,n15525,n15526,n15527,n15528 );
   nor U15317 ( n15528,n15529,n15403 );
   nor U15318 ( n15527,n15498,n14987 );
   nor U15319 ( n15526,n15529,n15404 );
   nor U15320 ( n15525,n15529,n15493 );
   nor U15321 ( n15523,n15530,n15531,n15532,n15533 );
   nor U15322 ( n15533,n15456,n15534 );
   nor U15323 ( n15532,n15491,n14987 );
   nor U15324 ( n15531,n15529,n15495 );
   nor U15325 ( n15529,n15535,n15536 );
   nor U15326 ( n15536,n15537,n15538 );
   nand U15327 ( n15538,n15539,n15540 );
   nand U15328 ( n15540,n15506,n15503 );
   not U15329 ( n15506,n15504 );
   nor U15330 ( n15535,n15541,n15542 );
   nor U15331 ( n15530,n15492,n14987 );
   nor U15332 ( n15517,n15090,n15543 );
   nand U15333 ( n15515,n15384,n14569 );
   nand U15334 ( n15514,n15082,n15544 );
   not U15335 ( n15544,n14988 );
   nand U15336 ( n14988,n15545,n15546 );
   nand U15337 ( n15546,n15547,n14990 );
   nand U15338 ( n15547,n15508,n15481 );
   or U15339 ( n15513,n15361,n14987 );
   xor U15340 ( n14987,n15539,n15548 );
   not U15341 ( n15539,n15549 );
   nor U15342 ( n15557,n15558,n15376 );
   and U15343 ( n15556,n15559,n15086 );
   nor U15344 ( n15555,n14969,n15089 );
   and U15345 ( n14969,n15560,n15561,n15562,n15563 );
   nor U15346 ( n15563,n15564,n15565,n15566,n15567 );
   nor U15347 ( n15567,n15491,n14975 );
   nor U15348 ( n15566,n15498,n14975 );
   nor U15349 ( n15565,n15492,n14975 );
   nor U15350 ( n15564,n15403,n15568 );
   nor U15351 ( n15562,n15569,n15570 );
   nor U15352 ( n15570,n15001,n15534 );
   nor U15353 ( n15569,n15495,n15568 );
   nand U15354 ( n15561,n15571,n15572 );
   nand U15355 ( n15560,n15571,n15573 );
   not U15356 ( n15571,n15568 );
   nand U15357 ( n15568,n15574,n15575 );
   nand U15358 ( n15575,n15576,n15577 );
   nand U15359 ( n15574,n15578,n15579 );
   nor U15360 ( n15554,n15090,n15580 );
   nand U15361 ( n15552,n15384,n14566 );
   nand U15362 ( n15551,n15082,n14976 );
   xor U15363 ( n14976,n15581,n15558 );
   or U15364 ( n15550,n15361,n14975 );
   nand U15365 ( n14975,n15582,n15583 );
   nand U15366 ( n15583,n15584,n15585,n15586 );
   not U15367 ( n15586,n15578 );
   nand U15368 ( n15582,n15587,n15588,n15578 );
   nand U15369 ( n15587,n15548,n15585 );
   not U15370 ( n15548,n15589 );
   nor U15371 ( n15597,n15598,n15376 );
   nor U15372 ( n15596,n15599,n15378 );
   nor U15373 ( n15595,n14957,n15089 );
   and U15374 ( n14957,n15600,n15601,n15602,n15603 );
   nor U15375 ( n15603,n15604,n15605,n15606,n15607 );
   nor U15376 ( n15607,n15608,n15404 );
   xor U15377 ( n15608,n15609,n15610 );
   nor U15378 ( n15606,n15611,n15403 );
   nor U15379 ( n15611,n15612,n15613 );
   not U15380 ( n15613,n15614 );
   nor U15381 ( n15612,n15609,n15610 );
   nor U15382 ( n15605,n15492,n14963 );
   nor U15383 ( n15604,n14989,n15534 );
   nand U15384 ( n15602,n15615,n15616 );
   nand U15385 ( n15601,n15095,n15617 );
   nand U15386 ( n15617,n15618,n15614 );
   nand U15387 ( n15614,n15609,n15610 );
   or U15388 ( n15618,n15610,n15609 );
   nor U15389 ( n15609,n15619,n15576 );
   nand U15390 ( n15600,n15615,n15620 );
   nor U15391 ( n15594,n15090,n15621 );
   nand U15392 ( n15592,n15384,n14563 );
   nand U15393 ( n15591,n15082,n15622 );
   not U15394 ( n15622,n14964 );
   nand U15395 ( n14964,n15623,n15624 );
   nand U15396 ( n15624,n15625,n14966 );
   nand U15397 ( n15625,n15581,n15558 );
   nand U15398 ( n15590,n15087,n15615 );
   not U15399 ( n15615,n14963 );
   xor U15400 ( n14963,n15610,n15626 );
   not U15401 ( n15610,n15627 );
   nor U15402 ( n15635,n14952,n15376 );
   and U15403 ( n15634,n15636,n15086 );
   and U15404 ( n15633,n14951,n15090 );
   nand U15405 ( n14951,n15637,n15638 );
   nand U15406 ( n15638,n15639,n15640,n15365 );
   nand U15407 ( n15640,n15641,n15642 );
   nand U15408 ( n15639,n15643,n15644,n15645 );
   nand U15409 ( n15637,n15122,n14566 );
   and U15410 ( n15632,n15089,p1_reg2_reg_9_ );
   nand U15411 ( n15630,n15384,n14560 );
   nand U15412 ( n15629,n15082,n14953 );
   xor U15413 ( n14953,n15646,n15623 );
   nand U15414 ( n15628,n14954,n15386 );
   xor U15415 ( n14954,n15641,n15647 );
   nor U15416 ( n15655,n14941,n15376 );
   nor U15417 ( n15654,n15656,n15378 );
   and U15418 ( n15653,n14940,n15090 );
   nand U15419 ( n14940,n15657,n15658,n15659,n15660 );
   nor U15420 ( n15660,n15661,n15662,n15663,n15664 );
   nor U15421 ( n15664,n15495,n15665 );
   nor U15422 ( n15663,n15491,n15666 );
   nor U15423 ( n15662,n15498,n15666 );
   nor U15424 ( n15661,n15492,n15666 );
   or U15425 ( n15659,n15665,n15493 );
   or U15426 ( n15658,n15665,n15109 );
   nand U15427 ( n15665,n15667,n15668 );
   nand U15428 ( n15668,n15669,n15670,n15671 );
   nand U15429 ( n15667,n15672,n15673 );
   nand U15430 ( n15657,n15122,n14563 );
   nor U15431 ( n15652,n15090,n15674 );
   nand U15432 ( n15650,n15384,n14557 );
   nand U15433 ( n15649,n15082,n14942 );
   and U15434 ( n14942,n15675,n15676 );
   nand U15435 ( n15676,n15677,n15678 );
   nand U15436 ( n15677,n15679,n14952 );
   nand U15437 ( n15648,n15087,n14943 );
   not U15438 ( n14943,n15666 );
   nand U15439 ( n15666,n15680,n15681 );
   nand U15440 ( n15681,n15682,n15683,n15684 );
   not U15441 ( n15684,n15672 );
   nand U15442 ( n15682,n15685,n15647 );
   not U15443 ( n15647,n15686 );
   nand U15444 ( n15680,n15687,n15685,n15672 );
   nand U15445 ( n15687,n15686,n15683 );
   nor U15446 ( n15686,n15688,n15689 );
   nor U15447 ( n15697,n15698,n15376 );
   nor U15448 ( n15696,n15699,n15378 );
   nor U15449 ( n15695,n14923,n15089 );
   and U15450 ( n14923,n15700,n15701 );
   nor U15451 ( n15701,n15702,n15703,n15704,n15705 );
   nor U15452 ( n15705,n15706,n15403 );
   nor U15453 ( n15704,n15492,n14929 );
   nor U15454 ( n15703,n15707,n15534 );
   nor U15455 ( n15702,n15706,n15493 );
   nor U15456 ( n15700,n15708,n15709,n15710,n15711 );
   nor U15457 ( n15711,n15706,n15495 );
   and U15458 ( n15706,n15712,n15713,n15714 );
   not U15459 ( n15714,n15715 );
   nand U15460 ( n15713,n15716,n15671 );
   nand U15461 ( n15712,n15673,n15717 );
   not U15462 ( n15673,n15671 );
   nor U15463 ( n15710,n15491,n14929 );
   nor U15464 ( n15709,n15498,n14929 );
   nor U15465 ( n15708,n15718,n15404 );
   nor U15466 ( n15718,n15715,n15719,n15720 );
   nor U15467 ( n15720,n15721,n15671 );
   and U15468 ( n15719,n15671,n15716 );
   nand U15469 ( n15671,n15644,n15722 );
   nand U15470 ( n15722,n15645,n15643 );
   nand U15471 ( n15715,n15723,n15724 );
   nand U15472 ( n15724,n15725,n15716 );
   nor U15473 ( n15716,n15726,n15727 );
   nand U15474 ( n15723,n15727,n15717 );
   not U15475 ( n15717,n15721 );
   nand U15476 ( n15721,n15728,n15729 );
   nor U15477 ( n15694,n15090,n15730 );
   nand U15478 ( n15692,n15384,n14554 );
   nand U15479 ( n15691,n15082,n14930 );
   xor U15480 ( n14930,n15731,n15698 );
   or U15481 ( n15690,n15361,n14929 );
   xor U15482 ( n14929,n15732,n15726 );
   not U15483 ( n15726,n15733 );
   nor U15484 ( n15741,n14918,n15376 );
   nor U15485 ( n15740,n15742,n15378 );
   and U15486 ( n15739,n14917,n15090 );
   nand U15487 ( n14917,n15743,n15744 );
   nand U15488 ( n15744,n15745,n15365 );
   nand U15489 ( n15365,n15405,n15109 );
   not U15490 ( n15405,n15095 );
   xor U15491 ( n15745,n15746,n15747 );
   nand U15492 ( n15743,n15122,n14557 );
   nor U15493 ( n15738,n15090,n15748 );
   nand U15494 ( n15736,n15384,n14551 );
   nand U15495 ( n15735,n14919,n15386 );
   xor U15496 ( n14919,n15749,n15747 );
   nand U15497 ( n15734,n15082,n14920 );
   and U15498 ( n14920,n15750,n15751 );
   nand U15499 ( n15751,n15752,n15753 );
   nand U15500 ( n15752,n15731,n15698 );
   nor U15501 ( n15761,n15762,n15376 );
   nor U15502 ( n15760,n15763,n15378 );
   nor U15503 ( n15759,n14900,n15089 );
   and U15504 ( n14900,n15764,n15765,n15766,n15767 );
   nor U15505 ( n15767,n15768,n15769,n15770,n15771 );
   nor U15506 ( n15771,n15403,n15772 );
   nor U15507 ( n15770,n15493,n15772 );
   nor U15508 ( n15769,n14931,n15534 );
   nor U15509 ( n15768,n15495,n15772 );
   nor U15510 ( n15766,n15773,n15774 );
   nor U15511 ( n15774,n15492,n14906 );
   nor U15512 ( n15773,n15404,n15772 );
   xor U15513 ( n15772,n15775,n15776 );
   nand U15514 ( n15765,n15777,n15620 );
   nand U15515 ( n15764,n15777,n15616 );
   nor U15516 ( n15758,n15090,n15778 );
   nand U15517 ( n15756,n15384,n14548 );
   nand U15518 ( n15755,n15082,n14907 );
   xor U15519 ( n14907,n15762,n15779 );
   nand U15520 ( n15754,n15087,n15777 );
   not U15521 ( n15777,n14906 );
   nand U15522 ( n14906,n15780,n15781 );
   nand U15523 ( n15781,n15782,n15783,n15775 );
   nand U15524 ( n15782,n15784,n15749 );
   not U15525 ( n15749,n15785 );
   nand U15526 ( n15780,n15786,n15784,n15787 );
   nand U15527 ( n15786,n15785,n15783 );
   nor U15528 ( n15785,n15788,n15789 );
   nor U15529 ( n15797,n14895,n15376 );
   and U15530 ( n15796,n15798,n15086 );
   and U15531 ( n15795,n14894,n15090 );
   nand U15532 ( n14894,n15799,n15800 );
   nand U15533 ( n15800,n15801,n15802,n15803 );
   nand U15534 ( n15802,n15804,n15805 );
   nand U15535 ( n15801,n15806,n15807,n15808 );
   nand U15536 ( n15799,n15122,n14551 );
   nor U15537 ( n15794,n15090,n15809 );
   nand U15538 ( n15792,n15384,n14545 );
   nand U15539 ( n15791,n14896,n15386 );
   xor U15540 ( n14896,n15804,n15810 );
   nand U15541 ( n15790,n15082,n14897 );
   and U15542 ( n14897,n15811,n15812 );
   nand U15543 ( n15812,n15813,n15814 );
   nand U15544 ( n15813,n15779,n15762 );
   nor U15545 ( n15822,n14884,n15376 );
   nor U15546 ( n15821,n15823,n15378 );
   and U15547 ( n15820,n14883,n15090 );
   nand U15548 ( n14883,n15824,n15825 );
   nand U15549 ( n15825,n15826,n15827,n15803 );
   nand U15550 ( n15803,n15828,n15493 );
   and U15551 ( n15828,n15109,n15495 );
   nand U15552 ( n15827,n15829,n15830,n15831 );
   nand U15553 ( n15826,n15832,n15833 );
   nand U15554 ( n15824,n15122,n14548 );
   nor U15555 ( n15819,n15090,n15834 );
   nand U15556 ( n15817,n15384,n14542 );
   nand U15557 ( n15816,n15082,n14885 );
   xor U15558 ( n14885,n15811,n15835 );
   nand U15559 ( n15815,n14886,n15386 );
   xor U15560 ( n14886,n15836,n15837 );
   not U15561 ( n15836,n15832 );
   nor U15562 ( n15845,n15846,n15376 );
   nor U15563 ( n15844,n15847,n15378 );
   nor U15564 ( n15843,n14867,n15089 );
   and U15565 ( n14867,n15848,n15849 );
   nor U15566 ( n15849,n15850,n15851,n15852,n15853 );
   nor U15567 ( n15853,n15403,n15854,n15855 );
   nor U15568 ( n15855,n15856,n15857 );
   and U15569 ( n15857,n15858,n15859 );
   nor U15570 ( n15856,n15860,n15861,n15862 );
   nor U15571 ( n15862,n15863,n15831 );
   nor U15572 ( n15854,n15833,n15861,n15864 );
   nor U15573 ( n15852,n15865,n15404 );
   nor U15574 ( n15851,n14873,n15491 );
   nor U15575 ( n15850,n15865,n15493 );
   nor U15576 ( n15848,n15866,n15867,n15868,n15869 );
   nor U15577 ( n15869,n14873,n15498 );
   nor U15578 ( n15868,n14873,n15492 );
   nor U15579 ( n15867,n15865,n15495 );
   and U15580 ( n15865,n15870,n15871,n15872,n15873 );
   nand U15581 ( n15873,n15864,n15829,n15831 );
   nand U15582 ( n15872,n15859,n15858,n15833 );
   not U15583 ( n15833,n15831 );
   nand U15584 ( n15871,n15859,n15858,n15861 );
   nand U15585 ( n15870,n15863,n15864 );
   nor U15586 ( n15866,n15874,n15534 );
   nor U15587 ( n15842,n15090,n15875 );
   nand U15588 ( n15840,n15384,n14539 );
   nand U15589 ( n15839,n15082,n15876 );
   not U15590 ( n15876,n14874 );
   nand U15591 ( n14874,n15877,n15878 );
   nand U15592 ( n15878,n15879,n14875 );
   nand U15593 ( n15879,n15880,n14884 );
   or U15594 ( n15838,n15361,n14873 );
   xor U15595 ( n14873,n15881,n15864 );
   not U15596 ( n15864,n15860 );
   nor U15597 ( n15889,n15890,n15376 );
   nor U15598 ( n15888,n15891,n15378 );
   nor U15599 ( n15887,n14855,n15089 );
   and U15600 ( n14855,n15892,n15893,n15894,n15895 );
   nor U15601 ( n15895,n15896,n15897,n15898,n15899 );
   nor U15602 ( n15899,n15403,n15900 );
   nor U15603 ( n15898,n15493,n15900 );
   nor U15604 ( n15897,n15901,n15534 );
   nor U15605 ( n15896,n15495,n15900 );
   nor U15606 ( n15894,n15902,n15903 );
   nor U15607 ( n15903,n15492,n14861 );
   nor U15608 ( n15902,n15404,n15900 );
   xor U15609 ( n15900,n15904,n15905 );
   nand U15610 ( n15893,n15906,n15620 );
   nand U15611 ( n15892,n15906,n15616 );
   nor U15612 ( n15886,n15090,n15907 );
   nand U15613 ( n15884,n15384,n14536 );
   nand U15614 ( n15883,n15082,n14862 );
   xor U15615 ( n14862,n15890,n15908 );
   nand U15616 ( n15882,n15087,n15906 );
   not U15617 ( n15906,n14861 );
   nand U15618 ( n14861,n15909,n15910 );
   nand U15619 ( n15910,n15911,n15912,n15904 );
   nand U15620 ( n15909,n15913,n15914,n15915 );
   nand U15621 ( n15913,n15912,n15881 );
   nor U15622 ( n15919,n15920,n15921,n15922,n15923 );
   nor U15623 ( n15923,n14850,n15376 );
   nor U15624 ( n15922,n15924,n15378 );
   and U15625 ( n15921,n14849,n15090 );
   nand U15626 ( n14849,n15925,n15926 );
   nand U15627 ( n15926,n15927,n15928 );
   xor U15628 ( n15927,n15929,n15930 );
   nand U15629 ( n15925,n15122,n14539 );
   nor U15630 ( n15920,n15090,n15931 );
   nand U15631 ( n15918,n15384,n14533 );
   nand U15632 ( n15917,n14851,n15386 );
   xor U15633 ( n14851,n15929,n15932 );
   nand U15634 ( n15916,n15082,n14852 );
   and U15635 ( n14852,n15933,n15934 );
   nand U15636 ( n15934,n15935,n15936 );
   nand U15637 ( n15935,n15908,n15890 );
   nor U15638 ( n15940,n15941,n15942,n15943,n15944 );
   nor U15639 ( n15944,n14839,n15376 );
   nor U15640 ( n15943,n15945,n15378 );
   and U15641 ( n15942,n14838,n15090 );
   nand U15642 ( n14838,n15946,n15947,n15948 );
   nand U15643 ( n15948,n15122,n14536 );
   nand U15644 ( n15947,n14841,n15048 );
   nand U15645 ( n15946,n15949,n15928 );
   nand U15646 ( n15928,n15495,n15403,n15493,n15404 );
   xor U15647 ( n15949,n15950,n15951 );
   nor U15648 ( n15941,n15090,n15952 );
   nand U15649 ( n15939,n15384,n14530 );
   nand U15650 ( n15938,n15082,n14840 );
   xor U15651 ( n14840,n15933,n15953 );
   nand U15652 ( n15937,n15087,n14841 );
   xor U15653 ( n14841,n15950,n15954 );
   nor U15654 ( n15958,n15959,n15960,n15961,n15962 );
   nor U15655 ( n15962,n14828,n15376 );
   nor U15656 ( n15961,n15963,n15378 );
   and U15657 ( n15960,n14827,n15090 );
   nand U15658 ( n14827,n15964,n15965 );
   nor U15659 ( n15965,n15966,n15967,n15968,n15969 );
   nor U15660 ( n15969,n15491,n15970 );
   nor U15661 ( n15968,n15498,n15970 );
   nor U15662 ( n15967,n15492,n15970 );
   nor U15663 ( n15966,n15404,n15971 );
   nor U15664 ( n15964,n15972,n15973,n15974,n15975 );
   nor U15665 ( n15975,n15403,n15971 );
   nor U15666 ( n15974,n15493,n15971 );
   nor U15667 ( n15973,n15976,n15534 );
   nor U15668 ( n15972,n15495,n15971 );
   xor U15669 ( n15971,n15977,n15978 );
   and U15670 ( n15959,n15089,p1_reg2_reg_20_ );
   nand U15671 ( n15957,n15384,n14527 );
   nand U15672 ( n15956,n15082,n14829 );
   and U15673 ( n14829,n15979,n15980 );
   nand U15674 ( n15980,n15981,n15982 );
   nand U15675 ( n15981,n15983,n14839 );
   nand U15676 ( n15955,n15087,n14830 );
   not U15677 ( n14830,n15970 );
   nand U15678 ( n15970,n15984,n15985 );
   nand U15679 ( n15985,n15986,n15987,n15988 );
   nand U15680 ( n15986,n15989,n15990 );
   nand U15681 ( n15984,n15977,n15990,n15991 );
   nand U15682 ( n15991,n15954,n15992 );
   nor U15683 ( n15996,n15997,n15998,n15999,n16000 );
   nor U15684 ( n16000,n16001,n15376 );
   and U15685 ( n15999,n16002,n15086 );
   nor U15686 ( n15998,n14810,n15089 );
   and U15687 ( n14810,n16003,n16004,n16005,n16006 );
   nor U15688 ( n16006,n16007,n16008,n16009,n16010 );
   nor U15689 ( n16010,n15495,n16011 );
   nor U15690 ( n16009,n15403,n16011 );
   nor U15691 ( n16008,n16012,n15534 );
   nor U15692 ( n16007,n15493,n16011 );
   nor U15693 ( n16005,n16013,n16014 );
   nor U15694 ( n16014,n16015,n16016,n16017,n15491 );
   nor U15695 ( n16016,n16018,n16019,n16020 );
   nor U15696 ( n16020,n15989,n16021 );
   nor U15697 ( n16015,n16022,n16023 );
   nor U15698 ( n16013,n15492,n14816 );
   or U15699 ( n16004,n16011,n15404 );
   nand U15700 ( n16011,n16024,n16025 );
   nand U15701 ( n16025,n16019,n16026 );
   nand U15702 ( n16024,n16027,n16028,n16029 );
   nand U15703 ( n16003,n16030,n15620 );
   and U15704 ( n15997,n15089,p1_reg2_reg_21_ );
   nand U15705 ( n15995,n15384,n14524 );
   nand U15706 ( n15994,n15082,n14817 );
   xor U15707 ( n14817,n16001,n16031 );
   nand U15708 ( n15993,n15087,n16030 );
   not U15709 ( n16030,n14816 );
   nand U15710 ( n14816,n16032,n16033,n16034 );
   not U15711 ( n16034,n16017 );
   nor U15712 ( n16017,n16021,n15989,n16023 );
   nand U15713 ( n16033,n16019,n16018 );
   not U15714 ( n16019,n16023 );
   nand U15715 ( n16032,n16035,n16023,n16022 );
   nand U15716 ( n16035,n15988,n15954 );
   not U15717 ( n15954,n15989 );
   nor U15718 ( n15989,n16036,n16037 );
   nor U15719 ( n16041,n16042,n16043,n16044,n16045 );
   nor U15720 ( n16045,n14804,n15376 );
   nor U15721 ( n16044,n16046,n15378 );
   and U15722 ( n16043,n14802,n15090 );
   nand U15723 ( n14802,n16047,n16048 );
   nand U15724 ( n16048,n16049,n16050,n16051 );
   nand U15725 ( n16051,n15495,n15493,n15109 );
   nand U15726 ( n16050,n16052,n16053,n16054 );
   nand U15727 ( n16049,n16055,n16056 );
   nand U15728 ( n16047,n15122,n14527 );
   and U15729 ( n16042,n15089,p1_reg2_reg_22_ );
   nand U15730 ( n16040,n15384,n14521 );
   nand U15731 ( n16039,n14805,n15386 );
   nand U15732 ( n15386,n15361,n16057 );
   nand U15733 ( n16057,n15090,n15048 );
   nand U15734 ( n15048,n16058,n15491 );
   nor U15735 ( n16058,n16059,n15620 );
   xor U15736 ( n14805,n16055,n16060 );
   nand U15737 ( n16038,n15082,n14807 );
   and U15738 ( n14807,n16061,n16062 );
   nand U15739 ( n16062,n16063,n16064 );
   nand U15740 ( n16063,n16031,n16001 );
   nor U15741 ( n16072,n16073,n15376 );
   and U15742 ( n16071,n16074,n15086 );
   nor U15743 ( n16070,n14785,n15089 );
   and U15744 ( n14785,n16075,n16076,n16077,n16078 );
   nor U15745 ( n16078,n16079,n16080,n16081,n16082 );
   nor U15746 ( n16082,n15403,n16083,n16084 );
   nor U15747 ( n16084,n16085,n16086 );
   nor U15748 ( n16086,n16087,n16088 );
   not U15749 ( n16088,n16089 );
   nor U15750 ( n16087,n16090,n16054 );
   nor U15751 ( n16083,n16089,n16091,n16056 );
   nor U15752 ( n16081,n14791,n15498 );
   nor U15753 ( n16080,n16092,n15404 );
   nor U15754 ( n16079,n14791,n15491 );
   not U15755 ( n14791,n16093 );
   nor U15756 ( n16077,n16094,n16095 );
   nor U15757 ( n16095,n16092,n15495 );
   not U15758 ( n16092,n16096 );
   nor U15759 ( n16094,n14818,n15534 );
   nand U15760 ( n16076,n15572,n16096 );
   nand U15761 ( n16096,n16097,n16098 );
   nand U15762 ( n16098,n16089,n16099 );
   nand U15763 ( n16099,n16056,n16053 );
   nor U15764 ( n16089,n16100,n16091 );
   nand U15765 ( n16097,n16085,n16101 );
   nand U15766 ( n16101,n16052,n16054 );
   not U15767 ( n16054,n16056 );
   nor U15768 ( n16056,n16102,n16103 );
   and U15769 ( n16085,n16104,n16105 );
   nand U15770 ( n16075,n16059,n16093 );
   and U15771 ( n16069,n15089,p1_reg2_reg_23_ );
   nand U15772 ( n16067,n15384,n14518 );
   nand U15773 ( n16066,n15082,n14792 );
   xor U15774 ( n14792,n16106,n16073 );
   nand U15775 ( n16065,n15087,n16093 );
   xor U15776 ( n16093,n16107,n16100 );
   nor U15777 ( n16111,n16112,n16113,n16114,n16115 );
   nor U15778 ( n16115,n16116,n15376 );
   and U15779 ( n16114,n16117,n15086 );
   nor U15780 ( n16113,n14774,n15089 );
   and U15781 ( n14774,n16118,n16119,n16120,n16121 );
   nor U15782 ( n16121,n16122,n16123,n16124,n16125 );
   nor U15783 ( n16125,n16126,n15534 );
   nor U15784 ( n16124,n16127,n15495 );
   nor U15785 ( n16123,n14780,n15498 );
   nor U15786 ( n16122,n16127,n15404 );
   nor U15787 ( n16120,n16128,n16129 );
   nor U15788 ( n16129,n16127,n15493 );
   nor U15789 ( n16128,n14780,n15492 );
   not U15790 ( n14780,n16130 );
   or U15791 ( n16119,n15403,n16127 );
   xor U15792 ( n16127,n16131,n16132 );
   nand U15793 ( n16118,n15616,n16130 );
   and U15794 ( n16112,n15089,p1_reg2_reg_24_ );
   nand U15795 ( n16110,n15384,n14515 );
   nand U15796 ( n16109,n15082,n16133 );
   not U15797 ( n16133,n14781 );
   nand U15798 ( n14781,n16134,n16135 );
   nand U15799 ( n16135,n16136,n14782 );
   nand U15800 ( n16136,n16106,n16073 );
   nand U15801 ( n16108,n15087,n16130 );
   xor U15802 ( n16130,n16137,n16131 );
   nor U15803 ( n16141,n16142,n16143,n16144,n16145 );
   nor U15804 ( n16145,n16146,n15376 );
   and U15805 ( n16144,n16147,n15086 );
   nor U15806 ( n16143,n14762,n15089 );
   and U15807 ( n14762,n16148,n16149,n16150,n16151 );
   nor U15808 ( n16151,n16152,n16153,n16154,n16155 );
   nor U15809 ( n16155,n15404,n16156 );
   nor U15810 ( n16154,n14769,n15491 );
   nor U15811 ( n16153,n15493,n16156 );
   nor U15812 ( n16152,n15495,n16156 );
   nor U15813 ( n16150,n16157,n16158 );
   nor U15814 ( n16158,n15403,n16156 );
   xor U15815 ( n16156,n16159,n16160 );
   nor U15816 ( n16157,n14769,n15492 );
   not U15817 ( n14769,n16161 );
   nand U15818 ( n16149,n15122,n14518 );
   nand U15819 ( n16148,n15620,n16161 );
   and U15820 ( n16142,n15089,p1_reg2_reg_25_ );
   nand U15821 ( n16140,n15384,n14512 );
   nand U15822 ( n16139,n15082,n14770 );
   xor U15823 ( n14770,n16162,n16146 );
   nand U15824 ( n16138,n15087,n16161 );
   xor U15825 ( n16161,n16159,n16163 );
   nor U15826 ( n16167,n16168,n16169,n16170,n16171 );
   nor U15827 ( n16171,n16172,n15376 );
   nor U15828 ( n16170,n16173,n15378 );
   nor U15829 ( n16169,n14749,n15089 );
   and U15830 ( n14749,n16174,n16175,n16176,n16177 );
   nor U15831 ( n16177,n16178,n16179,n16180,n16181 );
   nor U15832 ( n16181,n15491,n14755 );
   nor U15833 ( n16180,n15498,n14755 );
   nor U15834 ( n16179,n15492,n14755 );
   and U15835 ( n16178,n15437,n16182,n16183 );
   nor U15836 ( n16176,n16184,n16185 );
   nor U15837 ( n16185,n15493,n16186 );
   nor U15838 ( n16184,n15495,n16186 );
   nand U15839 ( n16186,n16187,n16183 );
   nand U15840 ( n16187,n16188,n16189 );
   nand U15841 ( n16175,n15122,n14515 );
   nand U15842 ( n16174,n16183,n16182,n15573 );
   nand U15843 ( n16182,n16190,n16189 );
   nand U15844 ( n16183,n16191,n16192 );
   and U15845 ( n16168,n15089,p1_reg2_reg_26_ );
   nand U15846 ( n16166,n15384,n14509 );
   nand U15847 ( n16165,n15082,n16193 );
   not U15848 ( n16193,n14757 );
   nand U15849 ( n14757,n16194,n16195 );
   nand U15850 ( n16195,n16196,n14759 );
   nand U15851 ( n16196,n16162,n16146 );
   or U15852 ( n16164,n15361,n14755 );
   nand U15853 ( n14755,n16197,n16198 );
   nand U15854 ( n16198,n16199,n16200,n16201 );
   nand U15855 ( n16199,n16202,n16203 );
   not U15856 ( n16202,n16163 );
   nand U15857 ( n16197,n16204,n16203,n16191 );
   nand U15858 ( n16204,n16200,n16163 );
   nand U15859 ( n16163,n16205,n16206 );
   nand U15860 ( n16206,n16207,n16137 );
   nor U15861 ( n16211,n16212,n16213,n16214,n16215 );
   nor U15862 ( n16215,n16216,n15376 );
   and U15863 ( n16214,n16217,n15086 );
   nor U15864 ( n16213,n14737,n15089 );
   and U15865 ( n14737,n16218,n16219,n16220,n16221 );
   nor U15866 ( n16221,n16222,n16223,n16224,n16225 );
   nor U15867 ( n16225,n15492,n14743 );
   nor U15868 ( n16224,n16226,n15493 );
   nor U15869 ( n16223,n16226,n15495 );
   nor U15870 ( n16226,n16227,n16228 );
   and U15871 ( n16228,n16229,n16230 );
   nand U15872 ( n16230,n16231,n16232 );
   nand U15873 ( n16229,n16188,n16233 );
   nor U15874 ( n16222,n16234,n15534 );
   nor U15875 ( n16220,n16235,n16236 );
   nor U15876 ( n16236,n16237,n15404 );
   nor U15877 ( n16237,n16227,n16238,n16239 );
   and U15878 ( n16239,n16190,n16240 );
   nor U15879 ( n16238,n16190,n16231 );
   nor U15880 ( n16227,n16233,n16189 );
   nor U15881 ( n16235,n15491,n14743 );
   nand U15882 ( n16219,n16241,n15620 );
   nand U15883 ( n16218,n16242,n16243,n15437 );
   nand U15884 ( n16243,n16190,n16233 );
   nand U15885 ( n16242,n16244,n16231 );
   nand U15886 ( n16231,n16233,n16189 );
   nand U15887 ( n16244,n16245,n16246,n16240 );
   nand U15888 ( n16245,n16192,n16189 );
   and U15889 ( n16212,n15089,p1_reg2_reg_27_ );
   nand U15890 ( n16210,n15384,n14506 );
   nand U15891 ( n16209,n15082,n14744 );
   xor U15892 ( n14744,n16247,n16216 );
   nand U15893 ( n16208,n15087,n16241 );
   not U15894 ( n16241,n14743 );
   xor U15895 ( n14743,n16233,n16248 );
   nand U15896 ( n16248,n16249,n16250,n16251 );
   nand U15897 ( n16249,n16252,n16203,n16253 );
   nor U15898 ( n16257,n16258,n16259,n16260,n16261 );
   nor U15899 ( n16261,n16262,n15376 );
   and U15900 ( n16260,n16263,n15086 );
   nor U15901 ( n15086,n15089,n16264 );
   nor U15902 ( n16259,n14723,n15089 );
   and U15903 ( n14723,n16265,n16266,n16267,n16268 );
   nor U15904 ( n16268,n16269,n16270,n16271,n16272 );
   nor U15905 ( n16272,n14730,n15491 );
   nor U15906 ( n16271,n14730,n15498 );
   nor U15907 ( n16270,n16273,n15495 );
   nor U15908 ( n16269,n14758,n15534 );
   not U15909 ( n15534,n15122 );
   nor U15910 ( n15122,n16274,n16275 );
   nor U15911 ( n16267,n16276,n16277 );
   nor U15912 ( n16277,n16273,n15493 );
   xor U15913 ( n16273,n15101,n16278 );
   nand U15914 ( n15101,n16279,n16280 );
   nand U15915 ( n16280,n16188,n16281 );
   not U15916 ( n16188,n16232 );
   nand U15917 ( n16232,n16282,n16246,n16283 );
   nor U15918 ( n16276,n14730,n15492 );
   nand U15919 ( n16266,n15437,n16284 );
   nand U15920 ( n16265,n15573,n16284 );
   xor U15921 ( n16284,n15113,n16285 );
   nand U15922 ( n15113,n16279,n16286 );
   nand U15923 ( n16286,n16190,n16281 );
   nor U15924 ( n16190,n16192,n16287 );
   not U15925 ( n16287,n16246 );
   nand U15926 ( n16192,n16282,n16283 );
   nand U15927 ( n16283,n16160,n16288 );
   nand U15928 ( n16160,n16289,n16290 );
   nand U15929 ( n16290,n16132,n16291 );
   and U15930 ( n16132,n16292,n16293 );
   nand U15931 ( n16293,n16105,n16294 );
   nand U15932 ( n16294,n16104,n16295 );
   nand U15933 ( n16295,n16103,n16052 );
   and U15934 ( n16104,n16053,n16296 );
   nand U15935 ( n16296,n16073,n14521 );
   nand U15936 ( n16292,n16105,n16052,n16102 );
   and U15937 ( n16102,n16029,n16027 );
   not U15938 ( n16029,n16026 );
   nand U15939 ( n16026,n16297,n16298 );
   nand U15940 ( n16298,n16012,n16299 );
   or U15941 ( n16299,n15978,n15982 );
   nand U15942 ( n16297,n15978,n15982 );
   nand U15943 ( n15978,n16300,n16301 );
   nand U15944 ( n16301,n15951,n16302 );
   nand U15945 ( n15951,n16303,n16304 );
   nand U15946 ( n16304,n16305,n15930 );
   nand U15947 ( n15930,n16306,n16307 );
   nand U15948 ( n16307,n16308,n15905 );
   nand U15949 ( n15905,n16309,n15858 );
   nand U15950 ( n16309,n15859,n16310 );
   nand U15951 ( n16310,n15831,n15829 );
   nand U15952 ( n15831,n16311,n15807 );
   nand U15953 ( n16311,n15808,n15806 );
   not U15954 ( n15808,n15805 );
   nand U15955 ( n15805,n16312,n16313 );
   nand U15956 ( n16313,n16314,n15776 );
   nand U15957 ( n15776,n16315,n16316 );
   nand U15958 ( n16316,n15746,n16317 );
   nand U15959 ( n16317,n14918,n14554 );
   and U15960 ( n15746,n16318,n16319 );
   nand U15961 ( n16319,n15729,n16320 );
   nand U15962 ( n16320,n15728,n16321 );
   or U15963 ( n16321,n15644,n15727 );
   and U15964 ( n15728,n15670,n16322 );
   nand U15965 ( n16322,n15698,n14557 );
   nand U15966 ( n16318,n15645,n16323 );
   not U15967 ( n15645,n15642 );
   nand U15968 ( n15642,n16324,n16325 );
   nand U15969 ( n16324,n16326,n16327 );
   not U15970 ( n16327,n15576 );
   nor U15971 ( n15576,n15579,n16328 );
   nand U15972 ( n15579,n15541,n16329 );
   nand U15973 ( n15541,n16330,n15503,n16331 );
   nand U15974 ( n16331,n15502,n15504 );
   nand U15975 ( n15504,n16332,n15462 );
   nand U15976 ( n16332,n15463,n15461 );
   nand U15977 ( n15463,n16333,n16334 );
   nand U15978 ( n16334,n16335,n14581 );
   or U15979 ( n16335,n15441,n15022 );
   nand U15980 ( n16333,n15022,n15441 );
   nand U15981 ( n15441,n16336,n15407 );
   not U15982 ( n16336,n15406 );
   nor U15983 ( n15406,n15409,n15419 );
   not U15984 ( n16308,n16337 );
   and U15985 ( n16279,n16338,n16339 );
   or U15986 ( n16339,n16189,n16340 );
   and U15987 ( n16258,n15089,p1_reg2_reg_28_ );
   or U15988 ( n16256,n15361,n14730 );
   xor U15989 ( n14730,n16285,n15121 );
   nand U15990 ( n15121,n16341,n16342,n16343,n16344 );
   nand U15991 ( n16343,n16253,n16345,n16252,n16203 );
   nand U15992 ( n16253,n16200,n16207 );
   nand U15993 ( n16342,n16346,n16345 );
   not U15994 ( n16346,n16250 );
   nand U15995 ( n16250,n16347,n16205,n16252,n16203 );
   not U15996 ( n16347,n16137 );
   nand U15997 ( n16137,n16348,n16349 );
   nand U15998 ( n16349,n16126,n16350 );
   or U15999 ( n16350,n16107,n16073 );
   nand U16000 ( n16348,n16073,n16107 );
   nand U16001 ( n16107,n16351,n16352 );
   nand U16002 ( n16352,n14818,n16353 );
   nand U16003 ( n16353,n16064,n16060 );
   or U16004 ( n16351,n16060,n16064 );
   nand U16005 ( n16060,n16354,n16355,n16356 );
   nand U16006 ( n16356,n16357,n16358 );
   nand U16007 ( n16358,n16022,n16359 );
   nand U16008 ( n16359,n16036,n15988 );
   not U16009 ( n16022,n16018 );
   nand U16010 ( n16018,n15987,n16360 );
   nand U16011 ( n16360,n16361,n16362 );
   nand U16012 ( n16354,n15988,n16357,n16037 );
   and U16013 ( n16037,n16363,n15932 );
   nand U16014 ( n15932,n16364,n16365 );
   nand U16015 ( n16365,n16366,n16367 );
   nand U16016 ( n16366,n15912,n15911 );
   nand U16017 ( n15911,n16368,n15914 );
   not U16018 ( n16368,n15881 );
   nand U16019 ( n15881,n16369,n16370 );
   nand U16020 ( n16370,n15874,n16371 );
   or U16021 ( n16371,n15837,n14884 );
   nand U16022 ( n16369,n14884,n15837 );
   nand U16023 ( n15837,n16372,n16373 );
   nand U16024 ( n16373,n14908,n16374 );
   nand U16025 ( n16374,n15814,n15810 );
   or U16026 ( n16372,n15810,n15814 );
   nand U16027 ( n15810,n16375,n16376 );
   nand U16028 ( n16376,n16377,n15784,n15788 );
   and U16029 ( n15788,n15732,n16378 );
   nand U16030 ( n16378,n16379,n15698 );
   nand U16031 ( n15732,n16380,n16381,n16382 );
   nand U16032 ( n16382,n16383,n15678 );
   nand U16033 ( n16381,n16384,n15685,n15688 );
   and U16034 ( n15688,n15626,n16385 );
   nand U16035 ( n16385,n14977,n15598 );
   nand U16036 ( n15626,n16386,n16387 );
   nand U16037 ( n16387,n16388,n16389 );
   nand U16038 ( n16389,n14989,n15558 );
   nand U16039 ( n16388,n15585,n15584 );
   nand U16040 ( n15584,n15589,n15588 );
   nand U16041 ( n15589,n16390,n16391,n16392 );
   nand U16042 ( n16392,n15512,n15002 );
   nand U16043 ( n16391,n15472,n16393,n16394 );
   nand U16044 ( n16394,n15456,n15481 );
   not U16045 ( n16393,n15511 );
   nand U16046 ( n15472,n16395,n16396,n16397 );
   nand U16047 ( n16397,n16398,n15443 );
   nand U16048 ( n16396,n16399,n15447,n15417 );
   nor U16049 ( n15417,n15387,n16400 );
   nor U16050 ( n16400,n14587,n15385 );
   nand U16051 ( n16399,n16401,n15022 );
   nand U16052 ( n16395,n16402,n14581 );
   nand U16053 ( n16402,n15445,n15022 );
   not U16054 ( n15445,n16398 );
   nand U16055 ( n16398,n16403,n16404 );
   nand U16056 ( n16404,n15418,n15447 );
   nand U16057 ( n16390,n16405,n14575 );
   or U16058 ( n16405,n15002,n15512 );
   nand U16059 ( n16386,n14978,n14569 );
   nand U16060 ( n16384,n15707,n14941 );
   nand U16061 ( n16380,n16406,n14560 );
   or U16062 ( n16406,n16383,n15678 );
   nand U16063 ( n16383,n15683,n16407 );
   nand U16064 ( n16407,n15689,n15685 );
   nand U16065 ( n16375,n16377,n16408 );
   nand U16066 ( n16408,n16409,n15783,n16410 );
   nand U16067 ( n16410,n15789,n15784 );
   nand U16068 ( n16363,n14863,n14850 );
   not U16069 ( n15988,n16021 );
   nand U16070 ( n16021,n15992,n16362 );
   nand U16071 ( n16341,n14512,n16345,n14759 );
   not U16072 ( n15361,n15087 );
   nor U16073 ( n15087,n16411,n15089 );
   nand U16074 ( n16255,n15384,n14503 );
   not U16075 ( n14733,n14766 );
   nand U16076 ( n16254,n15082,n14731 );
   nor U16077 ( n14731,n15083,n16412 );
   and U16078 ( n16412,n16413,n14734 );
   nand U16079 ( n16413,n16247,n16216 );
   nand U16080 ( n16417,p1_reg2_reg_30_,n15089 );
   nand U16081 ( n16415,n14708,n14709,n15082 );
   nand U16082 ( n14708,n14706,n16418 );
   nand U16083 ( n16418,n15083,n15084 );
   nand U16084 ( n16414,n15088,n14706 );
   nand U16085 ( n16421,p1_reg2_reg_31_,n15089 );
   nand U16086 ( n16416,n14707,n15090 );
   nor U16087 ( n14707,n15108,n16422 );
   and U16088 ( n15108,n16423,n16424 );
   nand U16089 ( n16424,n14766,n16425 );
   nand U16090 ( n16423,n16427,n16428 );
   nand U16091 ( n16420,n15082,n14700 );
   xor U16092 ( n14700,n14697,n14709 );
   nand U16093 ( n14709,n15084,n16429,n15083 );
   nor U16094 ( n15083,n14746,n14734,n16194 );
   not U16095 ( n16194,n16247 );
   nor U16096 ( n16247,n14771,n14759,n16134 );
   not U16097 ( n16134,n16162 );
   nor U16098 ( n16162,n14782,n14794,n16061 );
   not U16099 ( n16061,n16106 );
   nor U16100 ( n16106,n14819,n16064,n15979 );
   not U16101 ( n15979,n16031 );
   nor U16102 ( n16031,n15953,n15982,n15933 );
   not U16103 ( n15933,n15983 );
   nor U16104 ( n15983,n14864,n15936,n15877 );
   not U16105 ( n15877,n15908 );
   nor U16106 ( n15908,n14875,n15835,n15811 );
   not U16107 ( n15811,n15880 );
   nor U16108 ( n15880,n14909,n15814,n15750 );
   not U16109 ( n15750,n15779 );
   nor U16110 ( n15779,n14932,n15753,n15675 );
   not U16111 ( n15675,n15731 );
   nor U16112 ( n15731,n15678,n15646,n15623 );
   not U16113 ( n15623,n15679 );
   nor U16114 ( n15679,n14978,n14966,n15545 );
   not U16115 ( n15545,n15581 );
   nor U16116 ( n15581,n15002,n14990,n15465 );
   not U16117 ( n15465,n15508 );
   nor U16118 ( n15508,n15468,n15443,n15421 );
   not U16119 ( n15421,n15469 );
   nor U16120 ( n15469,n15385,n15056,n15036 );
   not U16121 ( n15084,n14719 );
   nand U16122 ( n16419,n15088,n14697 );
   nor U16123 ( n15088,n16431,n15089 );
   nand U16124 ( n16432,n16264,n16433 );
   nand U16125 ( n16433,n15064,n15060,n16434,n15059 );
   nor U16126 ( n16438,n16439,n16440 );
   and U16127 ( n16439,p1_addr_reg_19_,n16441 );
   nand U16128 ( n16437,n16442,n16443 );
   nand U16129 ( n16436,n16444,n16445,n16446 );
   nand U16130 ( n16445,n16447,n16448,n16449 );
   xor U16131 ( n16449,p1_reg1_reg_19_,n16443 );
   nand U16132 ( n16448,n16450,n16451 );
   nand U16133 ( n16444,n16450,n16452,n16453 );
   xor U16134 ( n16453,n16454,p1_reg1_reg_19_ );
   nand U16135 ( n16452,p1_reg1_reg_18_,n16447 );
   nand U16136 ( n16447,n16455,n16456 );
   not U16137 ( n16455,n16457 );
   nand U16138 ( n16450,n16458,n16457 );
   nand U16139 ( n16460,n16462,n16463,n16464 );
   xor U16140 ( n16464,n15952,n16454 );
   not U16141 ( n15952,p1_reg2_reg_19_ );
   nand U16142 ( n16463,n16465,n15931 );
   nand U16143 ( n16459,n16465,n16466,n16467 );
   xor U16144 ( n16467,n16454,p1_reg2_reg_19_ );
   nand U16145 ( n16466,p1_reg2_reg_18_,n16462 );
   nand U16146 ( n16462,n16468,n16456 );
   nand U16147 ( n16465,n16458,n16469 );
   nand U16148 ( n16474,n16475,n16476,n16477 );
   nand U16149 ( n16477,n16461,n16478 );
   xor U16150 ( n16478,n16468,p1_reg2_reg_18_ );
   nand U16151 ( n16475,n16446,n16479 );
   xor U16152 ( n16479,n16451,n16457 );
   not U16153 ( n16451,p1_reg1_reg_18_ );
   nand U16154 ( n16472,n16480,n16456 );
   nand U16155 ( n16480,n16481,n16482 );
   nand U16156 ( n16482,n16483,n16446 );
   xor U16157 ( n16483,n16457,p1_reg1_reg_18_ );
   nand U16158 ( n16457,n16484,n16485,n16486 );
   nand U16159 ( n16486,n16487,n16488 );
   nand U16160 ( n16485,p1_reg1_reg_17_,n16489 );
   nand U16161 ( n16489,n16490,n16491 );
   or U16162 ( n16484,n16491,n16490 );
   nand U16163 ( n16481,n16492,n16461 );
   xor U16164 ( n16492,n15931,n16468 );
   not U16165 ( n16468,n16469 );
   nand U16166 ( n16469,n16493,n16494,n16495 );
   nand U16167 ( n16495,n16496,n16497 );
   nand U16168 ( n16494,p1_reg2_reg_17_,n16498 );
   nand U16169 ( n16498,n16490,n16499 );
   or U16170 ( n16493,n16499,n16490 );
   not U16171 ( n15931,p1_reg2_reg_18_ );
   nand U16172 ( n16471,p1_addr_reg_18_,n16441 );
   nand U16173 ( n16470,p1_reg3_reg_18_,p1_u3084 );
   nor U16174 ( n16503,n16504,n16505 );
   nor U16175 ( n16504,n16506,n16507 );
   nand U16176 ( n16502,n16442,n16508 );
   nand U16177 ( n16501,n16509,n16510,n16446 );
   nand U16178 ( n16510,n16511,n16512,n16488 );
   and U16179 ( n16488,n16513,n16514 );
   or U16180 ( n16513,n16508,p1_reg1_reg_17_ );
   nand U16181 ( n16512,n16515,n16491 );
   nand U16182 ( n16511,n16508,p1_reg1_reg_17_ );
   nand U16183 ( n16509,n16516,n16491,n16517 );
   xor U16184 ( n16517,p1_reg1_reg_17_,n16490 );
   nand U16185 ( n16491,n16518,p1_reg1_reg_16_ );
   nand U16186 ( n16516,n16487,n16514 );
   nand U16187 ( n16514,n16519,n16520 );
   nand U16188 ( n16522,n16523,n16524,n16497 );
   and U16189 ( n16497,n16525,n16526 );
   nand U16190 ( n16525,n16490,n15907 );
   nand U16191 ( n16524,n16527,n16499 );
   nand U16192 ( n16523,n16508,p1_reg2_reg_17_ );
   nand U16193 ( n16521,n16528,n16499,n16529 );
   xor U16194 ( n16529,n15907,n16508 );
   not U16195 ( n15907,p1_reg2_reg_17_ );
   nand U16196 ( n16499,n16518,p1_reg2_reg_16_ );
   nand U16197 ( n16528,n16496,n16526 );
   nand U16198 ( n16526,n16519,n15875 );
   nand U16199 ( n16534,n16535,n16536 );
   nand U16200 ( n16536,n16446,n16537 );
   xor U16201 ( n16537,n16487,p1_reg1_reg_16_ );
   nand U16202 ( n16535,n16461,n16538 );
   xor U16203 ( n16538,n16496,p1_reg2_reg_16_ );
   nand U16204 ( n16532,n16518,n16539 );
   nand U16205 ( n16539,n16540,n16476,n16541 );
   nand U16206 ( n16541,n16542,n16461 );
   xor U16207 ( n16542,n15875,n16496 );
   not U16208 ( n16496,n16527 );
   nand U16209 ( n16527,n16543,n16544 );
   nand U16210 ( n16544,n16545,n15834 );
   or U16211 ( n16545,n16546,n16547 );
   nand U16212 ( n16543,n16546,n16547 );
   not U16213 ( n15875,p1_reg2_reg_16_ );
   nand U16214 ( n16540,n16548,n16446 );
   xor U16215 ( n16548,n16520,n16487 );
   not U16216 ( n16487,n16515 );
   nand U16217 ( n16515,n16549,n16550 );
   nand U16218 ( n16550,n16551,n16552 );
   or U16219 ( n16551,n16553,n16547 );
   nand U16220 ( n16549,n16553,n16547 );
   not U16221 ( n16520,p1_reg1_reg_16_ );
   nand U16222 ( n16531,p1_addr_reg_16_,n16441 );
   nand U16223 ( n16530,p1_reg3_reg_16_,p1_u3084 );
   nand U16224 ( n16559,n16560,n16476,n16561 );
   nand U16225 ( n16561,n16562,n16461 );
   xor U16226 ( n16562,p1_reg2_reg_15_,n16546 );
   nand U16227 ( n16560,n16563,n16446 );
   xor U16228 ( n16563,p1_reg1_reg_15_,n16553 );
   nand U16229 ( n16556,n16564,n16547 );
   nand U16230 ( n16564,n16565,n16566 );
   nand U16231 ( n16566,n16446,n16567 );
   xor U16232 ( n16567,n16553,n16552 );
   not U16233 ( n16552,p1_reg1_reg_15_ );
   nand U16234 ( n16553,n16568,n16569 );
   nand U16235 ( n16569,n16570,n16571 );
   or U16236 ( n16570,n16572,n16573 );
   nand U16237 ( n16568,n16573,n16572 );
   nand U16238 ( n16565,n16461,n16574 );
   xor U16239 ( n16574,n16546,n15834 );
   not U16240 ( n15834,p1_reg2_reg_15_ );
   nand U16241 ( n16546,n16575,n16576 );
   nand U16242 ( n16576,n16577,n15809 );
   or U16243 ( n16577,n16578,n16573 );
   nand U16244 ( n16575,n16573,n16578 );
   nand U16245 ( n16555,p1_addr_reg_15_,n16441 );
   nand U16246 ( n16554,p1_reg3_reg_15_,p1_u3084 );
   nand U16247 ( n16583,n16584,n16585 );
   nand U16248 ( n16585,n16446,n16586 );
   xor U16249 ( n16586,n16572,n16571 );
   not U16250 ( n16571,p1_reg1_reg_14_ );
   nand U16251 ( n16584,n16461,n16587 );
   xor U16252 ( n16587,n15809,n16578 );
   not U16253 ( n15809,p1_reg2_reg_14_ );
   nand U16254 ( n16581,n16588,n16589 );
   nand U16255 ( n16589,n16590,n16476,n16591 );
   nand U16256 ( n16591,n16592,n16461 );
   xor U16257 ( n16592,n16578,p1_reg2_reg_14_ );
   nand U16258 ( n16578,n16593,n16594 );
   nand U16259 ( n16593,n16595,n16596,n16597 );
   nand U16260 ( n16590,n16598,n16446 );
   xor U16261 ( n16598,p1_reg1_reg_14_,n16572 );
   nand U16262 ( n16572,n16599,n16600 );
   nand U16263 ( n16599,n16601,n16602,n16603 );
   nand U16264 ( n16580,p1_addr_reg_14_,n16441 );
   nand U16265 ( n16579,p1_reg3_reg_14_,p1_u3084 );
   nor U16266 ( n16607,n16608,n16609 );
   nor U16267 ( n16608,n16506,n16610 );
   nand U16268 ( n16606,n16442,n16611 );
   nand U16269 ( n16605,n16612,n16613,n16446 );
   nand U16270 ( n16613,n16603,n16614,n16615,n16600 );
   or U16271 ( n16600,p1_reg1_reg_13_,n16611 );
   nand U16272 ( n16614,n16616,n16602 );
   nand U16273 ( n16603,n16611,p1_reg1_reg_13_ );
   nand U16274 ( n16612,n16601,n16602,n16617 );
   xor U16275 ( n16617,p1_reg1_reg_13_,n16618 );
   nand U16276 ( n16620,n16597,n16621,n16622,n16594 );
   nand U16277 ( n16594,n15778,n16618 );
   nand U16278 ( n16621,n16623,n16596 );
   nand U16279 ( n16597,n16611,p1_reg2_reg_13_ );
   nand U16280 ( n16619,n16595,n16596,n16624 );
   xor U16281 ( n16624,n15778,n16611 );
   not U16282 ( n15778,p1_reg2_reg_13_ );
   nor U16283 ( n16628,n16629,n16630 );
   nor U16284 ( n16629,n16506,n16631 );
   nand U16285 ( n16627,n16632,n16633 );
   nand U16286 ( n16633,n16634,n16476,n16635 );
   nand U16287 ( n16635,p1_reg2_reg_12_,n16636,n16461 );
   nand U16288 ( n16634,p1_reg1_reg_12_,n16637,n16446 );
   nand U16289 ( n16626,n16638,n16601,n16446 );
   nand U16290 ( n16601,n16615,n16637 );
   nand U16291 ( n16638,n16616,n16639 );
   nand U16292 ( n16639,n16602,n16615 );
   or U16293 ( n16615,n16632,p1_reg1_reg_12_ );
   nand U16294 ( n16602,n16632,p1_reg1_reg_12_ );
   not U16295 ( n16616,n16637 );
   nand U16296 ( n16637,n16640,n16641 );
   nand U16297 ( n16641,n16642,n16643 );
   nand U16298 ( n16643,n16644,n16645 );
   nand U16299 ( n16640,n16646,p1_reg1_reg_11_ );
   nand U16300 ( n16625,n16647,n16595,n16461 );
   nand U16301 ( n16595,n16622,n16636 );
   nand U16302 ( n16647,n16623,n16648 );
   nand U16303 ( n16648,n16596,n16622 );
   nand U16304 ( n16622,n16649,n15748 );
   not U16305 ( n15748,p1_reg2_reg_12_ );
   nand U16306 ( n16596,n16632,p1_reg2_reg_12_ );
   not U16307 ( n16623,n16636 );
   nand U16308 ( n16636,n16650,n16651 );
   nand U16309 ( n16651,n16652,n16653 );
   nand U16310 ( n16653,n16644,n15730 );
   nand U16311 ( n16650,n16646,p1_reg2_reg_11_ );
   nand U16312 ( n16658,n16659,n16660 );
   nand U16313 ( n16660,n16446,n16661 );
   xor U16314 ( n16661,n16642,p1_reg1_reg_11_ );
   nand U16315 ( n16659,n16461,n16662 );
   xor U16316 ( n16662,n16652,p1_reg2_reg_11_ );
   nand U16317 ( n16656,n16646,n16663 );
   nand U16318 ( n16663,n16664,n16476,n16665 );
   nand U16319 ( n16665,n16666,n16461 );
   xor U16320 ( n16666,n15730,n16652 );
   and U16321 ( n16652,n16667,n16668 );
   nand U16322 ( n16667,n16669,n16670,n16671 );
   not U16323 ( n15730,p1_reg2_reg_11_ );
   nand U16324 ( n16664,n16672,n16446 );
   xor U16325 ( n16672,n16645,n16642 );
   and U16326 ( n16642,n16673,n16674 );
   nand U16327 ( n16673,n16675,n16676,n16677 );
   not U16328 ( n16645,p1_reg1_reg_11_ );
   nand U16329 ( n16655,p1_addr_reg_11_,n16441 );
   nand U16330 ( n16654,p1_reg3_reg_11_,p1_u3084 );
   nor U16331 ( n16681,n16682,n16683 );
   nor U16332 ( n16682,n16506,n16684 );
   nand U16333 ( n16680,n16442,n16685 );
   nand U16334 ( n16679,n16686,n16687,n16446 );
   nand U16335 ( n16687,n16677,n16688,n16689,n16674 );
   or U16336 ( n16674,n16685,p1_reg1_reg_10_ );
   nand U16337 ( n16677,n16685,p1_reg1_reg_10_ );
   nand U16338 ( n16686,n16675,n16676,n16690 );
   xor U16339 ( n16690,p1_reg1_reg_10_,n16691 );
   nand U16340 ( n16675,n16689,n16692 );
   nand U16341 ( n16694,n16671,n16695,n16696,n16668 );
   nand U16342 ( n16668,n16691,n15674 );
   nand U16343 ( n16671,n16685,p1_reg2_reg_10_ );
   nand U16344 ( n16693,n16669,n16670,n16697 );
   xor U16345 ( n16697,n15674,n16685 );
   not U16346 ( n15674,p1_reg2_reg_10_ );
   nand U16347 ( n16669,n16696,n16698 );
   nor U16348 ( n16702,n16703,n16704 );
   nor U16349 ( n16703,n16506,n16705 );
   nand U16350 ( n16701,n16706,n16707 );
   nand U16351 ( n16707,n16708,n16476,n16709 );
   nand U16352 ( n16709,p1_reg2_reg_9_,n16698,n16461 );
   nand U16353 ( n16708,p1_reg1_reg_9_,n16692,n16446 );
   nand U16354 ( n16700,n16710,n16711,n16446 );
   nand U16355 ( n16711,n16712,n16713 );
   nand U16356 ( n16710,n16688,n16689 );
   not U16357 ( n16689,n16712 );
   nor U16358 ( n16712,n16706,p1_reg1_reg_9_ );
   nand U16359 ( n16688,n16713,n16676 );
   nand U16360 ( n16676,n16706,p1_reg1_reg_9_ );
   not U16361 ( n16713,n16692 );
   nand U16362 ( n16692,n16714,n16715 );
   nand U16363 ( n16714,n16716,n16717 );
   nand U16364 ( n16699,n16718,n16719,n16461 );
   nand U16365 ( n16719,n16720,n16721 );
   nand U16366 ( n16718,n16695,n16696 );
   not U16367 ( n16696,n16720 );
   nor U16368 ( n16720,n16706,p1_reg2_reg_9_ );
   nand U16369 ( n16695,n16721,n16670 );
   nand U16370 ( n16670,n16706,p1_reg2_reg_9_ );
   not U16371 ( n16721,n16698 );
   nand U16372 ( n16698,n16722,n16723 );
   nand U16373 ( n16722,n16724,n16725 );
   nor U16374 ( n16729,n16730,n16731 );
   nor U16375 ( n16730,n16506,n16732 );
   nand U16376 ( n16728,n16442,n16733 );
   or U16377 ( n16727,n16734,n16735 );
   xor U16378 ( n16734,n16717,n16736 );
   nand U16379 ( n16736,n16716,n16715 );
   nand U16380 ( n16715,n16733,p1_reg1_reg_8_ );
   or U16381 ( n16716,n16733,p1_reg1_reg_8_ );
   nand U16382 ( n16717,n16737,n16738 );
   nand U16383 ( n16738,p1_reg1_reg_7_,n16739 );
   nand U16384 ( n16739,n16740,n16741 );
   nand U16385 ( n16737,n16742,n16743 );
   nand U16386 ( n16726,n16744,n16461 );
   xor U16387 ( n16744,n16745,n16725 );
   nand U16388 ( n16725,n16746,n16747 );
   nand U16389 ( n16747,p1_reg2_reg_7_,n16748 );
   nand U16390 ( n16748,n16749,n16741 );
   nand U16391 ( n16746,n16742,n16750 );
   and U16392 ( n16745,n16723,n16724 );
   nand U16393 ( n16724,n16751,n15621 );
   not U16394 ( n15621,p1_reg2_reg_8_ );
   nand U16395 ( n16723,n16733,p1_reg2_reg_8_ );
   nor U16396 ( n16755,n16756,n16757 );
   nor U16397 ( n16756,n16506,n16758 );
   nand U16398 ( n16754,n16742,n16759 );
   nand U16399 ( n16759,n16760,n16476,n16761 );
   nand U16400 ( n16761,n16762,n15580,n16461 );
   not U16401 ( n15580,p1_reg2_reg_7_ );
   nand U16402 ( n16760,n16763,n16764,n16446 );
   not U16403 ( n16764,p1_reg1_reg_7_ );
   nand U16404 ( n16753,n16765,n16763,n16446 );
   nand U16405 ( n16763,n16766,n16767,n16768 );
   xor U16406 ( n16768,n16742,p1_reg1_reg_7_ );
   nand U16407 ( n16766,n16769,n16770 );
   nand U16408 ( n16765,n16740,n16771 );
   nand U16409 ( n16771,p1_reg1_reg_7_,n16741 );
   not U16410 ( n16740,n16743 );
   nand U16411 ( n16743,n16770,n16772 );
   nand U16412 ( n16752,n16773,n16762,n16461 );
   nand U16413 ( n16762,n16774,n16775,n16776 );
   xor U16414 ( n16776,n16742,p1_reg2_reg_7_ );
   nand U16415 ( n16774,n16777,n16778 );
   nand U16416 ( n16773,n16749,n16779 );
   nand U16417 ( n16779,p1_reg2_reg_7_,n16741 );
   not U16418 ( n16749,n16750 );
   nand U16419 ( n16750,n16778,n16780 );
   nor U16420 ( n16784,n16785,n16786 );
   nor U16421 ( n16785,n16506,n16787 );
   nand U16422 ( n16783,n16788,n16789 );
   nand U16423 ( n16789,n16790,n16476,n16791 );
   nand U16424 ( n16791,p1_reg2_reg_6_,n16792,n16461 );
   nand U16425 ( n16790,p1_reg1_reg_6_,n16793,n16446 );
   nand U16426 ( n16782,n16794,n16772,n16446 );
   nand U16427 ( n16772,n16793,n16767 );
   nand U16428 ( n16794,n16769,n16795 );
   nand U16429 ( n16795,n16770,n16767 );
   or U16430 ( n16767,n16788,p1_reg1_reg_6_ );
   nand U16431 ( n16770,n16788,p1_reg1_reg_6_ );
   not U16432 ( n16769,n16793 );
   nand U16433 ( n16793,n16796,n16797 );
   nand U16434 ( n16797,p1_reg1_reg_5_,n16798 );
   nand U16435 ( n16798,n16799,n16800 );
   nand U16436 ( n16796,n16801,n16802 );
   nand U16437 ( n16781,n16803,n16780,n16461 );
   nand U16438 ( n16780,n16792,n16775 );
   nand U16439 ( n16803,n16777,n16804 );
   nand U16440 ( n16804,n16778,n16775 );
   nand U16441 ( n16775,n16805,n15543 );
   not U16442 ( n15543,p1_reg2_reg_6_ );
   nand U16443 ( n16778,n16788,p1_reg2_reg_6_ );
   not U16444 ( n16777,n16792 );
   nand U16445 ( n16792,n16806,n16807 );
   nand U16446 ( n16807,p1_reg2_reg_5_,n16808 );
   nand U16447 ( n16808,n16809,n16800 );
   nand U16448 ( n16806,n16801,n16810 );
   nor U16449 ( n16814,n16815,n16816 );
   nor U16450 ( n16815,n16506,n16817 );
   nand U16451 ( n16813,n16801,n16818 );
   nand U16452 ( n16818,n16819,n16476,n16820 );
   nand U16453 ( n16820,n16821,n16822,n16446 );
   not U16454 ( n16822,p1_reg1_reg_5_ );
   nand U16455 ( n16819,n16823,n15507,n16461 );
   not U16456 ( n15507,p1_reg2_reg_5_ );
   nand U16457 ( n16812,n16824,n16821,n16446 );
   nand U16458 ( n16821,n16825,n16826,n16827 );
   xor U16459 ( n16827,n16801,p1_reg1_reg_5_ );
   nand U16460 ( n16825,n16828,n16829 );
   nand U16461 ( n16824,n16799,n16830 );
   nand U16462 ( n16830,p1_reg1_reg_5_,n16800 );
   not U16463 ( n16799,n16802 );
   nand U16464 ( n16802,n16829,n16831 );
   nand U16465 ( n16831,n16832,n16826 );
   nand U16466 ( n16811,n16833,n16823,n16461 );
   nand U16467 ( n16823,n16834,n16835,n16836 );
   xor U16468 ( n16836,n16801,p1_reg2_reg_5_ );
   nand U16469 ( n16834,n16837,n16838 );
   nand U16470 ( n16833,n16809,n16839 );
   nand U16471 ( n16839,p1_reg2_reg_5_,n16800 );
   not U16472 ( n16809,n16810 );
   nand U16473 ( n16810,n16838,n16840 );
   nand U16474 ( n16840,n16841,n16835 );
   nor U16475 ( n16848,n16735,n16849,n16850 );
   nor U16476 ( n16850,n16851,n16832 );
   and U16477 ( n16851,n16826,n16829 );
   nand U16478 ( n16829,n16852,p1_reg1_reg_4_ );
   not U16479 ( n16826,n16853 );
   nor U16480 ( n16849,n16853,n16828 );
   not U16481 ( n16828,n16832 );
   nor U16482 ( n16853,n16852,p1_reg1_reg_4_ );
   not U16483 ( n16847,n16854 );
   nor U16484 ( n16846,n16855,n16856,n16857 );
   nor U16485 ( n16857,n16858,n16841 );
   and U16486 ( n16858,n16835,n16838 );
   nand U16487 ( n16838,n16852,p1_reg2_reg_4_ );
   not U16488 ( n16835,n16859 );
   nor U16489 ( n16856,n16859,n16837 );
   not U16490 ( n16837,n16841 );
   nor U16491 ( n16859,n16852,p1_reg2_reg_4_ );
   nand U16492 ( n16844,p1_reg3_reg_4_,p1_u3084 );
   nand U16493 ( n16860,n16861,n16476,n16862 );
   nand U16494 ( n16862,p1_reg1_reg_4_,n16832,n16446 );
   nand U16495 ( n16832,n16863,n16864 );
   nand U16496 ( n16864,p1_reg1_reg_3_,n16865 );
   or U16497 ( n16865,n16866,n16867 );
   nand U16498 ( n16863,n16867,n16866 );
   nand U16499 ( n16861,p1_reg2_reg_4_,n16841,n16461 );
   nand U16500 ( n16841,n16868,n16869 );
   nand U16501 ( n16869,p1_reg2_reg_3_,n16870 );
   or U16502 ( n16870,n16871,n16867 );
   nand U16503 ( n16868,n16867,n16871 );
   nand U16504 ( n16842,p1_addr_reg_4_,n16441 );
   nor U16505 ( n16875,n16876,n16877 );
   nor U16506 ( n16876,n16506,n16878 );
   nand U16507 ( n16874,n16442,n16867 );
   nand U16508 ( n16873,n16446,n16879 );
   xor U16509 ( n16879,n16880,n16867 );
   xor U16510 ( n16880,n16866,p1_reg1_reg_3_ );
   nand U16511 ( n16866,n16881,n16882 );
   nand U16512 ( n16882,n16883,n16884 );
   xor U16513 ( n16885,n16886,n16887 );
   xor U16514 ( n16886,n16871,n15442 );
   not U16515 ( n15442,p1_reg2_reg_3_ );
   nand U16516 ( n16871,n16888,n16889 );
   nand U16517 ( n16889,n16890,n16891 );
   nor U16518 ( n16897,n16506,n16898 );
   nor U16519 ( n16896,n16899,n16476 );
   nor U16520 ( n16895,p1_state_reg,n15397 );
   not U16521 ( n15397,p1_reg3_reg_2_ );
   nand U16522 ( n16893,n16900,n16901,n16461 );
   nand U16523 ( n16901,n16888,n16891,n16890 );
   nand U16524 ( n16891,n16899,n15411 );
   nand U16525 ( n16888,n16902,p1_reg2_reg_2_ );
   nand U16526 ( n16900,n16903,n16904 );
   not U16527 ( n16904,n16890 );
   nand U16528 ( n16890,n16905,n16906 );
   nand U16529 ( n16906,n16907,n16908 );
   xor U16530 ( n16903,n15411,n16902 );
   not U16531 ( n15411,p1_reg2_reg_2_ );
   nand U16532 ( n16854,n16909,n16910,p1_u4006 );
   nand U16533 ( n16910,n16911,n16912,n16426 );
   nand U16534 ( n16912,n16913,n16914 );
   nand U16535 ( n16911,n16915,n16916 );
   nand U16536 ( n16909,n16917,n16918 );
   nand U16537 ( n16917,n16426,n16919 );
   nand U16538 ( n16919,n16913,n16920 );
   nand U16539 ( n16892,n16921,n16922,n16446 );
   nand U16540 ( n16922,n16881,n16884,n16883 );
   or U16541 ( n16884,n16902,p1_reg1_reg_2_ );
   nand U16542 ( n16881,n16902,p1_reg1_reg_2_ );
   nand U16543 ( n16921,n16923,n16924 );
   not U16544 ( n16924,n16883 );
   nand U16545 ( n16883,n16925,n16926 );
   nand U16546 ( n16926,p1_reg1_reg_0_,n16927,p1_ir_reg_0_ );
   xor U16547 ( n16923,p1_reg1_reg_2_,n16899 );
   nor U16548 ( n16931,n16932,n16933 );
   nor U16549 ( n16933,p1_state_reg,n15377 );
   not U16550 ( n15377,p1_reg3_reg_1_ );
   nor U16551 ( n16932,n16506,n16934 );
   nand U16552 ( n16930,n16442,n16935 );
   not U16553 ( n16442,n16476 );
   nand U16554 ( n16929,n16461,n16936 );
   xor U16555 ( n16936,n16937,n16914 );
   not U16556 ( n16914,n16907 );
   nor U16557 ( n16907,n16918,n16920 );
   nand U16558 ( n16937,n16905,n16908 );
   nand U16559 ( n16908,n16938,n15383 );
   not U16560 ( n15383,p1_reg2_reg_1_ );
   nand U16561 ( n16905,n16935,p1_reg2_reg_1_ );
   nand U16562 ( n16928,n16446,n16939 );
   xor U16563 ( n16939,n16940,n16941 );
   nand U16564 ( n16941,n16925,n16927 );
   or U16565 ( n16927,n16935,p1_reg1_reg_1_ );
   nand U16566 ( n16925,n16935,p1_reg1_reg_1_ );
   nand U16567 ( n16940,p1_ir_reg_0_,p1_reg1_reg_0_ );
   nand U16568 ( n16945,p1_ir_reg_0_,n16946 );
   nand U16569 ( n16946,n16947,n16476,n16948 );
   nand U16570 ( n16948,n16461,n16920 );
   not U16571 ( n16920,p1_reg2_reg_0_ );
   nand U16572 ( n16476,n16949,n16275 );
   or U16573 ( n16947,n16735,p1_reg1_reg_0_ );
   nand U16574 ( n16944,n16950,n16918 );
   nand U16575 ( n16950,n16951,n16952 );
   nand U16576 ( n16952,n16446,p1_reg1_reg_0_ );
   nand U16577 ( n16735,n16949,n16915 );
   nand U16578 ( n16951,n16461,p1_reg2_reg_0_ );
   nand U16579 ( n16855,n16913,n16426,n16949 );
   and U16580 ( n16949,n16953,n16506 );
   nand U16581 ( n16953,n16954,n16955 );
   nand U16582 ( n16955,n15061,n16956 );
   nand U16583 ( n16956,n16957,n16430,n16958,n16959 );
   and U16584 ( n16959,n16960,n16431,n16264,n16961 );
   not U16585 ( n16958,n16962 );
   nand U16586 ( n16954,n16963,p1_state_reg );
   not U16587 ( n16441,n16506 );
   nand U16588 ( n16964,n16966,n16967 );
   nand U16589 ( n16942,p1_reg3_reg_0_,p1_u3084 );
   nand U16590 ( n16970,n16971,n16972,n16973 );
   nor U16591 ( n16973,n16974,n16975,n16976,n16977 );
   nor U16592 ( n16977,n16978,n16979,n16980 );
   and U16593 ( n16976,n16978,n16979,n15573 );
   nand U16594 ( n16978,n16981,n16982,n16983,n16984 );
   nor U16595 ( n16984,n16985,n16986,n16987 );
   nor U16596 ( n16987,n16988,n16989 );
   nor U16597 ( n16988,n16990,n16991 );
   nor U16598 ( n16991,n16992,n16993 );
   nor U16599 ( n16990,n16994,n16995 );
   nor U16600 ( n16986,n16996,n16997,n16998,n16999 );
   not U16601 ( n16997,n17000 );
   not U16602 ( n16996,n17001 );
   nor U16603 ( n16985,n17002,n17003 );
   and U16604 ( n17002,n17004,n16422 );
   nand U16605 ( n16983,n17005,n17006 );
   nand U16606 ( n17006,n17007,n17008 );
   nand U16607 ( n17008,n17009,n17010,n17011 );
   nand U16608 ( n17011,n17012,n14512 );
   nand U16609 ( n17009,n17013,n14759 );
   nand U16610 ( n17007,n17014,n17015 );
   nand U16611 ( n16982,n17005,n17016,n17017,n17018 );
   nand U16612 ( n17018,n17019,n17020 );
   nand U16613 ( n17020,n17021,n17022 );
   nand U16614 ( n17019,n17023,n17024 );
   nand U16615 ( n17024,n17025,n17026 );
   nand U16616 ( n17026,n17027,n17028 );
   nand U16617 ( n17025,n17029,n17030 );
   nand U16618 ( n17030,n17031,n17032,n17033 );
   nand U16619 ( n17033,n17034,n17035 );
   nand U16620 ( n17032,n17036,n17037 );
   or U16621 ( n17037,n17035,n17034 );
   and U16622 ( n17034,n17038,n17039 );
   nand U16623 ( n17039,n17013,n14819 );
   nand U16624 ( n17038,n17012,n14527 );
   nand U16625 ( n17035,n17040,n17041 );
   nand U16626 ( n17041,n17042,n17043 );
   nand U16627 ( n17043,n14828,n17044 );
   not U16628 ( n17042,n17045 );
   nand U16629 ( n17040,n17046,n17047 );
   nand U16630 ( n17047,n17044,n17045,n17048 );
   nand U16631 ( n17048,n17012,n15982 );
   nand U16632 ( n17045,n17049,n17050 );
   nand U16633 ( n17050,n17013,n15982 );
   nand U16634 ( n17049,n17012,n14530 );
   nand U16635 ( n17044,n14530,n17013 );
   nand U16636 ( n17046,n17051,n17052 );
   nand U16637 ( n17052,n17053,n17054,n17055,n17056 );
   nand U16638 ( n17056,n17057,n17058 );
   nor U16639 ( n17055,n17059,n17060 );
   nor U16640 ( n17060,n17061,n17062 );
   nor U16641 ( n17059,n17063,n17064,n17065 );
   not U16642 ( n17064,n17066 );
   nand U16643 ( n17054,n17067,n17068,n17069 );
   nand U16644 ( n17053,n17069,n17070,n17071,n17072 );
   nand U16645 ( n17072,n17073,n17074 );
   nand U16646 ( n17074,n17075,n17076 );
   nand U16647 ( n17073,n17077,n17078 );
   nand U16648 ( n17078,n17079,n17080 );
   nand U16649 ( n17080,n17081,n17082 );
   nand U16650 ( n17079,n17083,n17084 );
   nand U16651 ( n17084,n17085,n17086 );
   nand U16652 ( n17083,n17087,n17088,n17089,n17090 );
   nand U16653 ( n17090,n17091,n17092,n17093 );
   nand U16654 ( n17089,n17094,n17091,n17095 );
   nand U16655 ( n17095,n17096,n17097 );
   nand U16656 ( n17097,n17098,n17099,n17100 );
   nor U16657 ( n17100,n17101,n17102,n17103 );
   nor U16658 ( n17103,n17104,n17105 );
   nor U16659 ( n17102,n17106,n17107,n17108 );
   not U16660 ( n17107,n17109 );
   nor U16661 ( n17101,n17110,n17111,n17112 );
   nand U16662 ( n17099,n17113,n17114,n17115,n17116 );
   nand U16663 ( n17116,n17117,n17118,n17119,n17120 );
   nand U16664 ( n17120,n17121,n17122 );
   nand U16665 ( n17119,n17123,n17124 );
   nand U16666 ( n17118,n17125,n17126,n17127,n17128 );
   nor U16667 ( n17128,n17129,n17130,n17131,n17132 );
   nor U16668 ( n17132,n17121,n17122 );
   nor U16669 ( n17131,n17133,n17134 );
   nor U16670 ( n17130,n17012,n15366 );
   nor U16671 ( n17129,n17135,n17013 );
   nand U16672 ( n17117,n17136,n17137 );
   or U16673 ( n17137,n17122,n17121 );
   and U16674 ( n17121,n17138,n17139 );
   nand U16675 ( n17139,n17013,n15002 );
   nand U16676 ( n17138,n17012,n14575 );
   nand U16677 ( n17122,n17140,n17141 );
   nand U16678 ( n17141,n17013,n14575 );
   nand U16679 ( n17140,n17012,n15002 );
   nand U16680 ( n17136,n17142,n17143 );
   nand U16681 ( n17143,n17144,n17127 );
   nand U16682 ( n17127,n17145,n17146 );
   nand U16683 ( n17144,n17147,n17148 );
   nand U16684 ( n17148,n17149,n17125 );
   nand U16685 ( n17125,n17150,n17151 );
   nand U16686 ( n17149,n17152,n17153 );
   nand U16687 ( n17153,n17134,n17126,n17133 );
   and U16688 ( n17133,n17154,n17155 );
   nand U16689 ( n17155,n17013,n15385 );
   nand U16690 ( n17154,n17012,n14587 );
   nand U16691 ( n17126,n17156,n17157 );
   nand U16692 ( n17134,n17158,n17159 );
   nand U16693 ( n17159,n17013,n14587 );
   nand U16694 ( n17158,n17012,n15385 );
   or U16695 ( n17152,n17157,n17156 );
   and U16696 ( n17156,n17160,n17161 );
   nand U16697 ( n17161,n17013,n14584 );
   nand U16698 ( n17160,n17012,n15036 );
   nand U16699 ( n17157,n17162,n17163 );
   nand U16700 ( n17163,n17013,n15036 );
   nand U16701 ( n17162,n17012,n14584 );
   or U16702 ( n17147,n17151,n17150 );
   and U16703 ( n17150,n17164,n17165 );
   nand U16704 ( n17165,n17013,n14581 );
   nand U16705 ( n17164,n17012,n15443 );
   nand U16706 ( n17151,n17166,n17167 );
   nand U16707 ( n17167,n17013,n15443 );
   nand U16708 ( n17166,n17012,n14581 );
   or U16709 ( n17142,n17146,n17145 );
   and U16710 ( n17145,n17168,n17169 );
   nand U16711 ( n17169,n17013,n14578 );
   nand U16712 ( n17168,n17012,n15468 );
   nand U16713 ( n17146,n17170,n17171 );
   nand U16714 ( n17171,n17013,n15468 );
   nand U16715 ( n17170,n17012,n14578 );
   or U16716 ( n17115,n17124,n17123 );
   and U16717 ( n17123,n17172,n17173 );
   nand U16718 ( n17173,n17013,n14990 );
   nand U16719 ( n17172,n17012,n14572 );
   nand U16720 ( n17124,n17174,n17175 );
   nand U16721 ( n17175,n17013,n14572 );
   nand U16722 ( n17174,n17012,n14990 );
   nand U16723 ( n17114,n17111,n17112 );
   nand U16724 ( n17112,n17176,n17177 );
   nand U16725 ( n17177,n17013,n14978 );
   nand U16726 ( n17176,n17012,n14569 );
   and U16727 ( n17111,n17178,n17179 );
   nand U16728 ( n17179,n17013,n14569 );
   nand U16729 ( n17178,n17012,n14978 );
   not U16730 ( n17113,n17110 );
   nand U16731 ( n17110,n17180,n17109 );
   nand U16732 ( n17109,n17104,n17105 );
   nand U16733 ( n17105,n17181,n17182 );
   nand U16734 ( n17182,n17013,n15646 );
   nand U16735 ( n17181,n17012,n14563 );
   and U16736 ( n17104,n17183,n17184 );
   nand U16737 ( n17184,n17013,n14563 );
   nand U16738 ( n17183,n17012,n15646 );
   nand U16739 ( n17180,n17108,n17106 );
   nand U16740 ( n17106,n17185,n17186 );
   nand U16741 ( n17186,n17013,n14966 );
   nand U16742 ( n17185,n17012,n14566 );
   and U16743 ( n17108,n17187,n17188 );
   nand U16744 ( n17188,n17013,n14566 );
   nand U16745 ( n17187,n17012,n14966 );
   nand U16746 ( n17098,n17189,n17190 );
   or U16747 ( n17096,n17190,n17189 );
   and U16748 ( n17189,n17191,n17192 );
   nand U16749 ( n17192,n15678,n17013 );
   nand U16750 ( n17191,n17012,n14560 );
   nand U16751 ( n17190,n17193,n17194 );
   nand U16752 ( n17194,n17013,n14560 );
   nand U16753 ( n17193,n17012,n15678 );
   nand U16754 ( n17091,n17195,n17196 );
   or U16755 ( n17094,n17092,n17093 );
   and U16756 ( n17093,n17197,n17198 );
   nand U16757 ( n17198,n17013,n14557 );
   nand U16758 ( n17197,n17012,n14932 );
   nand U16759 ( n17092,n17199,n17200 );
   nand U16760 ( n17200,n17013,n14932 );
   nand U16761 ( n17199,n17012,n14557 );
   or U16762 ( n17088,n17196,n17195 );
   and U16763 ( n17195,n17201,n17202 );
   nand U16764 ( n17202,n17013,n15753 );
   nand U16765 ( n17201,n17012,n14554 );
   nand U16766 ( n17196,n17203,n17204 );
   nand U16767 ( n17204,n17013,n14554 );
   nand U16768 ( n17203,n17012,n15753 );
   or U16769 ( n17087,n17086,n17085 );
   and U16770 ( n17085,n17205,n17206 );
   nand U16771 ( n17206,n17013,n14909 );
   nand U16772 ( n17205,n17012,n14551 );
   nand U16773 ( n17086,n17207,n17208 );
   nand U16774 ( n17208,n17013,n14551 );
   nand U16775 ( n17207,n17012,n14909 );
   or U16776 ( n17077,n17082,n17081 );
   and U16777 ( n17081,n17209,n17210 );
   nand U16778 ( n17210,n17013,n14548 );
   nand U16779 ( n17209,n17012,n15814 );
   nand U16780 ( n17082,n17211,n17212 );
   nand U16781 ( n17212,n17013,n15814 );
   nand U16782 ( n17211,n17012,n14548 );
   or U16783 ( n17071,n17076,n17075 );
   and U16784 ( n17075,n17213,n17214 );
   nand U16785 ( n17214,n17013,n14545 );
   nand U16786 ( n17213,n17012,n15835 );
   nand U16787 ( n17076,n17215,n17216 );
   nand U16788 ( n17216,n17013,n15835 );
   nand U16789 ( n17215,n17012,n14545 );
   or U16790 ( n17070,n17068,n17067 );
   and U16791 ( n17067,n17217,n17218 );
   nand U16792 ( n17218,n17013,n14542 );
   nand U16793 ( n17217,n17012,n14875 );
   nand U16794 ( n17068,n17219,n17220 );
   nand U16795 ( n17220,n17013,n14875 );
   nand U16796 ( n17219,n17012,n14542 );
   and U16797 ( n17069,n17221,n17066 );
   nand U16798 ( n17066,n17061,n17062 );
   nand U16799 ( n17062,n17222,n17223 );
   nand U16800 ( n17223,n17013,n14536 );
   nand U16801 ( n17222,n17012,n15936 );
   and U16802 ( n17061,n17224,n17225 );
   nand U16803 ( n17225,n17013,n15936 );
   nand U16804 ( n17224,n17012,n14536 );
   nand U16805 ( n17221,n17065,n17063 );
   nand U16806 ( n17063,n17226,n17227 );
   nand U16807 ( n17227,n17013,n14539 );
   nand U16808 ( n17226,n17012,n14864 );
   and U16809 ( n17065,n17228,n17229 );
   nand U16810 ( n17229,n17013,n14864 );
   nand U16811 ( n17228,n17012,n14539 );
   or U16812 ( n17051,n17058,n17057 );
   and U16813 ( n17057,n17230,n17231 );
   nand U16814 ( n17231,n17013,n14533 );
   nand U16815 ( n17230,n17012,n15953 );
   nand U16816 ( n17058,n17232,n17233 );
   nand U16817 ( n17233,n17013,n15953 );
   nand U16818 ( n17232,n17012,n14533 );
   nand U16819 ( n17036,n17234,n17235 );
   nand U16820 ( n17235,n17013,n14527 );
   nand U16821 ( n17234,n17012,n14819 );
   nand U16822 ( n17031,n17236,n17237 );
   or U16823 ( n17029,n17237,n17236 );
   and U16824 ( n17236,n17238,n17239 );
   nand U16825 ( n17239,n17013,n16064 );
   nand U16826 ( n17238,n17012,n14524 );
   nand U16827 ( n17237,n17240,n17241 );
   nand U16828 ( n17241,n17013,n14524 );
   nand U16829 ( n17240,n17012,n16064 );
   or U16830 ( n17023,n17028,n17027 );
   and U16831 ( n17027,n17242,n17243 );
   nand U16832 ( n17243,n17013,n14794 );
   nand U16833 ( n17242,n17012,n14521 );
   nand U16834 ( n17028,n17244,n17245 );
   nand U16835 ( n17245,n17013,n14521 );
   nand U16836 ( n17244,n17012,n14794 );
   or U16837 ( n17017,n17022,n17021 );
   and U16838 ( n17021,n17246,n17247 );
   nand U16839 ( n17247,n17013,n14782 );
   nand U16840 ( n17246,n17012,n14518 );
   nand U16841 ( n17022,n17248,n17249 );
   nand U16842 ( n17249,n17013,n14518 );
   nand U16843 ( n17248,n17012,n14782 );
   or U16844 ( n17016,n17015,n17014 );
   and U16845 ( n17014,n17250,n17251 );
   nand U16846 ( n17251,n17013,n14771 );
   nand U16847 ( n17250,n17012,n14515 );
   nand U16848 ( n17015,n17252,n17253 );
   nand U16849 ( n17253,n17013,n14515 );
   nand U16850 ( n17252,n17012,n14771 );
   and U16851 ( n17005,n17254,n17255,n17256 );
   not U16852 ( n17256,n16989 );
   nand U16853 ( n16989,n17257,n17258,n17000,n17001 );
   nand U16854 ( n17000,n17259,n17260,n17261 );
   nand U16855 ( n17261,n17012,n14706 );
   nand U16856 ( n17258,n16994,n16995 );
   nand U16857 ( n16995,n17262,n17263 );
   nand U16858 ( n17263,n17013,n14734 );
   nand U16859 ( n17262,n17012,n14506 );
   and U16860 ( n16994,n17264,n17265 );
   nand U16861 ( n17265,n17013,n14506 );
   nand U16862 ( n17264,n17012,n14734 );
   nand U16863 ( n17257,n16998,n16999 );
   nand U16864 ( n16999,n17266,n17267 );
   nand U16865 ( n17267,n17013,n14719 );
   nand U16866 ( n17266,n17012,n14503 );
   and U16867 ( n16998,n17268,n17269 );
   nand U16868 ( n17269,n17012,n14719 );
   nand U16869 ( n17268,n17013,n14503 );
   nand U16870 ( n17255,n17270,n17271,n17272 );
   not U16871 ( n17272,n17010 );
   nand U16872 ( n17010,n17273,n17274 );
   nand U16873 ( n17274,n17013,n14512 );
   nand U16874 ( n17273,n17012,n14759 );
   nand U16875 ( n17271,n16172,n17013 );
   nand U16876 ( n17270,n17012,n16234 );
   nand U16877 ( n17254,n16992,n16993 );
   nand U16878 ( n16993,n17275,n17276 );
   nand U16879 ( n17276,n17013,n14746 );
   nand U16880 ( n17275,n17012,n14509 );
   and U16881 ( n16992,n17277,n17278 );
   nand U16882 ( n17278,n17013,n14509 );
   nand U16883 ( n17277,n17012,n14746 );
   nand U16884 ( n16981,n17279,n17001,n17280 );
   not U16885 ( n17280,n17259 );
   nand U16886 ( n17259,n17281,n17282 );
   nand U16887 ( n17282,n14500,n14497,n17012 );
   nand U16888 ( n17281,n17013,n14706 );
   nand U16889 ( n17001,n17004,n17003,n17283 );
   nand U16890 ( n17283,n17012,n14497 );
   nand U16891 ( n17003,n17284,n17285 );
   nand U16892 ( n17285,n17013,n14497 );
   nand U16893 ( n17284,n17012,n14697 );
   nand U16894 ( n17004,n14697,n17013 );
   nand U16895 ( n17279,n16429,n17260 );
   nand U16896 ( n17260,n14500,n14497,n17013 );
   nor U16897 ( n16975,n17286,n17287,n17288 );
   nor U16898 ( n16974,n17289,n17290,n16454 );
   nand U16899 ( n16972,n17291,n17292 );
   nand U16900 ( n17292,n17293,n17294 );
   nand U16901 ( n17294,n17295,n17296,n17297,n17298 );
   nor U16902 ( n17298,n17299,n16274 );
   nor U16903 ( n17299,n17300,n17301,n17302 );
   nor U16904 ( n17301,n16429,n14497 );
   not U16905 ( n16429,n14706 );
   nand U16906 ( n17300,n17303,n15102,n17304 );
   nand U16907 ( n17303,n17305,n17306 );
   nand U16908 ( n17306,n17307,n16281 );
   not U16909 ( n16281,n16340 );
   nand U16910 ( n17307,n16338,n17308 );
   nand U16911 ( n17308,n17309,n16246 );
   nand U16912 ( n17309,n17310,n16189,n17311 );
   nand U16913 ( n17311,n17312,n16282 );
   nand U16914 ( n17312,n17313,n17314 );
   nand U16915 ( n17310,n17315,n16282,n17316 );
   nand U16916 ( n17315,n17317,n16053 );
   not U16917 ( n16053,n16090 );
   nand U16918 ( n17317,n17318,n17319 );
   nand U16919 ( n17319,n17320,n17321 );
   nand U16920 ( n17321,n15858,n16300,n17322,n17323 );
   nor U16921 ( n17323,n17324,n17325 );
   nor U16922 ( n17324,n17326,n15829 );
   nand U16923 ( n17322,n15859,n17327 );
   nand U16924 ( n17327,n15806,n17328 );
   nand U16925 ( n17328,n17329,n17330,n17331 );
   and U16926 ( n17331,n16314,n15807,n17332 );
   nand U16927 ( n17332,n14918,n16312,n14554 );
   nand U16928 ( n17330,n17333,n15729,n17334,n16315 );
   nor U16929 ( n17334,n15727,n17335 );
   nand U16930 ( n17333,n17336,n15670 );
   not U16931 ( n15670,n15725 );
   nand U16932 ( n17336,n15643,n17337 );
   nand U16933 ( n17337,n17338,n15644 );
   nand U16934 ( n17338,n17339,n16325,n17340 );
   nand U16935 ( n17340,n17341,n17342,n17343 );
   nand U16936 ( n17341,n17344,n17345 );
   nand U16937 ( n17345,n15409,n15407,n17346 );
   nand U16938 ( n15409,n17347,n17348 );
   nand U16939 ( n17348,n17135,n17349 );
   nand U16940 ( n17339,n17343,n17350 );
   nand U16941 ( n17350,n17351,n15502 );
   nand U16942 ( n17351,n17342,n17352 );
   nand U16943 ( n17352,n17353,n16329,n17354 );
   not U16944 ( n17353,n16328 );
   or U16945 ( n17342,n16328,n15542,n15503 );
   not U16946 ( n15542,n16329 );
   and U16947 ( n17343,n16326,n17355 );
   or U16948 ( n17355,n16330,n16328 );
   or U16949 ( n17329,n17356,n17335 );
   nor U16950 ( n15859,n17326,n15863 );
   nand U16951 ( n17296,n14497,n17357,n17358 );
   nand U16952 ( n17295,n17359,n17357,n17360 );
   nand U16953 ( n17359,n14706,n17361 );
   nand U16954 ( n17361,n14500,n14497 );
   nand U16955 ( n17293,n17287,n17362 );
   and U16956 ( n17287,n17363,n17364,n17365,n17366 );
   nor U16957 ( n17366,n17367,n17368,n17369,n17370 );
   or U16958 ( n17370,n15440,n17302,n15505,n15578 );
   xor U16959 ( n15578,n14989,n15558 );
   xor U16960 ( n15505,n15456,n15481 );
   xor U16961 ( n15440,n16401,n15022 );
   or U16962 ( n17369,n15672,n15804,n15832,n16055 );
   xor U16963 ( n16055,n14818,n14804 );
   xor U16964 ( n15832,n15874,n14884 );
   xor U16965 ( n15804,n14908,n14895 );
   xor U16966 ( n15672,n15707,n14941 );
   nand U16967 ( n17368,n16100,n16285,n15116,n17297 );
   not U16968 ( n15116,n15103 );
   nand U16969 ( n15103,n17371,n17304 );
   nand U16970 ( n17304,n14732,n14719 );
   not U16971 ( n16285,n16278 );
   xor U16972 ( n16278,n14745,n16262 );
   not U16973 ( n16262,n14734 );
   xor U16974 ( n16100,n14521,n16073 );
   nand U16975 ( n17367,n15382,n15410,n15464,n15549 );
   nand U16976 ( n15549,n15588,n15585 );
   nand U16977 ( n15585,n14990,n14572 );
   nand U16978 ( n15588,n15001,n15521 );
   not U16979 ( n15464,n15471 );
   nor U16980 ( n15471,n15512,n15511 );
   nor U16981 ( n15511,n14578,n15468 );
   nor U16982 ( n15512,n15011,n17372 );
   nand U16983 ( n15410,n15447,n16403 );
   nand U16984 ( n16403,n15036,n14584 );
   nand U16985 ( n15447,n17373,n15396 );
   nand U16986 ( n15382,n17374,n17375 );
   nand U16987 ( n17375,n15356,n15045 );
   not U16988 ( n17374,n15418 );
   nor U16989 ( n15418,n15356,n15045 );
   nor U16990 ( n17365,n17376,n17377,n16240,n16191 );
   not U16991 ( n16191,n16201 );
   nand U16992 ( n16201,n16252,n16251 );
   nand U16993 ( n16251,n14759,n14512 );
   nand U16994 ( n16252,n16234,n16172 );
   not U16995 ( n16240,n16233 );
   nand U16996 ( n16233,n16344,n16345 );
   nand U16997 ( n16345,n14758,n16216 );
   nand U16998 ( n16344,n14509,n14746 );
   nand U16999 ( n17377,n15360,n15860,n17378 );
   nand U17000 ( n15860,n15914,n15912 );
   nand U17001 ( n15912,n14875,n14542 );
   nand U17002 ( n15914,n15901,n15846 );
   not U17003 ( n15846,n14875 );
   nand U17004 ( n15360,n17379,n15387 );
   nand U17005 ( n15387,n15056,n14590 );
   or U17006 ( n17379,n14590,n15056 );
   nand U17007 ( n17376,n15977,n16023,n16131,n16159 );
   nand U17008 ( n16159,n16200,n16203 );
   nand U17009 ( n16203,n17380,n16146 );
   nand U17010 ( n16200,n14771,n14515 );
   nand U17011 ( n16131,n16205,n16207 );
   nand U17012 ( n16207,n14782,n14518 );
   nand U17013 ( n16205,n14793,n16116 );
   nand U17014 ( n16023,n16355,n16357 );
   nand U17015 ( n16357,n17381,n16001 );
   nand U17016 ( n16355,n14527,n14819 );
   nand U17017 ( n15977,n15987,n16362 );
   nand U17018 ( n16362,n16012,n14828 );
   nand U17019 ( n15987,n15982,n14530 );
   nor U17020 ( n17364,n15950,n15929,n15915,n15787 );
   not U17021 ( n15787,n15775 );
   nand U17022 ( n15775,n16409,n16377 );
   nand U17023 ( n16377,n17382,n15762 );
   nand U17024 ( n16409,n14551,n14909 );
   not U17025 ( n15915,n15904 );
   nand U17026 ( n15904,n16367,n16364 );
   nand U17027 ( n16364,n14864,n14539 );
   nand U17028 ( n16367,n17383,n15890 );
   nor U17029 ( n15929,n16036,n17384 );
   nor U17030 ( n17384,n14536,n15936 );
   nor U17031 ( n16036,n14863,n14850 );
   and U17032 ( n15950,n15990,n15992 );
   nand U17033 ( n15992,n15976,n14839 );
   not U17034 ( n15990,n16361 );
   nor U17035 ( n16361,n14839,n15976 );
   nor U17036 ( n17363,n15747,n15733,n15641,n15627 );
   nor U17037 ( n15627,n15689,n17385 );
   nor U17038 ( n17385,n14566,n14966 );
   nor U17039 ( n15689,n15598,n14977 );
   and U17040 ( n15641,n15683,n15685 );
   nand U17041 ( n15685,n14965,n14952 );
   nand U17042 ( n15683,n14563,n15646 );
   nor U17043 ( n15733,n15789,n17386 );
   nor U17044 ( n17386,n14557,n14932 );
   nor U17045 ( n15789,n15698,n16379 );
   and U17046 ( n15747,n15783,n15784 );
   nand U17047 ( n15784,n14931,n14918 );
   not U17048 ( n14918,n15753 );
   nand U17049 ( n15783,n14554,n15753 );
   nand U17050 ( n16971,n17290,n15066 );
   and U17051 ( n17290,n17297,n17387 );
   nand U17052 ( n17387,n17388,n17389,n17390 );
   not U17053 ( n17390,n17302 );
   nand U17054 ( n17302,n17357,n17391 );
   nand U17055 ( n17391,n15107,n14706 );
   or U17056 ( n17357,n14697,n16422 );
   nand U17057 ( n17389,n14719,n17378,n14732 );
   nand U17058 ( n17388,n17392,n17393,n17371,n17378 );
   not U17059 ( n17378,n17358 );
   nor U17060 ( n17358,n14706,n15107 );
   not U17061 ( n15107,n14500 );
   nand U17062 ( n14500,n17394,n17395,n17396 );
   nand U17063 ( n17396,p1_reg2_reg_30_,n17397 );
   nand U17064 ( n17395,p1_reg0_reg_30_,n17398 );
   nand U17065 ( n17394,p1_reg1_reg_30_,n17399 );
   nand U17066 ( n14706,n17400,n17401 );
   nand U17067 ( n17401,n17402,n11410 );
   not U17068 ( n11410,n13553 );
   xor U17069 ( n13553,n17403,n17404 );
   nand U17070 ( n17404,n17405,n17406 );
   nand U17071 ( n17400,n17407,p2_datao_reg_30_ );
   not U17072 ( n17371,n17360 );
   nor U17073 ( n17360,n14719,n14732 );
   not U17074 ( n14732,n14503 );
   nand U17075 ( n14719,n17408,n17409 );
   nand U17076 ( n17409,n17402,n11400 );
   xor U17077 ( n11400,n17410,n17411 );
   and U17078 ( n17410,n17412,n17413 );
   nand U17079 ( n17408,n17407,p2_datao_reg_29_ );
   nand U17080 ( n17393,n17414,n17415 );
   nand U17081 ( n17415,n17416,n17313,n17314,n17417 );
   nand U17082 ( n17417,n16105,n16289,n16090 );
   nor U17083 ( n16090,n16064,n14818 );
   not U17084 ( n14818,n14524 );
   nand U17085 ( n17314,n16289,n14521,n16073 );
   and U17086 ( n17313,n16291,n16288 );
   nand U17087 ( n16288,n16146,n14515 );
   nand U17088 ( n16291,n16116,n14518 );
   nand U17089 ( n17392,n17414,n17316,n17318,n17418 );
   nand U17090 ( n17418,n17320,n17419 );
   nand U17091 ( n17419,n17420,n16300 );
   nand U17092 ( n17420,n17421,n17422 );
   nand U17093 ( n17422,n17326,n17423 );
   nor U17094 ( n17326,n14875,n15901 );
   nand U17095 ( n17421,n17423,n17424,n15858,n15829 );
   not U17096 ( n15829,n15861 );
   nor U17097 ( n15861,n14545,n14884 );
   not U17098 ( n14884,n15835 );
   nand U17099 ( n15858,n15901,n14875 );
   nand U17100 ( n17424,n17425,n15830 );
   not U17101 ( n15830,n15863 );
   nor U17102 ( n15863,n15835,n15874 );
   nand U17103 ( n17425,n15806,n17426 );
   nand U17104 ( n17426,n17427,n15807 );
   nand U17105 ( n15807,n14895,n14548 );
   not U17106 ( n14895,n15814 );
   nand U17107 ( n17427,n17428,n16312 );
   not U17108 ( n16312,n17335 );
   nor U17109 ( n17335,n14551,n15762 );
   nand U17110 ( n17428,n16314,n17356,n17429,n17430 );
   nor U17111 ( n17430,n17431,n17432 );
   nor U17112 ( n17432,n14931,n15753 );
   and U17113 ( n17431,n15725,n16315,n15729 );
   nor U17114 ( n15725,n15678,n15707 );
   nand U17115 ( n17429,n16323,n17433,n17434,n16315 );
   nand U17116 ( n17434,n16326,n17435,n15644,n16330 );
   nand U17117 ( n16330,n15521,n14572 );
   not U17118 ( n15521,n14990 );
   nand U17119 ( n17435,n17436,n16329 );
   nand U17120 ( n16329,n15001,n14990 );
   nand U17121 ( n17436,n15503,n17437 );
   nand U17122 ( n17437,n17354,n17344,n17438,n15502 );
   not U17123 ( n15502,n15537 );
   nor U17124 ( n15537,n14575,n15481 );
   nand U17125 ( n17438,n17346,n17349,n17439,n15407 );
   nand U17126 ( n15407,n15396,n14584 );
   nand U17127 ( n17439,n17347,n15366,n17440 );
   nand U17128 ( n17440,n17441,n15367 );
   nand U17129 ( n15367,n15358,n14590 );
   not U17130 ( n15366,n17135 );
   nor U17131 ( n17135,n14590,n15358 );
   not U17132 ( n15358,n15056 );
   nand U17133 ( n17347,n15356,n15385 );
   nand U17134 ( n17349,n15045,n14587 );
   not U17135 ( n15045,n15385 );
   nand U17136 ( n17344,n15419,n17346 );
   and U17137 ( n17346,n15462,n17442 );
   nand U17138 ( n17442,n15022,n14581 );
   not U17139 ( n15022,n15443 );
   nor U17140 ( n15419,n14584,n15396 );
   not U17141 ( n15396,n15036 );
   and U17142 ( n17354,n15461,n17443 );
   nand U17143 ( n17443,n15443,n15462,n16401 );
   nand U17144 ( n15462,n15011,n14578 );
   not U17145 ( n15011,n15468 );
   nand U17146 ( n15461,n17372,n15468 );
   nand U17147 ( n15503,n15481,n14575 );
   not U17148 ( n15481,n15002 );
   and U17149 ( n16326,n17444,n15577 );
   not U17150 ( n15577,n15619 );
   nor U17151 ( n15619,n14978,n14989 );
   nand U17152 ( n17433,n17445,n15644 );
   nand U17153 ( n15644,n14952,n14563 );
   not U17154 ( n14952,n15646 );
   nand U17155 ( n17445,n16325,n17446 );
   nand U17156 ( n17446,n16328,n17444 );
   nand U17157 ( n17444,n15598,n14566 );
   not U17158 ( n15598,n14966 );
   nor U17159 ( n16328,n14569,n15558 );
   not U17160 ( n15558,n14978 );
   nand U17161 ( n16325,n14977,n14966 );
   and U17162 ( n16323,n15729,n15669,n15643 );
   nand U17163 ( n15643,n14965,n15646 );
   not U17164 ( n14965,n14563 );
   not U17165 ( n15669,n15727 );
   nor U17166 ( n15727,n14560,n14941 );
   not U17167 ( n14941,n15678 );
   nand U17168 ( n15729,n16379,n14932 );
   nand U17169 ( n17356,n16315,n14557,n15698 );
   nand U17170 ( n16315,n14931,n15753 );
   not U17171 ( n14931,n14554 );
   nand U17172 ( n16314,n15762,n14551 );
   nand U17173 ( n15806,n14908,n15814 );
   not U17174 ( n14908,n14548 );
   not U17175 ( n17423,n17325 );
   nand U17176 ( n17325,n16303,n16306 );
   nand U17177 ( n16306,n17383,n14864 );
   and U17178 ( n17320,n17447,n16028,n17448 );
   nand U17179 ( n17448,n14828,n14530 );
   not U17180 ( n14828,n15982 );
   nand U17181 ( n17447,n17449,n16300 );
   nand U17182 ( n16300,n15976,n15953 );
   nand U17183 ( n17449,n17450,n16302,n16305 );
   nand U17184 ( n16305,n14850,n14536 );
   not U17185 ( n14850,n15936 );
   nand U17186 ( n16302,n14839,n14533 );
   nand U17187 ( n17450,n16337,n16303 );
   nand U17188 ( n16303,n14863,n15936 );
   not U17189 ( n14863,n14536 );
   nor U17190 ( n16337,n14864,n17383 );
   and U17191 ( n17318,n16027,n17451 );
   nand U17192 ( n17451,n15982,n16028,n16012 );
   not U17193 ( n16028,n16103 );
   nor U17194 ( n16103,n14819,n17381 );
   nand U17195 ( n16027,n17381,n14819 );
   and U17196 ( n17316,n16289,n16052,n16105 );
   nand U17197 ( n16105,n16126,n14794 );
   not U17198 ( n16052,n16091 );
   nor U17199 ( n16091,n14524,n14804 );
   not U17200 ( n14804,n16064 );
   nand U17201 ( n16289,n14793,n14782 );
   and U17202 ( n17414,n17452,n15102,n17453 );
   nand U17203 ( n17453,n16340,n17305 );
   nor U17204 ( n16340,n14509,n16216 );
   nand U17205 ( n15102,n14745,n14734 );
   nand U17206 ( n17452,n17416,n17454 );
   nand U17207 ( n17454,n16246,n16282 );
   nand U17208 ( n16282,n17380,n14771 );
   nand U17209 ( n16246,n16234,n14759 );
   and U17210 ( n17416,n17305,n16189,n16338 );
   nand U17211 ( n16338,n16216,n14509 );
   nand U17212 ( n16189,n16172,n14512 );
   not U17213 ( n17305,n15104 );
   nor U17214 ( n15104,n14734,n14745 );
   not U17215 ( n14745,n14506 );
   nand U17216 ( n17297,n16422,n14697 );
   nand U17217 ( n14697,n17455,n17456 );
   nand U17218 ( n17456,n17402,n11415 );
   not U17219 ( n11415,n13563 );
   nand U17220 ( n13563,n17457,n17458,n17459,n17460 );
   nand U17221 ( n17460,n17403,n17406,n17461 );
   or U17222 ( n17459,n17403,n17462,n17461 );
   nand U17223 ( n17403,n17412,n17463 );
   nand U17224 ( n17463,n17411,n17413 );
   nand U17225 ( n17413,n17464,n17465,n17466 );
   not U17226 ( n17466,si_29_ );
   nand U17227 ( n17465,n11414,p1_datao_reg_29_ );
   nand U17228 ( n17464,n11416,p2_datao_reg_29_ );
   and U17229 ( n17411,n17467,n17468 );
   nand U17230 ( n17468,n17469,n17470 );
   not U17231 ( n17470,si_28_ );
   or U17232 ( n17469,n17471,n17472 );
   nand U17233 ( n17467,n17472,n17471 );
   nand U17234 ( n17412,n17473,n17474,si_29_ );
   or U17235 ( n17474,n11414,p2_datao_reg_29_ );
   nand U17236 ( n17473,n11414,n13540 );
   not U17237 ( n13540,p1_datao_reg_29_ );
   or U17238 ( n17458,n17406,n17461 );
   or U17239 ( n17406,n17475,si_30_ );
   nand U17240 ( n17457,n17462,n17461 );
   xor U17241 ( n17461,si_31_,n17476 );
   nand U17242 ( n17476,n17477,n17478 );
   nand U17243 ( n17478,n11414,p1_datao_reg_31_ );
   nand U17244 ( n17477,n11416,p2_datao_reg_31_ );
   not U17245 ( n17462,n17405 );
   nand U17246 ( n17405,si_30_,n17475 );
   nand U17247 ( n17475,n17479,n17480 );
   nand U17248 ( n17480,n11414,p1_datao_reg_30_ );
   nand U17249 ( n17479,n11416,p2_datao_reg_30_ );
   nand U17250 ( n17455,n17407,p2_datao_reg_31_ );
   not U17251 ( n16422,n14497 );
   nand U17252 ( n14497,n17481,n17482,n17483 );
   nand U17253 ( n17483,p1_reg2_reg_31_,n17397 );
   nand U17254 ( n17482,p1_reg0_reg_31_,n17398 );
   nand U17255 ( n17481,p1_reg1_reg_31_,n17399 );
   nand U17256 ( n16968,p1_b_reg,n17484 );
   nand U17257 ( n17484,n17485,n17486,p1_state_reg );
   nand U17258 ( n17486,n16967,n17487 );
   nand U17259 ( n17487,n16979,n17488,n16426,n17489 );
   nor U17260 ( n17489,n16915,n16960 );
   not U17261 ( n16915,n16913 );
   nand U17262 ( n17485,n16979,n16963 );
   nor U17263 ( n17493,n17494,n17495,n17496 );
   nor U17264 ( n17496,n15901,n17497 );
   not U17265 ( n15901,n14542 );
   nor U17266 ( n17495,n17498,n15823 );
   not U17267 ( n15823,n17499 );
   and U17268 ( n17494,p1_u3084,p1_reg3_reg_15_ );
   nand U17269 ( n17492,n17500,n15835 );
   xor U17270 ( n17501,n17503,n17504 );
   xor U17271 ( n17504,n17505,n17506 );
   nand U17272 ( n17490,n17507,n14548 );
   nor U17273 ( n17511,n17512,n17513,n17514 );
   nor U17274 ( n17514,n14758,n17497 );
   nor U17275 ( n17513,n17380,n17515 );
   nor U17276 ( n17512,p1_state_reg,n17516 );
   nand U17277 ( n17510,n17500,n14759 );
   nand U17278 ( n17509,n17517,n17518 );
   xor U17279 ( n17518,n17519,n17520 );
   nand U17280 ( n17520,n17521,n17522 );
   nand U17281 ( n17519,n17523,n17524 );
   nand U17282 ( n17508,n17525,n17526 );
   nor U17283 ( n17530,n16786,n17531,n17532 );
   nor U17284 ( n17532,n15456,n17515 );
   nor U17285 ( n17531,n14989,n17497 );
   nor U17286 ( n16786,p1_state_reg,n17533 );
   nand U17287 ( n17529,n17534,n17535 );
   nand U17288 ( n17528,n17536,n17517 );
   xor U17289 ( n17536,n17537,n17538 );
   xor U17290 ( n17537,n17539,n17540 );
   nand U17291 ( n17527,n17500,n14990 );
   nor U17292 ( n17544,n17545,n17546,n17547 );
   nor U17293 ( n17547,n15976,n17497 );
   nor U17294 ( n17546,n17383,n17515 );
   nor U17295 ( n17545,p1_state_reg,n17548 );
   nand U17296 ( n17543,n17549,n17535 );
   or U17297 ( n17542,n17550,n17502 );
   xor U17298 ( n17550,n17551,n17552 );
   xor U17299 ( n17551,n17553,n17554 );
   nand U17300 ( n17541,n17500,n15936 );
   nor U17301 ( n17558,n17559,n17560 );
   nor U17302 ( n17560,n15356,n17515 );
   not U17303 ( n15356,n14587 );
   nor U17304 ( n17559,n16401,n17497 );
   nand U17305 ( n17557,n17500,n15036 );
   or U17306 ( n17556,n17561,n17502 );
   xor U17307 ( n17561,n17562,n17563 );
   xor U17308 ( n17562,n17564,n17565 );
   nand U17309 ( n17555,p1_reg3_reg_2_,n17566 );
   nor U17310 ( n17570,n17571,n17572,n17573 );
   nor U17311 ( n17573,n17498,n15699 );
   not U17312 ( n15699,n17574 );
   nor U17313 ( n17572,n15698,n17575 );
   not U17314 ( n15698,n14932 );
   and U17315 ( n17571,p1_u3084,p1_reg3_reg_11_ );
   nand U17316 ( n17569,n17576,n14554 );
   xor U17317 ( n17577,n17578,n17579 );
   xor U17318 ( n17579,n17580,n17581 );
   nand U17319 ( n17567,n17507,n14560 );
   nor U17320 ( n17585,n17586,n17587,n17588 );
   nor U17321 ( n17588,n16126,n17497 );
   not U17322 ( n16126,n14521 );
   nor U17323 ( n17587,n17381,n17515 );
   nor U17324 ( n17586,p1_state_reg,n17589 );
   nand U17325 ( n17584,n17500,n16064 );
   or U17326 ( n17583,n17590,n17502 );
   xor U17327 ( n17590,n17591,n17592 );
   xor U17328 ( n17591,n17593,n17594 );
   nand U17329 ( n17582,n17595,n17526 );
   nor U17330 ( n17599,n16609,n17600,n17601 );
   nor U17331 ( n17601,n17498,n15763 );
   not U17332 ( n15763,n17602 );
   nor U17333 ( n17600,n15762,n17575 );
   not U17334 ( n15762,n14909 );
   nor U17335 ( n16609,p1_state_reg,n17603 );
   nand U17336 ( n17598,n17507,n14554 );
   nand U17337 ( n17605,n17606,n17607 );
   nand U17338 ( n17607,n17608,n17609 );
   nand U17339 ( n17604,n17608,n17609,n17610 );
   nand U17340 ( n17596,n17576,n14548 );
   nor U17341 ( n17614,n17615,n17616,n17617 );
   nor U17342 ( n17617,n17381,n17497 );
   not U17343 ( n17381,n14527 );
   nor U17344 ( n17616,n15976,n17515 );
   not U17345 ( n15976,n14533 );
   nor U17346 ( n17615,p1_state_reg,n17618 );
   nand U17347 ( n17613,n17500,n15982 );
   nand U17348 ( n17612,n17517,n17619 );
   xor U17349 ( n17619,n17620,n17621 );
   xor U17350 ( n17620,n17622,n17623 );
   nand U17351 ( n17611,n17624,n17526 );
   nand U17352 ( n17628,p1_reg3_reg_0_,n17566 );
   nand U17353 ( n17627,n17517,n16916 );
   xor U17354 ( n16916,n17629,n17630 );
   xor U17355 ( n17630,n17631,n17632 );
   not U17356 ( n17629,n17633 );
   nand U17357 ( n17626,n17500,n15056 );
   nand U17358 ( n17625,n17576,n14587 );
   nor U17359 ( n17637,n16704,n17638,n17639 );
   nor U17360 ( n17639,n14977,n17515 );
   nor U17361 ( n17638,n15707,n17497 );
   not U17362 ( n15707,n14560 );
   nor U17363 ( n16704,p1_state_reg,n17640 );
   nand U17364 ( n17636,n15636,n17535 );
   nand U17365 ( n17635,n17641,n17517 );
   xor U17366 ( n17641,n17642,n17643 );
   xor U17367 ( n17642,n17644,n17645 );
   nand U17368 ( n17634,n17500,n15646 );
   nor U17369 ( n17649,n17650,n17651,n17652 );
   nor U17370 ( n17652,n16401,n17515 );
   not U17371 ( n16401,n14581 );
   nor U17372 ( n17651,n15456,n17497 );
   not U17373 ( n15456,n14575 );
   nor U17374 ( n17650,p1_state_reg,n17653 );
   nand U17375 ( n17648,n17500,n15468 );
   nand U17376 ( n17647,n15470,n17535 );
   xor U17377 ( n17654,n17655,n17656 );
   xor U17378 ( n17655,n17657,n17658 );
   nor U17379 ( n17662,n17663,n17664,n17665 );
   nor U17380 ( n17665,n17380,n17497 );
   not U17381 ( n17380,n14515 );
   nor U17382 ( n17664,n16116,n17575 );
   not U17383 ( n16116,n14782 );
   nor U17384 ( n17663,p1_state_reg,n17666 );
   nand U17385 ( n17661,n17507,n14521 );
   nand U17386 ( n17660,n17517,n17667 );
   xor U17387 ( n17667,n17668,n17669 );
   nand U17388 ( n17668,n17670,n17671 );
   nand U17389 ( n17659,n16117,n17526 );
   nor U17390 ( n17675,n16505,n17676,n17677 );
   nor U17391 ( n17677,n17498,n15891 );
   not U17392 ( n15891,n17678 );
   nor U17393 ( n17676,n15890,n17575 );
   not U17394 ( n15890,n14864 );
   nor U17395 ( n16505,p1_state_reg,n17679 );
   nand U17396 ( n17674,n17507,n14542 );
   nand U17397 ( n17681,n17682,n17683 );
   nand U17398 ( n17683,n17684,n17685 );
   nand U17399 ( n17680,n17684,n17685,n17686 );
   nand U17400 ( n17672,n17576,n14536 );
   nor U17401 ( n17690,n16816,n17691,n17692 );
   nor U17402 ( n17692,n17372,n17515 );
   not U17403 ( n17372,n14578 );
   nor U17404 ( n17691,n15001,n17497 );
   nor U17405 ( n16816,p1_state_reg,n17693 );
   nand U17406 ( n17689,n15482,n17535 );
   nand U17407 ( n17688,n17694,n17517 );
   xor U17408 ( n17694,n17695,n17696 );
   xor U17409 ( n17695,n17697,n17698 );
   nand U17410 ( n17687,n17500,n15002 );
   nor U17411 ( n17702,n17703,n17704,n17705 );
   nor U17412 ( n17705,n17383,n17497 );
   not U17413 ( n17383,n14539 );
   nor U17414 ( n17704,n17498,n15847 );
   nor U17415 ( n17703,p1_state_reg,n17706 );
   nand U17416 ( n17701,n17500,n14875 );
   xor U17417 ( n17707,n17708,n17709 );
   xor U17418 ( n17709,n17710,n17711 );
   nand U17419 ( n17699,n17507,n14545 );
   nor U17420 ( n17715,n17716,n17717,n17718 );
   nor U17421 ( n17718,n16234,n17497 );
   nor U17422 ( n17717,n16146,n17575 );
   not U17423 ( n16146,n14771 );
   and U17424 ( n17716,p1_u3084,p1_reg3_reg_25_ );
   nand U17425 ( n17714,n17507,n14518 );
   nand U17426 ( n17713,n17517,n17719 );
   nand U17427 ( n17719,n17720,n17721 );
   nand U17428 ( n17721,n17722,n17524 );
   not U17429 ( n17722,n17523 );
   nand U17430 ( n17720,n17723,n17724 );
   nand U17431 ( n17724,n17725,n17670 );
   not U17432 ( n17723,n17726 );
   xor U17433 ( n17726,n17727,n17728 );
   nand U17434 ( n17712,n16147,n17526 );
   nor U17435 ( n17732,n16630,n17733,n17734 );
   nor U17436 ( n17734,n17382,n17497 );
   nor U17437 ( n17733,n16379,n17515 );
   nor U17438 ( n16630,p1_state_reg,n17735 );
   nand U17439 ( n17731,n17736,n17535 );
   nand U17440 ( n17730,n17517,n17737 );
   xor U17441 ( n17737,n17738,n17739 );
   xor U17442 ( n17738,n17740,n17741 );
   nand U17443 ( n17729,n17500,n15753 );
   nor U17444 ( n17745,n17746,n17747,n17748 );
   nor U17445 ( n17748,n16001,n17575 );
   not U17446 ( n16001,n14819 );
   nor U17447 ( n17747,n16012,n17515 );
   not U17448 ( n16012,n14530 );
   nor U17449 ( n17746,p1_state_reg,n17749 );
   nand U17450 ( n17744,n17576,n14524 );
   nand U17451 ( n17743,n17750,n17751,n17517 );
   nand U17452 ( n17751,n17752,n17753 );
   nand U17453 ( n17753,n17754,n17755 );
   nand U17454 ( n17750,n17754,n17755,n17756 );
   nand U17455 ( n17742,n16002,n17526 );
   nand U17456 ( n17760,n17500,n15385 );
   nor U17457 ( n17759,n17761,n17762 );
   and U17458 ( n17762,n17566,p1_reg3_reg_1_ );
   nand U17459 ( n17566,n17498,p1_state_reg );
   nor U17460 ( n17761,n17502,n17763 );
   xor U17461 ( n17763,n17764,n17765 );
   xor U17462 ( n17764,n17766,n17767 );
   nand U17463 ( n17758,n17576,n14584 );
   nand U17464 ( n17757,n17507,n14590 );
   nor U17465 ( n17771,n16731,n17772,n17773 );
   nor U17466 ( n17773,n14989,n17515 );
   not U17467 ( n14989,n14569 );
   nor U17468 ( n17772,n17498,n15599 );
   nor U17469 ( n16731,p1_state_reg,n17774 );
   nand U17470 ( n17770,n17576,n14563 );
   or U17471 ( n17769,n17775,n17502 );
   xor U17472 ( n17775,n17776,n17777 );
   xor U17473 ( n17776,n17778,n17779 );
   nand U17474 ( n17768,n17500,n14966 );
   nor U17475 ( n17783,n17784,n17785,n17786 );
   nor U17476 ( n17786,n14758,n17515 );
   not U17477 ( n14758,n14509 );
   and U17478 ( n17785,n17526,n16263 );
   nor U17479 ( n17784,p1_state_reg,n17787 );
   nand U17480 ( n17782,n17500,n14734 );
   nand U17481 ( n17789,n17790,n17791 );
   nand U17482 ( n17791,n17792,n17793 );
   or U17483 ( n17793,n17794,n17795 );
   not U17484 ( n17790,n17796 );
   nand U17485 ( n17788,n17796,n17797 );
   nand U17486 ( n17797,n17798,n17799 );
   nand U17487 ( n17799,n17794,n17792 );
   not U17488 ( n17792,n17800 );
   xor U17489 ( n17796,n17801,n17802 );
   nand U17490 ( n17802,n17803,n17804 );
   nand U17491 ( n17804,n17805,n14734 );
   nand U17492 ( n17803,n17806,n14506 );
   nand U17493 ( n17807,n17809,n17810 );
   nand U17494 ( n17810,n17811,n14734 );
   nand U17495 ( n14734,n17812,n17813 );
   nand U17496 ( n17813,n17402,n11390 );
   xor U17497 ( n11390,n17472,n17814 );
   xor U17498 ( n17814,si_28_,n17471 );
   nand U17499 ( n17471,n17815,n17816 );
   nand U17500 ( n17816,n17817,n17818 );
   not U17501 ( n17818,si_27_ );
   or U17502 ( n17817,n17819,n17820 );
   nand U17503 ( n17815,n17820,n17819 );
   nand U17504 ( n17472,n17821,n17822 );
   or U17505 ( n17822,n11414,p2_datao_reg_28_ );
   nand U17506 ( n17821,n11414,n13901 );
   not U17507 ( n13901,p1_datao_reg_28_ );
   nand U17508 ( n17812,n17407,p2_datao_reg_28_ );
   nand U17509 ( n17809,n17805,n14506 );
   nand U17510 ( n17780,n17576,n14503 );
   nand U17511 ( n14503,n17823,n17824,n17825,n17826 );
   nand U17512 ( n17826,n17827,n15085 );
   nor U17513 ( n15085,n17828,n17829,n17787 );
   not U17514 ( n17787,p1_reg3_reg_28_ );
   nand U17515 ( n17825,p1_reg0_reg_29_,n17398 );
   nand U17516 ( n17824,p1_reg1_reg_29_,n17399 );
   nand U17517 ( n17823,p1_reg2_reg_29_,n17397 );
   nor U17518 ( n17833,n16440,n17834,n17835 );
   nor U17519 ( n17835,n17498,n15945 );
   not U17520 ( n15945,n17836 );
   nor U17521 ( n17834,n14839,n17575 );
   not U17522 ( n14839,n15953 );
   nor U17523 ( n16440,p1_state_reg,n17837 );
   nand U17524 ( n17832,n17576,n14530 );
   xor U17525 ( n17838,n17839,n17840 );
   xor U17526 ( n17840,n17841,n17842 );
   nand U17527 ( n17830,n17507,n14536 );
   nor U17528 ( n17846,n17847,n16877,n17848 );
   nor U17529 ( n17848,p1_reg3_reg_3_,n17498 );
   nor U17530 ( n16877,p1_state_reg,n17849 );
   nor U17531 ( n17847,n17373,n17515 );
   not U17532 ( n17373,n14584 );
   nand U17533 ( n17845,n17576,n14578 );
   nand U17534 ( n17844,n17850,n17851,n17517 );
   nand U17535 ( n17851,n17852,n17853 );
   nand U17536 ( n17853,n17854,n17855 );
   nand U17537 ( n17850,n17854,n17855,n17856 );
   nand U17538 ( n17843,n17500,n15443 );
   nor U17539 ( n17860,n16683,n17861,n17862 );
   nor U17540 ( n17862,n16379,n17497 );
   not U17541 ( n16379,n14557 );
   nor U17542 ( n17861,n17498,n15656 );
   not U17543 ( n15656,n17863 );
   not U17544 ( n17498,n17535 );
   nor U17545 ( n16683,p1_state_reg,n17864 );
   nand U17546 ( n17859,n17500,n15678 );
   xor U17547 ( n17865,n17866,n17867 );
   xor U17548 ( n17867,n17868,n17869 );
   nand U17549 ( n17857,n17507,n14563 );
   nor U17550 ( n17873,n17874,n17875,n17876 );
   nor U17551 ( n17876,n14793,n17497 );
   not U17552 ( n14793,n14518 );
   nor U17553 ( n17875,n16073,n17575 );
   not U17554 ( n16073,n14794 );
   nor U17555 ( n17874,p1_state_reg,n17877 );
   nand U17556 ( n17872,n17507,n14524 );
   or U17557 ( n17871,n17878,n17502 );
   xor U17558 ( n17878,n17879,n17880 );
   xor U17559 ( n17880,n17881,n17882 );
   nand U17560 ( n17870,n16074,n17526 );
   nor U17561 ( n17886,n17887,n17888,n17889 );
   nor U17562 ( n17889,n15874,n17497 );
   not U17563 ( n15874,n14545 );
   nor U17564 ( n17888,n17382,n17515 );
   not U17565 ( n17382,n14551 );
   nor U17566 ( n17887,p1_state_reg,n17890 );
   nand U17567 ( n17885,n15798,n17535 );
   or U17568 ( n17884,n17891,n17502 );
   xor U17569 ( n17891,n17892,n17893 );
   xor U17570 ( n17892,n17894,n17895 );
   nand U17571 ( n17883,n17500,n15814 );
   nor U17572 ( n17899,n17900,n17901,n17902 );
   nor U17573 ( n17902,n16234,n17515 );
   not U17574 ( n16234,n14512 );
   nor U17575 ( n17901,n16216,n17575 );
   not U17576 ( n16216,n14746 );
   nor U17577 ( n17900,p1_state_reg,n17828 );
   nand U17578 ( n17898,n17576,n14506 );
   nand U17579 ( n14506,n17903,n17904,n17905,n17906 );
   nand U17580 ( n17906,n17827,n16263 );
   xor U17581 ( n16263,n17907,p1_reg3_reg_28_ );
   nor U17582 ( n17907,n17829,n17828 );
   nand U17583 ( n17905,p1_reg0_reg_28_,n17398 );
   nand U17584 ( n17904,p1_reg1_reg_28_,n17399 );
   nand U17585 ( n17903,p1_reg2_reg_28_,n17397 );
   nand U17586 ( n17897,n17908,n17517 );
   xor U17587 ( n17908,n17909,n17794 );
   nand U17588 ( n17794,n17522,n17910 );
   nand U17589 ( n17910,n17521,n17524,n17523 );
   nand U17590 ( n17523,n17725,n17670,n17911 );
   nand U17591 ( n17911,n17727,n17728 );
   nand U17592 ( n17670,n17912,n17913 );
   nand U17593 ( n17725,n17915,n17671 );
   nand U17594 ( n17671,n17916,n17917 );
   not U17595 ( n17917,n17913 );
   nand U17596 ( n17913,n17918,n17919 );
   nand U17597 ( n17919,n17805,n14782 );
   nand U17598 ( n17918,n17806,n14518 );
   xor U17599 ( n17916,n17631,n17914 );
   nand U17600 ( n17914,n17920,n17921 );
   nand U17601 ( n17921,n17811,n14782 );
   nand U17602 ( n14782,n17922,n17923 );
   nand U17603 ( n17923,n17402,n11354 );
   xor U17604 ( n11354,n17924,n17925 );
   xor U17605 ( n17925,si_24_,n17926 );
   nand U17606 ( n17922,n17407,p2_datao_reg_24_ );
   nand U17607 ( n17920,n17805,n14518 );
   nand U17608 ( n14518,n17927,n17928,n17929,n17930 );
   nand U17609 ( n17930,n16117,n17827 );
   nor U17610 ( n16117,n17931,n17932 );
   and U17611 ( n17931,n17666,n17933 );
   nand U17612 ( n17933,p1_reg3_reg_23_,n17934 );
   nand U17613 ( n17929,p1_reg0_reg_24_,n17398 );
   nand U17614 ( n17928,p1_reg1_reg_24_,n17399 );
   nand U17615 ( n17927,p1_reg2_reg_24_,n17397 );
   not U17616 ( n17915,n17669 );
   nand U17617 ( n17669,n17935,n17936 );
   nand U17618 ( n17936,n17879,n17937 );
   or U17619 ( n17937,n17882,n17881 );
   xor U17620 ( n17879,n17631,n17938 );
   nand U17621 ( n17938,n17939,n17940 );
   nand U17622 ( n17940,n17811,n14794 );
   nand U17623 ( n17939,n17805,n14521 );
   nand U17624 ( n17935,n17881,n17882 );
   nand U17625 ( n17882,n17941,n17942 );
   nand U17626 ( n17942,n17943,n17594 );
   nand U17627 ( n17594,n17944,n17755 );
   nand U17628 ( n17755,n17945,n17946 );
   not U17629 ( n17946,n17947 );
   xor U17630 ( n17945,n17631,n17948 );
   nand U17631 ( n17944,n17752,n17754 );
   nand U17632 ( n17754,n17949,n17947 );
   nand U17633 ( n17947,n17950,n17951 );
   nand U17634 ( n17951,n17805,n14819 );
   nand U17635 ( n17950,n17806,n14527 );
   nand U17636 ( n17948,n17952,n17953 );
   nand U17637 ( n17953,n17811,n14819 );
   nand U17638 ( n14819,n17954,n17955 );
   nand U17639 ( n17955,n17402,n11328 );
   xor U17640 ( n11328,n17956,n17957 );
   xor U17641 ( n17957,si_21_,n17958 );
   nand U17642 ( n17954,n17407,p2_datao_reg_21_ );
   nand U17643 ( n17952,n17805,n14527 );
   nand U17644 ( n14527,n17959,n17960,n17961,n17962 );
   nand U17645 ( n17962,n17827,n16002 );
   xor U17646 ( n16002,p1_reg3_reg_21_,n17963 );
   nand U17647 ( n17961,p1_reg0_reg_21_,n17398 );
   nand U17648 ( n17960,p1_reg1_reg_21_,n17399 );
   nand U17649 ( n17959,p1_reg2_reg_21_,n17397 );
   not U17650 ( n17752,n17756 );
   nand U17651 ( n17756,n17964,n17965 );
   nand U17652 ( n17965,n17966,n17623 );
   nand U17653 ( n17623,n17967,n17968 );
   nand U17654 ( n17968,n17805,n15982 );
   nand U17655 ( n17967,n17806,n14530 );
   nand U17656 ( n17966,n17622,n17621 );
   or U17657 ( n17964,n17621,n17622 );
   and U17658 ( n17622,n17969,n17970 );
   nand U17659 ( n17970,n17842,n17971 );
   or U17660 ( n17971,n17841,n17839 );
   and U17661 ( n17842,n17972,n17973 );
   nand U17662 ( n17973,n17974,n17554 );
   nand U17663 ( n17554,n17975,n17685 );
   nand U17664 ( n17685,n17976,n17977 );
   not U17665 ( n17977,n17978 );
   xor U17666 ( n17976,n17631,n17979 );
   nand U17667 ( n17975,n17682,n17684 );
   nand U17668 ( n17684,n17980,n17978 );
   nand U17669 ( n17978,n17981,n17982 );
   nand U17670 ( n17982,n17805,n14864 );
   nand U17671 ( n17981,n17806,n14539 );
   nand U17672 ( n17979,n17983,n17984 );
   nand U17673 ( n17984,n17811,n14864 );
   nand U17674 ( n14864,n17985,n17986,n17987 );
   nand U17675 ( n17987,n17407,p2_datao_reg_17_ );
   nand U17676 ( n17986,n16508,n16427 );
   not U17677 ( n16508,n16490 );
   nand U17678 ( n16490,n17988,n17989,n15248 );
   nand U17679 ( n17989,n15240,n17990 );
   not U17680 ( n15240,p1_ir_reg_17_ );
   nand U17681 ( n17988,p1_ir_reg_17_,n15232,p1_ir_reg_31_ );
   nand U17682 ( n17985,n17402,n11295 );
   not U17683 ( n11295,n14058 );
   xor U17684 ( n14058,n17991,n17992 );
   xor U17685 ( n17991,n17993,n17994 );
   nand U17686 ( n17983,n17805,n14539 );
   nand U17687 ( n14539,n17995,n17996,n17997,n17998 );
   nand U17688 ( n17998,n17827,n17678 );
   xor U17689 ( n17678,n17679,n17999 );
   nand U17690 ( n17997,p1_reg0_reg_17_,n17398 );
   nand U17691 ( n17996,p1_reg1_reg_17_,n17399 );
   nand U17692 ( n17995,p1_reg2_reg_17_,n17397 );
   not U17693 ( n17682,n17686 );
   nand U17694 ( n17686,n18000,n18001 );
   nand U17695 ( n18001,n17708,n18002 );
   nand U17696 ( n18002,n17710,n17711 );
   xor U17697 ( n17708,n17808,n18003 );
   nand U17698 ( n18003,n18004,n18005 );
   nand U17699 ( n18005,n17811,n14875 );
   nand U17700 ( n18004,n17805,n14542 );
   or U17701 ( n18000,n17711,n17710 );
   and U17702 ( n17710,n18006,n18007 );
   nand U17703 ( n18007,n17805,n14875 );
   nand U17704 ( n14875,n18008,n18009,n18010 );
   nand U17705 ( n18010,n17407,p2_datao_reg_16_ );
   nand U17706 ( n18009,n16518,n16427 );
   not U17707 ( n16518,n16519 );
   nand U17708 ( n16519,n18011,n18012 );
   or U17709 ( n18012,p1_ir_reg_16_,p1_ir_reg_31_ );
   nand U17710 ( n18011,p1_ir_reg_31_,n18013 );
   nand U17711 ( n18013,n15231,n15232 );
   nand U17712 ( n15231,p1_ir_reg_16_,n18014 );
   nand U17713 ( n18008,n17402,n11285 );
   not U17714 ( n11285,n14202 );
   xor U17715 ( n14202,n18015,n18016 );
   xor U17716 ( n18015,n18017,n18018 );
   nand U17717 ( n18006,n17806,n14542 );
   nand U17718 ( n14542,n18019,n18020,n18021,n18022 );
   nand U17719 ( n18022,n18023,n17827 );
   not U17720 ( n18023,n15847 );
   nand U17721 ( n15847,n18024,n17999 );
   nand U17722 ( n18024,n17706,n18025 );
   nand U17723 ( n18025,p1_reg3_reg_15_,n18026 );
   not U17724 ( n17706,p1_reg3_reg_16_ );
   nand U17725 ( n18021,p1_reg0_reg_16_,n17398 );
   nand U17726 ( n18020,p1_reg1_reg_16_,n17399 );
   nand U17727 ( n18019,p1_reg2_reg_16_,n17397 );
   nand U17728 ( n17711,n18027,n18028 );
   nand U17729 ( n18028,n17503,n18029 );
   nand U17730 ( n18029,n17506,n17505 );
   xor U17731 ( n17503,n17631,n18030 );
   nand U17732 ( n18030,n18031,n18032 );
   nand U17733 ( n18032,n17811,n15835 );
   nand U17734 ( n18031,n17805,n14545 );
   or U17735 ( n18027,n17505,n17506 );
   and U17736 ( n17506,n18033,n18034 );
   nand U17737 ( n18034,n18035,n17895 );
   nand U17738 ( n17895,n18036,n17609 );
   nand U17739 ( n17609,n18037,n18038 );
   not U17740 ( n18038,n18039 );
   xor U17741 ( n18037,n17631,n18040 );
   nand U17742 ( n18036,n17606,n17608 );
   nand U17743 ( n17608,n18041,n18039 );
   nand U17744 ( n18039,n18042,n18043 );
   nand U17745 ( n18043,n17805,n14909 );
   nand U17746 ( n18042,n17806,n14551 );
   nand U17747 ( n18040,n18044,n18045 );
   nand U17748 ( n18045,n17811,n14909 );
   nand U17749 ( n14909,n18046,n18047,n18048 );
   nand U17750 ( n18048,n17407,p2_datao_reg_13_ );
   nand U17751 ( n18047,n16611,n16427 );
   not U17752 ( n16611,n16618 );
   nand U17753 ( n16618,n18049,n18050,n18051 );
   nand U17754 ( n18050,n15211,n17990 );
   nand U17755 ( n18049,p1_ir_reg_13_,n15203,p1_ir_reg_31_ );
   nand U17756 ( n18046,n17402,n11261 );
   nand U17757 ( n11261,n18052,n18053 );
   nand U17758 ( n18053,n18054,n18055 );
   nand U17759 ( n18054,n18056,n18057 );
   nand U17760 ( n18052,n18058,n18059 );
   xor U17761 ( n18059,si_13_,n18060 );
   not U17762 ( n18058,n18055 );
   nand U17763 ( n18055,n18061,n18062 );
   nand U17764 ( n18062,n18063,n18064 );
   nand U17765 ( n18044,n17805,n14551 );
   nand U17766 ( n14551,n18065,n18066,n18067,n18068 );
   nand U17767 ( n18068,n17827,n17602 );
   xor U17768 ( n17602,n17603,n18069 );
   nand U17769 ( n18067,p1_reg0_reg_13_,n17398 );
   nand U17770 ( n18066,p1_reg1_reg_13_,n17399 );
   nand U17771 ( n18065,p1_reg2_reg_13_,n17397 );
   not U17772 ( n17606,n17610 );
   nand U17773 ( n17610,n18070,n18071 );
   nand U17774 ( n18071,n18072,n17741 );
   nand U17775 ( n17741,n18073,n18074 );
   nand U17776 ( n18074,n17805,n15753 );
   nand U17777 ( n18073,n17806,n14554 );
   nand U17778 ( n18072,n17740,n17739 );
   or U17779 ( n18070,n17739,n17740 );
   and U17780 ( n17740,n18075,n18076 );
   nand U17781 ( n18076,n17581,n18077 );
   or U17782 ( n18077,n17580,n17578 );
   and U17783 ( n17581,n18078,n18079 );
   nand U17784 ( n18079,n17866,n18080 );
   or U17785 ( n18080,n17869,n17868 );
   xor U17786 ( n17866,n17631,n18081 );
   nand U17787 ( n18081,n18082,n18083 );
   nand U17788 ( n18083,n17811,n15678 );
   nand U17789 ( n18082,n17805,n14560 );
   nand U17790 ( n18078,n17868,n17869 );
   nand U17791 ( n17869,n18084,n18085 );
   nand U17792 ( n18085,n18086,n18087 );
   or U17793 ( n18087,n17644,n17643 );
   not U17794 ( n18086,n17645 );
   nand U17795 ( n17645,n18088,n18089 );
   nand U17796 ( n18089,n17806,n14563 );
   nand U17797 ( n18088,n17805,n15646 );
   nand U17798 ( n18084,n17643,n17644 );
   nand U17799 ( n17644,n18090,n18091 );
   nand U17800 ( n18091,n18092,n17778 );
   nand U17801 ( n17778,n18093,n18094 );
   nand U17802 ( n18093,n18095,n18096 );
   nand U17803 ( n18092,n17777,n17779 );
   or U17804 ( n18090,n17779,n17777 );
   xor U17805 ( n17777,n17808,n18097 );
   nand U17806 ( n18097,n18098,n18099 );
   nand U17807 ( n18099,n17811,n14966 );
   nand U17808 ( n18098,n17805,n14566 );
   nand U17809 ( n17779,n18100,n18101 );
   nand U17810 ( n18101,n17805,n14966 );
   nand U17811 ( n14966,n18102,n18103,n18104 );
   nand U17812 ( n18104,n17407,p2_datao_reg_8_ );
   nand U17813 ( n18103,n16733,n16427 );
   not U17814 ( n16733,n16751 );
   nand U17815 ( n16751,n18105,n18106 );
   or U17816 ( n18106,p1_ir_reg_31_,p1_ir_reg_8_ );
   nand U17817 ( n18105,p1_ir_reg_31_,n18107 );
   nand U17818 ( n18107,n15180,n15181 );
   nand U17819 ( n15180,p1_ir_reg_8_,n18108 );
   nand U17820 ( n18102,n17402,n11218 );
   xor U17821 ( n11218,n18109,n18110 );
   and U17822 ( n18109,n18111,n18112 );
   nand U17823 ( n18100,n17806,n14566 );
   xor U17824 ( n17643,n17631,n18113 );
   nand U17825 ( n18113,n18114,n18115 );
   nand U17826 ( n18115,n17811,n15646 );
   nand U17827 ( n15646,n18116,n18117,n18118 );
   nand U17828 ( n18118,n17407,p2_datao_reg_9_ );
   nand U17829 ( n18117,n16706,n16427 );
   and U17830 ( n16706,n18119,n18120 );
   nand U17831 ( n18120,n17990,n18121 );
   or U17832 ( n18119,n15186,n17990 );
   xor U17833 ( n15186,n18121,n18122 );
   nand U17834 ( n18116,n17402,n11227 );
   xor U17835 ( n11227,n18123,n18124 );
   and U17836 ( n18123,n18125,n18126 );
   nand U17837 ( n18114,n17805,n14563 );
   nand U17838 ( n14563,n18127,n18128,n18129,n18130 );
   nand U17839 ( n18130,n17827,n15636 );
   xor U17840 ( n15636,p1_reg3_reg_9_,n18131 );
   nand U17841 ( n18129,p1_reg0_reg_9_,n17398 );
   nand U17842 ( n18128,p1_reg1_reg_9_,n17399 );
   nand U17843 ( n18127,p1_reg2_reg_9_,n17397 );
   and U17844 ( n17868,n18132,n18133 );
   nand U17845 ( n18133,n17806,n14560 );
   nand U17846 ( n14560,n18134,n18135,n18136,n18137 );
   nand U17847 ( n18137,n17863,n17827 );
   nor U17848 ( n17863,n18138,n18139 );
   and U17849 ( n18138,n17864,n18140 );
   nand U17850 ( n18140,p1_reg3_reg_9_,n18131 );
   nand U17851 ( n18136,p1_reg0_reg_10_,n17398 );
   nand U17852 ( n18135,p1_reg1_reg_10_,n17399 );
   nand U17853 ( n18134,p1_reg2_reg_10_,n17397 );
   nand U17854 ( n18132,n17805,n15678 );
   nand U17855 ( n15678,n18141,n18142,n18143 );
   nand U17856 ( n18143,n17407,p2_datao_reg_10_ );
   nand U17857 ( n18142,n16685,n16427 );
   not U17858 ( n16685,n16691 );
   nand U17859 ( n16691,n18144,n18145 );
   or U17860 ( n18145,p1_ir_reg_10_,p1_ir_reg_31_ );
   nand U17861 ( n18144,p1_ir_reg_31_,n15192 );
   nand U17862 ( n15192,n18146,n18147 );
   nand U17863 ( n18147,p1_ir_reg_10_,n18148 );
   nand U17864 ( n18148,n18122,n18121 );
   not U17865 ( n18121,p1_ir_reg_9_ );
   nand U17866 ( n18141,n17402,n11234 );
   xor U17867 ( n11234,n18149,n18150 );
   xor U17868 ( n18150,si_10_,n18151 );
   nand U17869 ( n18075,n17578,n17580 );
   nand U17870 ( n17580,n18152,n18153 );
   nand U17871 ( n18153,n17806,n14557 );
   nand U17872 ( n18152,n17805,n14932 );
   xor U17873 ( n17578,n17808,n18154 );
   nand U17874 ( n18154,n18155,n18156 );
   nand U17875 ( n18156,n17811,n14932 );
   nand U17876 ( n14932,n18157,n18158,n18159 );
   nand U17877 ( n18159,n17407,p2_datao_reg_11_ );
   nand U17878 ( n18158,n16646,n16427 );
   not U17879 ( n16646,n16644 );
   nand U17880 ( n16644,n18160,n18161 );
   nand U17881 ( n18161,n18162,n17990 );
   or U17882 ( n18160,n15197,n17990 );
   xor U17883 ( n15197,n18146,p1_ir_reg_11_ );
   nand U17884 ( n18157,n17402,n11244 );
   xor U17885 ( n11244,n18163,n18164 );
   nor U17886 ( n18163,n18165,n18166 );
   nand U17887 ( n18155,n17805,n14557 );
   nand U17888 ( n14557,n18167,n18168,n18169,n18170 );
   nand U17889 ( n18170,n17827,n17574 );
   xor U17890 ( n17574,p1_reg3_reg_11_,n18139 );
   nand U17891 ( n18169,p1_reg0_reg_11_,n17398 );
   nand U17892 ( n18168,p1_reg1_reg_11_,n17399 );
   nand U17893 ( n18167,p1_reg2_reg_11_,n17397 );
   xor U17894 ( n17739,n17631,n18171 );
   nand U17895 ( n18171,n18172,n18173 );
   nand U17896 ( n18173,n17811,n15753 );
   nand U17897 ( n15753,n18174,n18175,n18176 );
   nand U17898 ( n18176,n17407,p2_datao_reg_12_ );
   nand U17899 ( n18175,n16632,n16427 );
   not U17900 ( n16632,n16649 );
   nand U17901 ( n16649,n18177,n18178 );
   or U17902 ( n18178,p1_ir_reg_12_,p1_ir_reg_31_ );
   nand U17903 ( n18177,p1_ir_reg_31_,n18179 );
   nand U17904 ( n18179,n15202,n15203 );
   not U17905 ( n15203,n15210 );
   nand U17906 ( n15202,p1_ir_reg_12_,n18180 );
   nand U17907 ( n18180,n18181,n18162 );
   not U17908 ( n18162,p1_ir_reg_11_ );
   nand U17909 ( n18174,n17402,n11251 );
   xor U17910 ( n11251,n18182,n18063 );
   nand U17911 ( n18063,n18183,n18184 );
   nand U17912 ( n18184,n18185,n18164 );
   and U17913 ( n18182,n18061,n18064 );
   nand U17914 ( n18172,n17805,n14554 );
   nand U17915 ( n14554,n18186,n18187,n18188,n18189 );
   nand U17916 ( n18189,n17736,n17827 );
   not U17917 ( n17736,n15742 );
   nand U17918 ( n15742,n18190,n18069 );
   nand U17919 ( n18190,n17735,n18191 );
   nand U17920 ( n18191,p1_reg3_reg_11_,n18139 );
   not U17921 ( n17735,p1_reg3_reg_12_ );
   nand U17922 ( n18188,p1_reg0_reg_12_,n17398 );
   nand U17923 ( n18187,p1_reg1_reg_12_,n17399 );
   nand U17924 ( n18186,p1_reg2_reg_12_,n17397 );
   nand U17925 ( n18035,n17893,n17894 );
   or U17926 ( n18033,n17894,n17893 );
   xor U17927 ( n17893,n17808,n18192 );
   nand U17928 ( n18192,n18193,n18194 );
   nand U17929 ( n18194,n17811,n15814 );
   nand U17930 ( n18193,n17805,n14548 );
   nand U17931 ( n17894,n18195,n18196 );
   nand U17932 ( n18196,n17805,n15814 );
   nand U17933 ( n15814,n18197,n18198,n18199 );
   nand U17934 ( n18199,n17407,p2_datao_reg_14_ );
   nand U17935 ( n18198,n16588,n16427 );
   not U17936 ( n16588,n16573 );
   nand U17937 ( n16573,n18200,n18201 );
   or U17938 ( n18201,p1_ir_reg_14_,p1_ir_reg_31_ );
   nand U17939 ( n18200,p1_ir_reg_31_,n15217 );
   nand U17940 ( n15217,n15225,n18202 );
   nand U17941 ( n18202,p1_ir_reg_14_,n18051 );
   nand U17942 ( n18197,n17402,n11268 );
   xor U17943 ( n11268,n18203,n18204 );
   xor U17944 ( n18204,si_14_,n18205 );
   nand U17945 ( n18205,n18206,n18207 );
   nand U17946 ( n18195,n17806,n14548 );
   nand U17947 ( n14548,n18208,n18209,n18210,n18211 );
   nand U17948 ( n18211,n15798,n17827 );
   nor U17949 ( n15798,n18212,n18026 );
   and U17950 ( n18212,n17890,n18213 );
   or U17951 ( n18213,n17603,n18069 );
   nand U17952 ( n18210,p1_reg0_reg_14_,n17398 );
   nand U17953 ( n18209,p1_reg1_reg_14_,n17399 );
   nand U17954 ( n18208,p1_reg2_reg_14_,n17397 );
   nand U17955 ( n17505,n18214,n18215 );
   nand U17956 ( n18215,n17806,n14545 );
   nand U17957 ( n14545,n18216,n18217,n18218,n18219 );
   nand U17958 ( n18219,n17827,n17499 );
   xor U17959 ( n17499,p1_reg3_reg_15_,n18026 );
   nand U17960 ( n18218,p1_reg0_reg_15_,n17398 );
   nand U17961 ( n18217,p1_reg1_reg_15_,n17399 );
   nand U17962 ( n18216,p1_reg2_reg_15_,n17397 );
   nand U17963 ( n18214,n17805,n15835 );
   nand U17964 ( n15835,n18220,n18221,n18222 );
   nand U17965 ( n18222,n17407,p2_datao_reg_15_ );
   nand U17966 ( n18221,n16558,n16427 );
   not U17967 ( n16558,n16547 );
   nand U17968 ( n16547,n18223,n18224,n18014 );
   nand U17969 ( n18224,n15226,n17990 );
   nand U17970 ( n18223,p1_ir_reg_15_,n15225,p1_ir_reg_31_ );
   not U17971 ( n15225,n15224 );
   nand U17972 ( n18220,n17402,n11278 );
   not U17973 ( n11278,n14076 );
   xor U17974 ( n14076,n18225,n18226 );
   xor U17975 ( n18225,n18227,n18228 );
   nand U17976 ( n17974,n17552,n17553 );
   or U17977 ( n17972,n17553,n17552 );
   xor U17978 ( n17552,n17808,n18229 );
   nand U17979 ( n18229,n18230,n18231 );
   nand U17980 ( n18231,n17811,n15936 );
   nand U17981 ( n18230,n17805,n14536 );
   nand U17982 ( n17553,n18232,n18233 );
   nand U17983 ( n18233,n17805,n15936 );
   nand U17984 ( n15936,n18234,n18235,n18236 );
   nand U17985 ( n18236,n17407,p2_datao_reg_18_ );
   nand U17986 ( n18235,n16458,n16427 );
   not U17987 ( n16458,n16456 );
   nand U17988 ( n16456,n18237,n18238,n18239 );
   nand U17989 ( n18238,n15249,n17990 );
   nand U17990 ( n18237,p1_ir_reg_18_,n15248,p1_ir_reg_31_ );
   not U17991 ( n15248,n15247 );
   nand U17992 ( n18234,n17402,n11305 );
   xor U17993 ( n11305,n18240,n18241 );
   xor U17994 ( n18241,si_18_,n18242 );
   nand U17995 ( n18232,n17806,n14536 );
   nand U17996 ( n14536,n18243,n18244,n18245,n18246 );
   nand U17997 ( n18246,n17549,n17827 );
   not U17998 ( n17549,n15924 );
   nand U17999 ( n15924,n18247,n18248 );
   nand U18000 ( n18247,n17548,n18249 );
   or U18001 ( n18249,n17679,n17999 );
   nand U18002 ( n18245,p1_reg0_reg_18_,n17398 );
   nand U18003 ( n18244,p1_reg1_reg_18_,n17399 );
   nand U18004 ( n18243,p1_reg2_reg_18_,n17397 );
   nand U18005 ( n17969,n17839,n17841 );
   nand U18006 ( n17841,n18250,n18251 );
   nand U18007 ( n18251,n17806,n14533 );
   nand U18008 ( n18250,n17805,n15953 );
   xor U18009 ( n17839,n17808,n18252 );
   nand U18010 ( n18252,n18253,n18254 );
   nand U18011 ( n18254,n17811,n15953 );
   nand U18012 ( n15953,n18255,n18256,n18257 );
   nand U18013 ( n18257,n16427,n16443 );
   nand U18014 ( n18256,n17402,n11312 );
   xor U18015 ( n11312,n18258,n18259 );
   xor U18016 ( n18259,si_19_,n18260 );
   nand U18017 ( n18255,n17407,p2_datao_reg_19_ );
   nand U18018 ( n18253,n17805,n14533 );
   nand U18019 ( n14533,n18261,n18262,n18263,n18264 );
   nand U18020 ( n18264,n17827,n17836 );
   xor U18021 ( n17836,p1_reg3_reg_19_,n18265 );
   nand U18022 ( n18263,p1_reg0_reg_19_,n17398 );
   nand U18023 ( n18262,p1_reg1_reg_19_,n17399 );
   nand U18024 ( n18261,p1_reg2_reg_19_,n17397 );
   xor U18025 ( n17621,n17631,n18266 );
   nand U18026 ( n18266,n18267,n18268 );
   nand U18027 ( n18268,n17811,n15982 );
   nand U18028 ( n15982,n18269,n18270 );
   nand U18029 ( n18270,n17402,n11319 );
   xor U18030 ( n11319,n18271,n18272 );
   xor U18031 ( n18272,si_20_,n18273 );
   nand U18032 ( n18269,n17407,p2_datao_reg_20_ );
   nand U18033 ( n18267,n17805,n14530 );
   nand U18034 ( n14530,n18274,n18275,n18276,n18277 );
   nand U18035 ( n18277,n17624,n17827 );
   not U18036 ( n17624,n15963 );
   nand U18037 ( n15963,n18278,n18279 );
   nand U18038 ( n18278,n17618,n18280 );
   nand U18039 ( n18280,p1_reg3_reg_19_,n18265 );
   nand U18040 ( n18276,p1_reg0_reg_20_,n17398 );
   nand U18041 ( n18275,p1_reg1_reg_20_,n17399 );
   nand U18042 ( n18274,p1_reg2_reg_20_,n17397 );
   nand U18043 ( n17943,n17592,n17593 );
   or U18044 ( n17941,n17593,n17592 );
   xor U18045 ( n17592,n17808,n18281 );
   nand U18046 ( n18281,n18282,n18283 );
   nand U18047 ( n18283,n17811,n16064 );
   nand U18048 ( n18282,n17805,n14524 );
   nand U18049 ( n17593,n18284,n18285 );
   nand U18050 ( n18285,n17805,n16064 );
   nand U18051 ( n16064,n18286,n18287 );
   nand U18052 ( n18287,n17402,n11338 );
   xor U18053 ( n11338,n18288,n18289 );
   xor U18054 ( n18289,si_22_,n18290 );
   nand U18055 ( n18286,n17407,p2_datao_reg_22_ );
   nand U18056 ( n18284,n17806,n14524 );
   nand U18057 ( n14524,n18291,n18292,n18293,n18294 );
   nand U18058 ( n18294,n17595,n17827 );
   not U18059 ( n17595,n16046 );
   nand U18060 ( n16046,n18295,n18296 );
   nand U18061 ( n18295,n17589,n18297 );
   nand U18062 ( n18297,p1_reg3_reg_21_,n17963 );
   nand U18063 ( n18293,p1_reg0_reg_22_,n17398 );
   nand U18064 ( n18292,p1_reg1_reg_22_,n17399 );
   nand U18065 ( n18291,p1_reg2_reg_22_,n17397 );
   and U18066 ( n17881,n18298,n18299 );
   nand U18067 ( n18299,n17806,n14521 );
   nand U18068 ( n14521,n18300,n18301,n18302,n18303 );
   nand U18069 ( n18303,n17827,n16074 );
   xor U18070 ( n16074,p1_reg3_reg_23_,n17934 );
   nand U18071 ( n18302,p1_reg0_reg_23_,n17398 );
   nand U18072 ( n18301,p1_reg1_reg_23_,n17399 );
   nand U18073 ( n18300,p1_reg2_reg_23_,n17397 );
   nand U18074 ( n18298,n17805,n14794 );
   nand U18075 ( n14794,n18304,n18305 );
   nand U18076 ( n18305,n17402,n11345 );
   xor U18077 ( n11345,n18306,n18307 );
   xor U18078 ( n18307,si_23_,n18308 );
   nand U18079 ( n18304,n17407,p2_datao_reg_23_ );
   or U18080 ( n17524,n17728,n17727 );
   xor U18081 ( n17727,n17808,n18309 );
   nand U18082 ( n18309,n18310,n18311 );
   nand U18083 ( n18311,n17811,n14771 );
   nand U18084 ( n18310,n17805,n14515 );
   nand U18085 ( n17728,n18312,n18313 );
   nand U18086 ( n18313,n17805,n14771 );
   nand U18087 ( n14771,n18314,n18315 );
   nand U18088 ( n18315,n17402,n11364 );
   xor U18089 ( n11364,n18316,n18317 );
   xor U18090 ( n18317,si_25_,n18318 );
   nand U18091 ( n18314,n17407,p2_datao_reg_25_ );
   nand U18092 ( n18312,n17806,n14515 );
   nand U18093 ( n14515,n18319,n18320,n18321,n18322 );
   nand U18094 ( n18322,n17827,n16147 );
   xor U18095 ( n16147,p1_reg3_reg_25_,n17932 );
   nand U18096 ( n18321,p1_reg0_reg_25_,n17398 );
   nand U18097 ( n18320,p1_reg1_reg_25_,n17399 );
   nand U18098 ( n18319,p1_reg2_reg_25_,n17397 );
   nand U18099 ( n17521,n18323,n18324,n18325 );
   xor U18100 ( n18325,n17631,n18326 );
   nand U18101 ( n18324,n17805,n14759 );
   nand U18102 ( n17522,n18327,n18328,n18329 );
   nand U18103 ( n18326,n18330,n18331 );
   nand U18104 ( n18331,n17811,n14759 );
   nand U18105 ( n18330,n17805,n14512 );
   nand U18106 ( n18328,n18323,n18332 );
   nand U18107 ( n18323,n17806,n14512 );
   nand U18108 ( n14512,n18333,n18334,n18335,n18336 );
   nand U18109 ( n18336,n17525,n17827 );
   not U18110 ( n17525,n16173 );
   nand U18111 ( n16173,n17829,n18337 );
   nand U18112 ( n18337,n18338,n17516 );
   nand U18113 ( n18335,p1_reg0_reg_26_,n17398 );
   nand U18114 ( n18334,p1_reg1_reg_26_,n17399 );
   nand U18115 ( n18333,p1_reg2_reg_26_,n17397 );
   nand U18116 ( n18327,n16172,n18339 );
   not U18117 ( n16172,n14759 );
   nand U18118 ( n14759,n18340,n18341 );
   nand U18119 ( n18341,n17402,n11371 );
   xor U18120 ( n11371,n18342,n18343 );
   xor U18121 ( n18343,si_26_,n18344 );
   nand U18122 ( n18340,n17407,p2_datao_reg_26_ );
   nor U18123 ( n17909,n17795,n17800 );
   nor U18124 ( n17800,n18345,n18346 );
   not U18125 ( n17795,n17798 );
   nand U18126 ( n17798,n18346,n18345 );
   nand U18127 ( n18345,n18347,n18348 );
   nand U18128 ( n18348,n17805,n14746 );
   nand U18129 ( n18347,n17806,n14509 );
   xor U18130 ( n18346,n17808,n18349 );
   nand U18131 ( n18349,n18350,n18351 );
   nand U18132 ( n18351,n17811,n14746 );
   nand U18133 ( n14746,n18352,n18353 );
   nand U18134 ( n18353,n17402,n11380 );
   xor U18135 ( n11380,n17820,n18354 );
   xor U18136 ( n18354,si_27_,n17819 );
   nand U18137 ( n17819,n18355,n18356 );
   nand U18138 ( n18356,n18357,n18358 );
   not U18139 ( n18358,si_26_ );
   or U18140 ( n18357,n18344,n18342 );
   nand U18141 ( n18355,n18342,n18344 );
   nand U18142 ( n18344,n18359,n18360 );
   nand U18143 ( n18360,n18361,n18362 );
   not U18144 ( n18362,si_25_ );
   or U18145 ( n18361,n18318,n18316 );
   nand U18146 ( n18359,n18316,n18318 );
   nand U18147 ( n18318,n18363,n18364 );
   nand U18148 ( n18364,n18365,n18366 );
   not U18149 ( n18366,si_24_ );
   or U18150 ( n18365,n17926,n17924 );
   nand U18151 ( n18363,n17924,n17926 );
   nand U18152 ( n17926,n18367,n18368 );
   nand U18153 ( n18368,n18369,n18370 );
   not U18154 ( n18370,si_23_ );
   or U18155 ( n18369,n18308,n18306 );
   nand U18156 ( n18367,n18306,n18308 );
   nand U18157 ( n18308,n18371,n18372 );
   nand U18158 ( n18372,n18373,n18374 );
   not U18159 ( n18374,si_22_ );
   or U18160 ( n18373,n18290,n18288 );
   nand U18161 ( n18371,n18288,n18290 );
   nand U18162 ( n18290,n18375,n18376 );
   nand U18163 ( n18376,n18377,n18378 );
   not U18164 ( n18378,si_21_ );
   or U18165 ( n18377,n17958,n17956 );
   nand U18166 ( n18375,n17956,n17958 );
   nand U18167 ( n17958,n18379,n18380 );
   nand U18168 ( n18380,n18381,n18382 );
   not U18169 ( n18382,si_20_ );
   or U18170 ( n18381,n18273,n18271 );
   nand U18171 ( n18379,n18271,n18273 );
   nand U18172 ( n18273,n18383,n18384 );
   nand U18173 ( n18384,n18385,n18386 );
   not U18174 ( n18386,si_19_ );
   or U18175 ( n18385,n18260,n18258 );
   nand U18176 ( n18383,n18258,n18260 );
   nand U18177 ( n18260,n18387,n18388 );
   nand U18178 ( n18388,n18389,n18390 );
   not U18179 ( n18390,si_18_ );
   or U18180 ( n18389,n18242,n18240 );
   nand U18181 ( n18387,n18240,n18242 );
   nand U18182 ( n18242,n18391,n18392 );
   nand U18183 ( n18392,n18393,n17994 );
   not U18184 ( n17994,si_17_ );
   or U18185 ( n18393,n17993,n17992 );
   nand U18186 ( n18391,n17992,n17993 );
   nand U18187 ( n17993,n18394,n18395 );
   nand U18188 ( n18395,n18396,n18018 );
   not U18189 ( n18018,si_16_ );
   or U18190 ( n18396,n18017,n18016 );
   nand U18191 ( n18394,n18016,n18017 );
   nand U18192 ( n18017,n18397,n18398 );
   nand U18193 ( n18398,n18399,n18227 );
   not U18194 ( n18227,si_15_ );
   nand U18195 ( n18399,n18226,n18228 );
   or U18196 ( n18397,n18228,n18226 );
   nand U18197 ( n18226,n18400,n18401 );
   nand U18198 ( n18401,n11414,p1_datao_reg_15_ );
   nand U18199 ( n18400,n11416,p2_datao_reg_15_ );
   nand U18200 ( n18228,n18402,n18403,n18404 );
   or U18201 ( n18404,n18206,n18405 );
   nand U18202 ( n18403,n18406,n18407 );
   or U18203 ( n18407,n18203,si_14_ );
   not U18204 ( n18203,n18405 );
   not U18205 ( n18406,n18207 );
   nand U18206 ( n18207,n18185,n18164,n18064,n18057 );
   nand U18207 ( n18164,n18408,n18409 );
   nand U18208 ( n18409,si_10_,n18410 );
   or U18209 ( n18410,n18151,n18149 );
   nand U18210 ( n18408,n18149,n18151 );
   nand U18211 ( n18151,n18125,n18411 );
   nand U18212 ( n18411,n18124,n18126 );
   nand U18213 ( n18126,n18412,n18413,n18414 );
   not U18214 ( n18414,si_9_ );
   nand U18215 ( n18413,n11414,p1_datao_reg_9_ );
   nand U18216 ( n18412,n11416,p2_datao_reg_9_ );
   nand U18217 ( n18124,n18111,n18415 );
   nand U18218 ( n18415,n18110,n18112 );
   nand U18219 ( n18112,n18416,n18417,n18418 );
   not U18220 ( n18418,si_8_ );
   nand U18221 ( n18417,n11414,p1_datao_reg_8_ );
   nand U18222 ( n18416,n11416,p2_datao_reg_8_ );
   nand U18223 ( n18110,n18419,n18420 );
   nand U18224 ( n18420,n18421,n18422 );
   nand U18225 ( n18111,n18423,n18424,si_8_ );
   or U18226 ( n18424,n11414,p2_datao_reg_8_ );
   nand U18227 ( n18423,n11414,n14137 );
   not U18228 ( n14137,p1_datao_reg_8_ );
   nand U18229 ( n18125,n18425,n18426,si_9_ );
   or U18230 ( n18426,n11414,p2_datao_reg_9_ );
   nand U18231 ( n18425,n11414,n14121 );
   not U18232 ( n14121,p1_datao_reg_9_ );
   and U18233 ( n18149,n18427,n18428 );
   or U18234 ( n18428,n11414,p2_datao_reg_10_ );
   or U18235 ( n18427,n11416,p1_datao_reg_10_ );
   not U18236 ( n18185,n18165 );
   nor U18237 ( n18165,n18429,si_11_ );
   nand U18238 ( n18402,si_14_,n18430 );
   nand U18239 ( n18430,n18405,n18206 );
   nand U18240 ( n18206,n18057,n18431 );
   nand U18241 ( n18431,n18056,n18061,n18432 );
   nand U18242 ( n18432,n18166,n18064 );
   nand U18243 ( n18064,n18433,n18434,n18435 );
   not U18244 ( n18435,si_12_ );
   nand U18245 ( n18434,n11414,p1_datao_reg_12_ );
   nand U18246 ( n18433,n11416,p2_datao_reg_12_ );
   not U18247 ( n18166,n18183 );
   nand U18248 ( n18183,si_11_,n18429 );
   nand U18249 ( n18429,n18436,n18437 );
   nand U18250 ( n18437,n11414,p1_datao_reg_11_ );
   nand U18251 ( n18436,n11416,p2_datao_reg_11_ );
   nand U18252 ( n18061,n18438,n18439,si_12_ );
   or U18253 ( n18439,n11414,p2_datao_reg_12_ );
   nand U18254 ( n18438,n11414,n14170 );
   not U18255 ( n14170,p1_datao_reg_12_ );
   nand U18256 ( n18056,si_13_,n18060 );
   or U18257 ( n18057,n18060,si_13_ );
   and U18258 ( n18060,n18440,n18441 );
   or U18259 ( n18441,n11414,p2_datao_reg_13_ );
   or U18260 ( n18440,n11416,p1_datao_reg_13_ );
   nand U18261 ( n18405,n18442,n18443 );
   or U18262 ( n18443,n11414,p2_datao_reg_14_ );
   or U18263 ( n18442,n11416,p1_datao_reg_14_ );
   nand U18264 ( n18016,n18444,n18445 );
   or U18265 ( n18445,n11414,p2_datao_reg_16_ );
   nand U18266 ( n18444,n11414,n14203 );
   not U18267 ( n14203,p1_datao_reg_16_ );
   nand U18268 ( n17992,n18446,n18447 );
   or U18269 ( n18447,n11414,p2_datao_reg_17_ );
   nand U18270 ( n18446,n11414,n14060 );
   not U18271 ( n14060,p1_datao_reg_17_ );
   nand U18272 ( n18240,n18448,n18449 );
   or U18273 ( n18449,n11414,p2_datao_reg_18_ );
   nand U18274 ( n18448,n11414,n14224 );
   not U18275 ( n14224,p1_datao_reg_18_ );
   nand U18276 ( n18258,n18450,n18451 );
   or U18277 ( n18451,n11414,p2_datao_reg_19_ );
   nand U18278 ( n18450,n11414,n14229 );
   not U18279 ( n14229,p1_datao_reg_19_ );
   nand U18280 ( n18271,n18452,n18453 );
   or U18281 ( n18453,n11414,p2_datao_reg_20_ );
   nand U18282 ( n18452,n11414,n14238 );
   not U18283 ( n14238,p1_datao_reg_20_ );
   nand U18284 ( n17956,n18454,n18455 );
   or U18285 ( n18455,n11414,p2_datao_reg_21_ );
   nand U18286 ( n18454,n11414,n14032 );
   not U18287 ( n14032,p1_datao_reg_21_ );
   nand U18288 ( n18288,n18456,n18457 );
   or U18289 ( n18457,n11414,p2_datao_reg_22_ );
   nand U18290 ( n18456,n11414,n14254 );
   not U18291 ( n14254,p1_datao_reg_22_ );
   nand U18292 ( n18306,n18458,n18459 );
   or U18293 ( n18459,n11414,p2_datao_reg_23_ );
   nand U18294 ( n18458,n11414,n14022 );
   not U18295 ( n14022,p1_datao_reg_23_ );
   nand U18296 ( n17924,n18460,n18461 );
   or U18297 ( n18461,n11414,p2_datao_reg_24_ );
   nand U18298 ( n18460,n11414,n14263 );
   not U18299 ( n14263,p1_datao_reg_24_ );
   nand U18300 ( n18316,n18462,n18463 );
   or U18301 ( n18463,n11414,p2_datao_reg_25_ );
   nand U18302 ( n18462,n11414,n14279 );
   not U18303 ( n14279,p1_datao_reg_25_ );
   nand U18304 ( n18342,n18464,n18465 );
   or U18305 ( n18465,n11414,p2_datao_reg_26_ );
   nand U18306 ( n18464,n11414,n14290 );
   not U18307 ( n14290,p1_datao_reg_26_ );
   nand U18308 ( n17820,n18466,n18467 );
   or U18309 ( n18467,n11414,p2_datao_reg_27_ );
   nand U18310 ( n18466,n11414,n14010 );
   not U18311 ( n14010,p1_datao_reg_27_ );
   nand U18312 ( n18352,n17407,p2_datao_reg_27_ );
   nand U18313 ( n18350,n17805,n14509 );
   nand U18314 ( n14509,n18468,n18469,n18470,n18471 );
   nand U18315 ( n18471,n17827,n16217 );
   nand U18316 ( n18470,p1_reg0_reg_27_,n17398 );
   nand U18317 ( n18469,p1_reg1_reg_27_,n17399 );
   nand U18318 ( n18468,p1_reg2_reg_27_,n17397 );
   nand U18319 ( n17896,n16217,n17526 );
   nand U18320 ( n17526,n18472,n18473 );
   nand U18321 ( n18472,n18474,p1_state_reg );
   xor U18322 ( n16217,n17828,n17829 );
   or U18323 ( n17829,n17516,n18338 );
   nand U18324 ( n18338,p1_reg3_reg_25_,n17932 );
   nor U18325 ( n17932,n17877,n18296,n17666 );
   not U18326 ( n17666,p1_reg3_reg_24_ );
   not U18327 ( n18296,n17934 );
   nor U18328 ( n17934,n17749,n18279,n17589 );
   not U18329 ( n17589,p1_reg3_reg_22_ );
   not U18330 ( n18279,n17963 );
   nor U18331 ( n17963,n17837,n18248,n17618 );
   not U18332 ( n17618,p1_reg3_reg_20_ );
   not U18333 ( n18248,n18265 );
   nor U18334 ( n18265,n17679,n17999,n17548 );
   not U18335 ( n17548,p1_reg3_reg_18_ );
   nand U18336 ( n17999,p1_reg3_reg_15_,n18026,p1_reg3_reg_16_ );
   nor U18337 ( n18026,n17603,n18069,n17890 );
   not U18338 ( n17890,p1_reg3_reg_14_ );
   nand U18339 ( n18069,p1_reg3_reg_11_,n18139,p1_reg3_reg_12_ );
   nor U18340 ( n18139,n17864,n18475,n17640 );
   not U18341 ( n17640,p1_reg3_reg_9_ );
   not U18342 ( n17864,p1_reg3_reg_10_ );
   not U18343 ( n17603,p1_reg3_reg_13_ );
   not U18344 ( n17679,p1_reg3_reg_17_ );
   not U18345 ( n17837,p1_reg3_reg_19_ );
   not U18346 ( n17749,p1_reg3_reg_21_ );
   not U18347 ( n17877,p1_reg3_reg_23_ );
   not U18348 ( n17516,p1_reg3_reg_26_ );
   not U18349 ( n17828,p1_reg3_reg_27_ );
   nor U18350 ( n18479,n16757,n18480,n18481 );
   nor U18351 ( n18481,n15001,n17515 );
   nor U18352 ( n17507,n18482,n16275,n18483 );
   not U18353 ( n16275,n16426 );
   not U18354 ( n15001,n14572 );
   nor U18355 ( n18480,n14977,n17497 );
   nor U18356 ( n17576,n16426,n18482,n18483 );
   not U18357 ( n14977,n14566 );
   nand U18358 ( n14566,n18484,n18485,n18486,n18487 );
   nand U18359 ( n18487,n18488,n17827 );
   not U18360 ( n18488,n15599 );
   nand U18361 ( n15599,n18489,n18475 );
   not U18362 ( n18475,n18131 );
   nor U18363 ( n18131,n18490,n18491,n17774 );
   nand U18364 ( n18489,n17774,n18492 );
   nand U18365 ( n18492,p1_reg3_reg_7_,n18493 );
   not U18366 ( n17774,p1_reg3_reg_8_ );
   nand U18367 ( n18486,p1_reg0_reg_8_,n17398 );
   nand U18368 ( n18485,p1_reg1_reg_8_,n17399 );
   nand U18369 ( n18484,p1_reg2_reg_8_,n17397 );
   nor U18370 ( n16757,p1_state_reg,n18490 );
   not U18371 ( n18490,p1_reg3_reg_7_ );
   nand U18372 ( n18478,n15559,n17535 );
   nand U18373 ( n17535,n18494,n18473 );
   nand U18374 ( n18473,n18495,p1_state_reg );
   nand U18375 ( n18495,n16967,n18496,n16434,n17488 );
   not U18376 ( n16434,n15065 );
   nor U18377 ( n15065,n16274,n15066 );
   not U18378 ( n16274,n16428 );
   nand U18379 ( n18496,n18497,n18482 );
   nand U18380 ( n18494,n18474,n15061 );
   and U18381 ( n18474,n18482,n18498 );
   nand U18382 ( n18498,n18483,n16431 );
   not U18383 ( n16431,n18499 );
   nand U18384 ( n18483,n16979,n15061,n18500 );
   not U18385 ( n18500,n16960 );
   nand U18386 ( n18477,n18501,n18502,n17517 );
   not U18387 ( n17517,n17502 );
   nand U18388 ( n17502,n15061,n18497,n18503 );
   nand U18389 ( n18497,n18504,n18505,n18506 );
   and U18390 ( n18506,n16430,n15491,n15498 );
   not U18391 ( n15498,n15620 );
   nor U18392 ( n15620,n16960,n16979 );
   nor U18393 ( n15616,n16961,n17441 );
   nand U18394 ( n16430,n14699,n16454 );
   nand U18395 ( n14756,n18507,n17286 );
   or U18396 ( n18505,n17441,n16957 );
   nor U18397 ( n16957,n15095,n16059 );
   nor U18398 ( n16059,n18508,n18509 );
   nand U18399 ( n15095,n15495,n15493 );
   nor U18400 ( n15572,n17286,n18509,n16454 );
   nand U18401 ( n18504,n18509,n16962 );
   nand U18402 ( n16962,n15109,n16411 );
   nor U18403 ( n15109,n15573,n15437 );
   nor U18404 ( n15437,n18508,n17362 );
   nand U18405 ( n18502,n18095,n18510 );
   nand U18406 ( n18510,n18096,n18094 );
   not U18407 ( n18095,n18511 );
   nand U18408 ( n18501,n18096,n18094,n18511 );
   nand U18409 ( n18511,n18512,n18513 );
   nand U18410 ( n18513,n17539,n18514 );
   nand U18411 ( n18514,n17540,n17538 );
   and U18412 ( n17539,n18515,n18516 );
   nand U18413 ( n18516,n17696,n18517 );
   nand U18414 ( n18517,n18518,n17697 );
   xor U18415 ( n17696,n17631,n18519 );
   nand U18416 ( n18519,n18520,n18521 );
   nand U18417 ( n18521,n17811,n15002 );
   nand U18418 ( n18520,n17805,n14575 );
   or U18419 ( n18515,n17697,n18518 );
   not U18420 ( n18518,n17698 );
   nand U18421 ( n17698,n18522,n18523 );
   nand U18422 ( n18523,n17658,n18524 );
   or U18423 ( n18524,n17657,n17656 );
   and U18424 ( n17658,n18525,n18526 );
   nand U18425 ( n18526,n17805,n15468 );
   nand U18426 ( n18525,n17806,n14578 );
   nand U18427 ( n18522,n17656,n17657 );
   nand U18428 ( n17657,n18527,n17855 );
   nand U18429 ( n17855,n18528,n18529 );
   not U18430 ( n18529,n18530 );
   xor U18431 ( n18528,n17631,n18531 );
   nand U18432 ( n18527,n17852,n17854 );
   nand U18433 ( n17854,n18532,n18530 );
   nand U18434 ( n18530,n18533,n18534 );
   nand U18435 ( n18534,n17805,n15443 );
   nand U18436 ( n18533,n17806,n14581 );
   nand U18437 ( n18531,n18535,n18536 );
   nand U18438 ( n18536,n17811,n15443 );
   nand U18439 ( n15443,n18537,n18538,n18539 );
   nand U18440 ( n18539,n17407,p2_datao_reg_3_ );
   nand U18441 ( n18538,n16867,n16427 );
   not U18442 ( n16867,n16887 );
   nand U18443 ( n16887,n18540,n18541 );
   or U18444 ( n18541,p1_ir_reg_31_,p1_ir_reg_3_ );
   or U18445 ( n18540,n15146,n17990 );
   xor U18446 ( n15146,p1_ir_reg_3_,n15141 );
   nand U18447 ( n18537,n17402,n11178 );
   xor U18448 ( n11178,n18542,n18543 );
   xor U18449 ( n18542,n18544,n18545 );
   nand U18450 ( n18544,n18546,n18547 );
   nand U18451 ( n18547,n18548,n18549 );
   nand U18452 ( n18535,n17805,n14581 );
   nand U18453 ( n14581,n18550,n18551,n18552,n18553 );
   nand U18454 ( n18553,p1_reg0_reg_3_,n17398 );
   nand U18455 ( n18552,p1_reg1_reg_3_,n17399 );
   nand U18456 ( n18551,p1_reg2_reg_3_,n17397 );
   nand U18457 ( n18550,n17827,n17849 );
   not U18458 ( n17852,n17856 );
   nand U18459 ( n17856,n18554,n18555 );
   nand U18460 ( n18555,n17563,n18556 );
   nand U18461 ( n18556,n18557,n17565 );
   xor U18462 ( n17563,n17808,n18558 );
   nand U18463 ( n18558,n18559,n18560 );
   nand U18464 ( n18560,n17811,n15036 );
   nand U18465 ( n18559,n17805,n14584 );
   or U18466 ( n18554,n17565,n18557 );
   not U18467 ( n18557,n17564 );
   nand U18468 ( n17564,n18561,n18562 );
   nand U18469 ( n18562,n17805,n15036 );
   nand U18470 ( n15036,n18563,n18564,n18565 );
   nand U18471 ( n18565,n17407,p2_datao_reg_2_ );
   nand U18472 ( n18564,n16902,n16427 );
   not U18473 ( n16902,n16899 );
   nand U18474 ( n16899,n18566,n18567 );
   or U18475 ( n18567,p1_ir_reg_2_,p1_ir_reg_31_ );
   nand U18476 ( n18566,p1_ir_reg_31_,n18568 );
   nand U18477 ( n18568,n15140,n15141 );
   nand U18478 ( n15140,p1_ir_reg_2_,n18569 );
   nand U18479 ( n18569,n16918,n18570 );
   not U18480 ( n16918,p1_ir_reg_0_ );
   nand U18481 ( n18563,n17402,n11172 );
   nand U18482 ( n11172,n18571,n18572,n18573 );
   nand U18483 ( n18573,n18574,n18549 );
   nand U18484 ( n18572,n18575,n18576,si_2_ );
   nand U18485 ( n18571,n18577,n18578 );
   xor U18486 ( n18577,n18576,n18575 );
   not U18487 ( n18575,n18549 );
   nand U18488 ( n18561,n17806,n14584 );
   nand U18489 ( n14584,n18579,n18580,n18581,n18582 );
   nand U18490 ( n18582,p1_reg0_reg_2_,n17398 );
   nand U18491 ( n18581,p1_reg1_reg_2_,n17399 );
   nand U18492 ( n18580,p1_reg2_reg_2_,n17397 );
   nand U18493 ( n18579,p1_reg3_reg_2_,n17827 );
   nand U18494 ( n17565,n18583,n18584 );
   nand U18495 ( n18584,n17765,n18585 );
   or U18496 ( n18585,n17767,n17766 );
   xor U18497 ( n17765,n17631,n18586 );
   nand U18498 ( n18586,n18587,n18588 );
   nand U18499 ( n18588,n17811,n15385 );
   nand U18500 ( n18587,n17805,n14587 );
   nand U18501 ( n18583,n17766,n17767 );
   nand U18502 ( n17767,n18589,n18590 );
   nand U18503 ( n18590,n17631,n18591 );
   nand U18504 ( n18591,n17633,n17632 );
   or U18505 ( n18589,n17633,n17632 );
   nand U18506 ( n17632,n18592,n18593,n18594 );
   nand U18507 ( n18594,p1_ir_reg_0_,n16966 );
   nand U18508 ( n18593,n17806,n14590 );
   nand U18509 ( n18592,n17805,n15056 );
   xor U18510 ( n17633,n17808,n18595 );
   nand U18511 ( n18595,n18596,n18597,n18598 );
   nand U18512 ( n18598,p1_reg1_reg_0_,n16966 );
   nand U18513 ( n18597,n17805,n14590 );
   nand U18514 ( n14590,n18599,n18600,n18601,n18602 );
   nand U18515 ( n18602,p1_reg0_reg_0_,n17398 );
   nand U18516 ( n18601,p1_reg1_reg_0_,n17399 );
   nand U18517 ( n18600,p1_reg2_reg_0_,n17397 );
   nand U18518 ( n18599,p1_reg3_reg_0_,n17827 );
   nand U18519 ( n18596,n17811,n15056 );
   nand U18520 ( n15056,n18603,n18604,n18605 );
   nand U18521 ( n18605,p1_ir_reg_0_,n16427 );
   nand U18522 ( n18604,n17402,n11159 );
   and U18523 ( n11159,n18606,n18607 );
   nand U18524 ( n18606,n18608,n18609 );
   nand U18525 ( n18603,n17407,p2_datao_reg_0_ );
   and U18526 ( n17766,n18610,n18611 );
   nand U18527 ( n18611,n17805,n15385 );
   nand U18528 ( n15385,n18612,n18613,n18614 );
   nand U18529 ( n18614,n17407,p2_datao_reg_1_ );
   nand U18530 ( n18613,n16935,n16427 );
   not U18531 ( n16935,n16938 );
   nand U18532 ( n16938,n18615,n18616 );
   nand U18533 ( n18616,n18570,n17990 );
   not U18534 ( n18570,p1_ir_reg_1_ );
   or U18535 ( n18615,n15135,n17990 );
   xor U18536 ( n15135,p1_ir_reg_0_,p1_ir_reg_1_ );
   nand U18537 ( n18612,n17402,n11165 );
   xor U18538 ( n11165,n18617,n18618 );
   xor U18539 ( n18617,si_1_,n18607 );
   nand U18540 ( n18610,n17806,n14587 );
   nand U18541 ( n14587,n18619,n18620,n18621,n18622 );
   nand U18542 ( n18622,p1_reg0_reg_1_,n17398 );
   nand U18543 ( n18621,p1_reg1_reg_1_,n17399 );
   nand U18544 ( n18620,p1_reg2_reg_1_,n17397 );
   nand U18545 ( n18619,p1_reg3_reg_1_,n17827 );
   xor U18546 ( n17656,n17631,n18623 );
   nand U18547 ( n18623,n18624,n18625 );
   nand U18548 ( n18625,n17811,n15468 );
   nand U18549 ( n15468,n18626,n18627,n18628 );
   nand U18550 ( n18628,n17407,p2_datao_reg_4_ );
   nand U18551 ( n18627,n17402,n11185 );
   xor U18552 ( n11185,n18629,n18630 );
   and U18553 ( n18629,n18631,n18632 );
   nand U18554 ( n18626,n16852,n16427 );
   and U18555 ( n16852,n18633,n18634 );
   or U18556 ( n18634,p1_ir_reg_31_,p1_ir_reg_4_ );
   nand U18557 ( n18633,p1_ir_reg_31_,n18635 );
   nand U18558 ( n18635,n15152,n15151 );
   nand U18559 ( n15151,p1_ir_reg_4_,n18636 );
   nand U18560 ( n18624,n17805,n14578 );
   nand U18561 ( n14578,n18637,n18638,n18639,n18640 );
   nand U18562 ( n18640,n15470,n17827 );
   and U18563 ( n15470,n18641,n18642 );
   nand U18564 ( n18641,n17653,n17849 );
   nand U18565 ( n18639,p1_reg0_reg_4_,n17398 );
   nand U18566 ( n18638,p1_reg1_reg_4_,n17399 );
   nand U18567 ( n18637,p1_reg2_reg_4_,n17397 );
   nand U18568 ( n17697,n18643,n18644 );
   nand U18569 ( n18644,n17805,n15002 );
   nand U18570 ( n15002,n18645,n18646,n18647 );
   nand U18571 ( n18647,n17407,p2_datao_reg_5_ );
   nand U18572 ( n18646,n17402,n11195 );
   xor U18573 ( n11195,n18648,n18649 );
   and U18574 ( n18648,n18650,n18651 );
   nand U18575 ( n18645,n16801,n16427 );
   not U18576 ( n16801,n16800 );
   nand U18577 ( n16800,n18652,n18653,n18654 );
   nand U18578 ( n18653,n17990,n15161 );
   nand U18579 ( n18652,p1_ir_reg_31_,n15152,p1_ir_reg_5_ );
   not U18580 ( n15152,n15160 );
   nand U18581 ( n18643,n17806,n14575 );
   nand U18582 ( n14575,n18655,n18656,n18657,n18658 );
   nand U18583 ( n18658,n17827,n15482 );
   xor U18584 ( n15482,p1_reg3_reg_5_,n18659 );
   nand U18585 ( n18657,p1_reg0_reg_5_,n17398 );
   nand U18586 ( n18656,p1_reg1_reg_5_,n17399 );
   nand U18587 ( n18655,p1_reg2_reg_5_,n17397 );
   or U18588 ( n18512,n17538,n17540 );
   and U18589 ( n17540,n18660,n18661 );
   nand U18590 ( n18661,n17805,n14990 );
   nand U18591 ( n18660,n17806,n14572 );
   xor U18592 ( n17538,n17631,n18662 );
   nand U18593 ( n18662,n18663,n18664 );
   nand U18594 ( n18664,n17811,n14990 );
   nand U18595 ( n14990,n18665,n18666,n18667 );
   nand U18596 ( n18667,n17407,p2_datao_reg_6_ );
   nand U18597 ( n18666,n16788,n16427 );
   not U18598 ( n16788,n16805 );
   nand U18599 ( n16805,n18668,n18669 );
   or U18600 ( n18669,p1_ir_reg_31_,p1_ir_reg_6_ );
   nand U18601 ( n18668,p1_ir_reg_31_,n18670 );
   nand U18602 ( n18670,n15166,n15167 );
   nand U18603 ( n15166,p1_ir_reg_6_,n18654 );
   nand U18604 ( n18665,n17402,n11202 );
   xor U18605 ( n11202,n18671,n18672 );
   xor U18606 ( n18671,n18673,si_6_ );
   nand U18607 ( n18663,n17805,n14572 );
   nand U18608 ( n14572,n18674,n18675,n18676,n18677 );
   nand U18609 ( n18677,p1_reg0_reg_6_,n17398 );
   nand U18610 ( n18676,p1_reg1_reg_6_,n17399 );
   nand U18611 ( n18675,p1_reg2_reg_6_,n17397 );
   nand U18612 ( n18674,n17534,n17827 );
   not U18613 ( n17534,n15522 );
   nand U18614 ( n15522,n18678,n18491 );
   not U18615 ( n18491,n18493 );
   nand U18616 ( n18678,n17533,n18679 );
   nand U18617 ( n18679,p1_reg3_reg_5_,n18659 );
   nand U18618 ( n18094,n18680,n18681 );
   not U18619 ( n18681,n18682 );
   xor U18620 ( n18680,n17631,n18683 );
   nand U18621 ( n18096,n18684,n18682 );
   nand U18622 ( n18682,n18685,n18686 );
   nand U18623 ( n18686,n17806,n14569 );
   nand U18624 ( n18685,n17805,n14978 );
   nand U18625 ( n18683,n18688,n18689 );
   nand U18626 ( n18689,n17805,n14569 );
   nand U18627 ( n14569,n18690,n18691,n18692,n18693 );
   nand U18628 ( n18693,n17827,n15559 );
   xor U18629 ( n15559,p1_reg3_reg_7_,n18493 );
   nor U18630 ( n18493,n17693,n18642,n17533 );
   not U18631 ( n17533,p1_reg3_reg_6_ );
   not U18632 ( n18642,n18659 );
   nor U18633 ( n18659,n17653,n17849 );
   not U18634 ( n17849,p1_reg3_reg_3_ );
   not U18635 ( n17653,p1_reg3_reg_4_ );
   not U18636 ( n17693,p1_reg3_reg_5_ );
   nand U18637 ( n18692,p1_reg0_reg_7_,n17398 );
   nand U18638 ( n18691,p1_reg1_reg_7_,n17399 );
   nand U18639 ( n18690,p1_reg2_reg_7_,n17397 );
   xor U18640 ( n18695,p1_ir_reg_31_,p1_ir_reg_30_ );
   not U18641 ( n18696,n18694 );
   xor U18642 ( n18694,p1_ir_reg_31_,p1_ir_reg_29_ );
   nand U18643 ( n18332,n18697,n17488 );
   nand U18644 ( n18697,n16960,n16411 );
   nand U18645 ( n16411,n16443,n17441,n17286 );
   nand U18646 ( n16960,n15066,n17441 );
   nand U18647 ( n18688,n17811,n14978 );
   nand U18648 ( n18687,n18507,n17488 );
   nand U18649 ( n18339,n18698,n17488 );
   nand U18650 ( n18698,n17288,n16961,n18508,n15404 );
   nor U18651 ( n15573,n16980,n16454 );
   nand U18652 ( n16980,n17289,n17441 );
   not U18653 ( n18508,n17291 );
   nand U18654 ( n16961,n15066,n16979 );
   nor U18655 ( n15066,n17289,n16443 );
   nand U18656 ( n17288,n17362,n16443 );
   nand U18657 ( n18476,n17500,n14978 );
   nand U18658 ( n14978,n18699,n18700,n18701 );
   nand U18659 ( n18701,n17407,p2_datao_reg_7_ );
   nand U18660 ( n18700,n16742,n16427 );
   not U18661 ( n16742,n16741 );
   nand U18662 ( n16741,n18702,n18703,n18108 );
   nand U18663 ( n18703,n17990,n15175 );
   nand U18664 ( n18702,p1_ir_reg_31_,n15167,p1_ir_reg_7_ );
   not U18665 ( n15167,n15174 );
   nand U18666 ( n18699,n17402,n11211 );
   xor U18667 ( n11211,n18704,n18421 );
   nand U18668 ( n18421,n18705,n18706 );
   nand U18669 ( n18706,si_6_,n18707 );
   nand U18670 ( n18707,n18673,n18672 );
   or U18671 ( n18705,n18672,n18673 );
   and U18672 ( n18673,n18651,n18708 );
   nand U18673 ( n18708,n18649,n18650 );
   nand U18674 ( n18650,n18709,n18710,n18711 );
   not U18675 ( n18711,si_5_ );
   nand U18676 ( n18710,n11414,p1_datao_reg_5_ );
   nand U18677 ( n18709,n11416,p2_datao_reg_5_ );
   nand U18678 ( n18649,n18631,n18712 );
   nand U18679 ( n18712,n18630,n18632 );
   or U18680 ( n18632,n18713,si_4_ );
   nand U18681 ( n18630,n18714,n18715,n18716 );
   or U18682 ( n18716,n18546,n18543 );
   nand U18683 ( n18715,n18717,n18549,n18548 );
   nand U18684 ( n18548,n18576,n18578 );
   nand U18685 ( n18549,n18718,n18719 );
   nand U18686 ( n18719,si_1_,n18720 );
   nand U18687 ( n18720,n18618,n18607 );
   or U18688 ( n18718,n18607,n18618 );
   nand U18689 ( n18618,n18721,n18722 );
   or U18690 ( n18722,n11414,p2_datao_reg_1_ );
   or U18691 ( n18721,n11416,p1_datao_reg_1_ );
   or U18692 ( n18607,n18609,n18608 );
   and U18693 ( n18608,n18723,n18724 );
   nand U18694 ( n18724,n11414,p1_datao_reg_0_ );
   nand U18695 ( n18723,n11416,p2_datao_reg_0_ );
   not U18696 ( n18609,si_0_ );
   nand U18697 ( n18717,n18543,n18545 );
   not U18698 ( n18545,si_3_ );
   nand U18699 ( n18714,si_3_,n18725 );
   nand U18700 ( n18725,n18543,n18546 );
   not U18701 ( n18546,n18574 );
   nor U18702 ( n18574,n18578,n18576 );
   and U18703 ( n18576,n18726,n18727 );
   nand U18704 ( n18727,n11414,p1_datao_reg_2_ );
   nand U18705 ( n18726,n11416,p2_datao_reg_2_ );
   not U18706 ( n18578,si_2_ );
   nand U18707 ( n18543,n18728,n18729 );
   or U18708 ( n18729,n11414,p2_datao_reg_3_ );
   or U18709 ( n18728,n11416,p1_datao_reg_3_ );
   nand U18710 ( n18631,si_4_,n18713 );
   nand U18711 ( n18713,n18730,n18731 );
   nand U18712 ( n18731,n11414,p1_datao_reg_4_ );
   nand U18713 ( n18730,n11416,p2_datao_reg_4_ );
   nand U18714 ( n18651,n18732,n18733,si_5_ );
   or U18715 ( n18733,n11414,p2_datao_reg_5_ );
   nand U18716 ( n18732,n11414,n14351 );
   not U18717 ( n14351,p1_datao_reg_5_ );
   nand U18718 ( n18672,n18734,n18735 );
   or U18719 ( n18735,n11414,p2_datao_reg_6_ );
   or U18720 ( n18734,n11416,p1_datao_reg_6_ );
   and U18721 ( n18704,n18419,n18422 );
   or U18722 ( n18422,n18736,si_7_ );
   nand U18723 ( n18419,si_7_,n18736 );
   nand U18724 ( n18736,n18737,n18738 );
   nand U18725 ( n18738,n11414,p1_datao_reg_7_ );
   nand U18726 ( n18737,n11416,p2_datao_reg_7_ );
   or U18727 ( n18740,p1_addr_reg_19_,p1_rd_reg,p2_addr_reg_19_ );
   nand U18728 ( n18739,p1_addr_reg_19_,n10565,p2_addr_reg_19_ );
   not U18729 ( n10565,p2_rd_reg );
   nand U18730 ( n17575,n18741,n15061 );
   nor U18731 ( n15061,n16966,p1_u3084,n16963 );
   nand U18732 ( n18741,n16264,n18742 );
   nand U18733 ( n18742,n18503,n18499 );
   nor U18734 ( n18499,n17286,n14803 );
   nand U18735 ( n14698,n18743,n18744 );
   nand U18736 ( n18744,n17291,n18507 );
   nor U18737 ( n18507,n17441,n16979 );
   nor U18738 ( n17291,n16443,n17286 );
   nand U18739 ( n18743,n17012,n17362 );
   not U18740 ( n17286,n17289 );
   not U18741 ( n18503,n18482 );
   nand U18742 ( n18482,n14689,n15060,n15064 );
   and U18743 ( n15064,n15071,n18745 );
   nand U18744 ( n15071,n18746,n18747 );
   and U18745 ( n15060,n18748,n18749,n18750,n18751 );
   nor U18746 ( n18751,n18752,n18753,n18754,n18755 );
   not U18747 ( n15339,p1_d_reg_6_ );
   not U18748 ( n15341,p1_d_reg_13_ );
   not U18749 ( n15343,p1_d_reg_17_ );
   nor U18750 ( n18756,p1_d_reg_22_,p1_d_reg_24_,p1_d_reg_23_ );
   nor U18751 ( n18750,n18757,n18758,n18759,n18760 );
   not U18752 ( n15345,p1_d_reg_19_ );
   not U18753 ( n15342,p1_d_reg_16_ );
   nor U18754 ( n18761,p1_d_reg_7_,p1_d_reg_9_,p1_d_reg_8_ );
   not U18755 ( n15340,p1_d_reg_10_ );
   nor U18756 ( n18749,n18762,n18763,n18764,n18765 );
   not U18757 ( n15347,p1_d_reg_29_ );
   not U18758 ( n15338,p1_d_reg_2_ );
   not U18759 ( n15346,p1_d_reg_27_ );
   not U18760 ( n15344,p1_d_reg_18_ );
   nor U18761 ( n18748,n18766,n18767,n18768,n18769 );
   nor U18762 ( n18770,p1_d_reg_5_,p1_d_reg_4_,p1_d_reg_3_,p1_d_reg_30_ );
   nor U18763 ( n18771,p1_d_reg_20_,p1_d_reg_26_,p1_d_reg_25_ );
   nor U18764 ( n18772,p1_d_reg_15_,p1_d_reg_14_,p1_d_reg_12_,p1_d_reg_11_ );
   nor U18765 ( n18773,p1_d_reg_21_,p1_d_reg_31_,p1_d_reg_28_ );
   not U18766 ( n14689,n15059 );
   nand U18767 ( n15059,n15074,n18774 );
   nand U18768 ( n15348,n18775,n18776,n18777 );
   nand U18769 ( n18776,n18778,n16425 );
   not U18770 ( n16425,p1_b_reg );
   nand U18771 ( n18775,n18779,n18747,p1_b_reg );
   nand U18772 ( n15074,n18746,n18779 );
   nand U18773 ( n16264,n14717,n17362 );
   nand U18774 ( n17289,n18780,n18781 );
   nand U18775 ( n18781,p1_ir_reg_20_,n17990 );
   nand U18776 ( n18780,n15260,n15261,p1_ir_reg_31_ );
   nand U18777 ( n15260,p1_ir_reg_20_,n15255 );
   not U18778 ( n16454,n16443 );
   nand U18779 ( n16443,n18782,n18783 );
   nand U18780 ( n18783,p1_ir_reg_19_,n17990 );
   nand U18781 ( n18782,n15254,n15255,p1_ir_reg_31_ );
   nand U18782 ( n15254,p1_ir_reg_19_,n18239 );
   not U18783 ( n17488,n16966 );
   nor U18784 ( n16966,n18747,n18779,n18746 );
   not U18785 ( n18746,n18777 );
   nand U18786 ( n18777,n18785,n18786 );
   nand U18787 ( n18786,p1_ir_reg_26_,n17990 );
   nand U18788 ( n18785,n15302,n15303,p1_ir_reg_31_ );
   nand U18789 ( n15302,p1_ir_reg_26_,n18787 );
   nand U18790 ( n18787,n15296,n15297 );
   not U18791 ( n15297,p1_ir_reg_25_ );
   not U18792 ( n18779,n18778 );
   nand U18793 ( n18778,n18788,n18789 );
   nand U18794 ( n18789,p1_ir_reg_24_,n17990 );
   nand U18795 ( n18788,n15288,n15289,p1_ir_reg_31_ );
   nand U18796 ( n15288,p1_ir_reg_24_,n18790 );
   nand U18797 ( n18790,n15282,n15283 );
   not U18798 ( n15283,p1_ir_reg_23_ );
   xor U18799 ( n18747,p1_ir_reg_25_,n18791 );
   nand U18800 ( n18791,p1_ir_reg_31_,n15289 );
   nand U18801 ( n18784,n18792,p1_state_reg );
   nand U18802 ( n18792,n18793,n18794 );
   not U18803 ( n18794,n16427 );
   nand U18804 ( n16426,n18795,n18796 );
   nand U18805 ( n18796,p1_ir_reg_28_,n17990 );
   nand U18806 ( n18795,n15316,n15317,p1_ir_reg_31_ );
   not U18807 ( n15317,n15324 );
   nor U18808 ( n15324,p1_ir_reg_27_,p1_ir_reg_28_,n15303 );
   not U18809 ( n15303,n15310 );
   nand U18810 ( n15316,p1_ir_reg_28_,n18797 );
   nand U18811 ( n18797,n15310,n15311 );
   not U18812 ( n15311,p1_ir_reg_27_ );
   xor U18813 ( n16913,n18798,p1_ir_reg_27_ );
   nor U18814 ( n18798,n15310,n17990 );
   nor U18815 ( n15310,p1_ir_reg_25_,p1_ir_reg_26_,n15289 );
   not U18816 ( n15289,n15296 );
   nor U18817 ( n15296,p1_ir_reg_23_,p1_ir_reg_24_,n15275 );
   nand U18818 ( n18793,n16428,n16967 );
   not U18819 ( n16967,n16963 );
   xor U18820 ( n16963,n18799,p1_ir_reg_23_ );
   nor U18821 ( n18799,n15282,n17990 );
   nor U18822 ( n16428,n18509,n17362 );
   not U18823 ( n17362,n17441 );
   xor U18824 ( n17441,n15269,n18800 );
   nand U18825 ( n18800,p1_ir_reg_31_,n15261 );
   not U18826 ( n18509,n16979 );
   nand U18827 ( n16979,n18801,n18802 );
   nand U18828 ( n18802,p1_ir_reg_22_,n17990 );
   not U18829 ( n17990,p1_ir_reg_31_ );
   nand U18830 ( n18801,n15274,n15275,p1_ir_reg_31_ );
   not U18831 ( n15275,n15282 );
   nor U18832 ( n15282,p1_ir_reg_21_,p1_ir_reg_22_,n15261 );
   not U18833 ( n15261,n15268 );
   nand U18834 ( n15274,p1_ir_reg_22_,n18803 );
   nand U18835 ( n18803,n15268,n15269 );
   not U18836 ( n15269,p1_ir_reg_21_ );
   nor U18837 ( n15268,n15255,p1_ir_reg_20_ );
   or U18838 ( n15255,n18239,p1_ir_reg_19_ );
   nand U18839 ( n18239,n15247,n15249 );
   not U18840 ( n15249,p1_ir_reg_18_ );
   nor U18841 ( n15247,n15232,p1_ir_reg_17_ );
   not U18842 ( n15232,n15239 );
   nor U18843 ( n15239,n18014,p1_ir_reg_16_ );
   nand U18844 ( n18014,n15224,n15226 );
   not U18845 ( n15226,p1_ir_reg_15_ );
   nor U18846 ( n15224,n18051,p1_ir_reg_14_ );
   nand U18847 ( n18051,n15210,n15211 );
   not U18848 ( n15211,p1_ir_reg_13_ );
   nor U18849 ( n15210,p1_ir_reg_11_,p1_ir_reg_12_,n18146 );
   not U18850 ( n18146,n18181 );
   nor U18851 ( n18181,p1_ir_reg_10_,p1_ir_reg_9_,n15181 );
   not U18852 ( n15181,n18122 );
   nor U18853 ( n18122,n18108,p1_ir_reg_8_ );
   nand U18854 ( n18108,n15174,n15175 );
   not U18855 ( n15175,p1_ir_reg_7_ );
   nor U18856 ( n15174,n18654,p1_ir_reg_6_ );
   nand U18857 ( n18654,n15160,n15161 );
   not U18858 ( n15161,p1_ir_reg_5_ );
   nor U18859 ( n15160,n18636,p1_ir_reg_4_ );
   or U18860 ( n18636,n15141,p1_ir_reg_3_ );
   or U18861 ( n15141,p1_ir_reg_1_,p1_ir_reg_2_,p1_ir_reg_0_ );
   xor U18862 ( n18804,n16684,p2_addr_reg_10_ );
   xor U18863 ( n18806,n18808,p2_addr_reg_11_ );
   xor U18864 ( n18809,n16631,p2_addr_reg_12_ );
   xor U18865 ( n18811,n16610,p2_addr_reg_13_ );
   xor U18866 ( n18813,n18815,p2_addr_reg_14_ );
   xor U18867 ( n18816,n18818,p2_addr_reg_15_ );
   xor U18868 ( n18819,n18821,p2_addr_reg_16_ );
   xor U18869 ( n18822,n16507,p2_addr_reg_17_ );
   xor U18870 ( n18824,n18826,p2_addr_reg_18_ );
   xor U18871 ( n18827,n16898,p2_addr_reg_2_ );
   xor U18872 ( n18829,n16878,p2_addr_reg_3_ );
   xor U18873 ( n18831,p1_addr_reg_4_,n12959 );
   xor U18874 ( n18833,n16817,p2_addr_reg_5_ );
   xor U18875 ( n18835,n16787,p2_addr_reg_6_ );
   xor U18876 ( n18840,n16758,p2_addr_reg_7_ );
   xor U18877 ( n18842,n16732,p2_addr_reg_8_ );
   xor U18878 ( n18844,n16705,p2_addr_reg_9_ );
   nand U18879 ( n18847,n18848,n18849 );
   nand U18880 ( n18849,p2_addr_reg_18_,n18850 );
   nand U18881 ( n18850,n18826,n18825 );
   or U18882 ( n18848,n18825,n18826 );
   not U18883 ( n18826,p1_addr_reg_18_ );
   nand U18884 ( n18825,n18851,n18852 );
   nand U18885 ( n18852,n18853,n18854 );
   not U18886 ( n18854,p2_addr_reg_17_ );
   or U18887 ( n18853,n18823,n16507 );
   nand U18888 ( n18851,n18823,n16507 );
   not U18889 ( n16507,p1_addr_reg_17_ );
   nand U18890 ( n18823,n18855,n18856 );
   nand U18891 ( n18856,n18857,n18858 );
   not U18892 ( n18858,p2_addr_reg_16_ );
   or U18893 ( n18857,n18820,n18821 );
   nand U18894 ( n18855,n18820,n18821 );
   not U18895 ( n18821,p1_addr_reg_16_ );
   nand U18896 ( n18820,n18859,n18860 );
   nand U18897 ( n18860,n18861,n18862 );
   not U18898 ( n18862,p2_addr_reg_15_ );
   or U18899 ( n18861,n18817,n18818 );
   nand U18900 ( n18859,n18817,n18818 );
   not U18901 ( n18818,p1_addr_reg_15_ );
   nand U18902 ( n18817,n18863,n18864 );
   nand U18903 ( n18864,n18865,n18866 );
   not U18904 ( n18866,p2_addr_reg_14_ );
   or U18905 ( n18865,n18814,n18815 );
   nand U18906 ( n18863,n18814,n18815 );
   not U18907 ( n18815,p1_addr_reg_14_ );
   nand U18908 ( n18814,n18867,n18868 );
   nand U18909 ( n18868,n18869,n18870 );
   not U18910 ( n18870,p2_addr_reg_13_ );
   or U18911 ( n18869,n18812,n16610 );
   nand U18912 ( n18867,n18812,n16610 );
   not U18913 ( n16610,p1_addr_reg_13_ );
   nand U18914 ( n18812,n18871,n18872 );
   nand U18915 ( n18872,n18873,n12736 );
   not U18916 ( n12736,p2_addr_reg_12_ );
   or U18917 ( n18873,n18810,n16631 );
   nand U18918 ( n18871,n18810,n16631 );
   not U18919 ( n16631,p1_addr_reg_12_ );
   nand U18920 ( n18810,n18874,n18875 );
   nand U18921 ( n18875,n18876,n18877 );
   not U18922 ( n18877,p2_addr_reg_11_ );
   or U18923 ( n18876,n18807,n18808 );
   nand U18924 ( n18874,n18807,n18808 );
   not U18925 ( n18808,p1_addr_reg_11_ );
   nand U18926 ( n18807,n18878,n18879 );
   nand U18927 ( n18879,n18880,n18881 );
   not U18928 ( n18881,p2_addr_reg_10_ );
   or U18929 ( n18880,n18805,n16684 );
   nand U18930 ( n18878,n18805,n16684 );
   not U18931 ( n16684,p1_addr_reg_10_ );
   nand U18932 ( n18805,n18882,n18883 );
   nand U18933 ( n18883,n18884,n12819 );
   not U18934 ( n12819,p2_addr_reg_9_ );
   or U18935 ( n18884,n18845,n16705 );
   nand U18936 ( n18882,n18845,n16705 );
   not U18937 ( n16705,p1_addr_reg_9_ );
   nand U18938 ( n18845,n18885,n18886 );
   nand U18939 ( n18886,n18887,n18888 );
   not U18940 ( n18888,p2_addr_reg_8_ );
   or U18941 ( n18887,n18843,n16732 );
   nand U18942 ( n18885,n18843,n16732 );
   not U18943 ( n16732,p1_addr_reg_8_ );
   nand U18944 ( n18843,n18889,n18890 );
   nand U18945 ( n18890,n18891,n12871 );
   not U18946 ( n12871,p2_addr_reg_7_ );
   or U18947 ( n18891,n18841,n16758 );
   nand U18948 ( n18889,n18841,n16758 );
   not U18949 ( n16758,p1_addr_reg_7_ );
   nand U18950 ( n18841,n18892,n18893 );
   nand U18951 ( n18893,n18894,n12900 );
   not U18952 ( n12900,p2_addr_reg_6_ );
   or U18953 ( n18894,n18836,n16787 );
   nand U18954 ( n18892,n18836,n16787 );
   not U18955 ( n16787,p1_addr_reg_6_ );
   nand U18956 ( n18836,n18895,n18896 );
   nand U18957 ( n18896,n18897,n12930 );
   not U18958 ( n12930,p2_addr_reg_5_ );
   or U18959 ( n18897,n18834,n16817 );
   nand U18960 ( n18895,n18834,n16817 );
   not U18961 ( n16817,p1_addr_reg_5_ );
   nand U18962 ( n18834,n18898,n18899 );
   nand U18963 ( n18899,n18900,n12959 );
   not U18964 ( n12959,p2_addr_reg_4_ );
   nand U18965 ( n18900,n18901,p1_addr_reg_4_ );
   or U18966 ( n18898,n18901,p1_addr_reg_4_ );
   not U18967 ( n18901,n18832 );
   nand U18968 ( n18832,n18902,n18903 );
   nand U18969 ( n18903,n18904,n18905 );
   not U18970 ( n18905,p2_addr_reg_3_ );
   or U18971 ( n18904,n18830,n16878 );
   nand U18972 ( n18902,n18830,n16878 );
   not U18973 ( n16878,p1_addr_reg_3_ );
   nand U18974 ( n18830,n18906,n18907 );
   nand U18975 ( n18907,n18908,n18909 );
   not U18976 ( n18909,p2_addr_reg_2_ );
   or U18977 ( n18908,n18828,n16898 );
   nand U18978 ( n18906,n18828,n16898 );
   not U18979 ( n16898,p1_addr_reg_2_ );
   nand U18980 ( n18828,n18910,n18911 );
   nand U18981 ( n18911,n18912,n18839 );
   not U18982 ( n18839,p2_addr_reg_1_ );
   nand U18983 ( n18912,n18837,p1_addr_reg_1_ );
   not U18984 ( n18837,n18913 );
   nand U18985 ( n18910,n18913,n16934 );
   not U18986 ( n16934,p1_addr_reg_1_ );
   nand U18987 ( n18913,p1_addr_reg_0_,p2_addr_reg_0_ );
   xor U18988 ( n18846,p2_addr_reg_19_,p1_addr_reg_19_ );
endmodule
