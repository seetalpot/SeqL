
module b22 ( si_31_, si_30_, si_29_, si_28_, si_27_, si_26_, si_25_, si_24_,         si_23_, si_22_, si_21_, si_20_, si_19_, si_18_, si_17_, si_16_, si_15_,         si_14_, si_13_, si_12_, si_11_, si_10_, si_9_, si_8_, si_7_, si_6_,         si_5_, si_4_, si_3_, si_2_, si_1_, si_0_, p1_ir_reg_0_, p1_ir_reg_1_,         p1_ir_reg_2_, p1_ir_reg_3_, p1_ir_reg_4_, p1_ir_reg_5_, p1_ir_reg_6_,         p1_ir_reg_7_, p1_ir_reg_8_, p1_ir_reg_9_, p1_ir_reg_10_, p1_ir_reg_11_,         p1_ir_reg_12_, p1_ir_reg_13_, p1_ir_reg_14_, p1_ir_reg_15_,         p1_ir_reg_16_, p1_ir_reg_17_, p1_ir_reg_18_, p1_ir_reg_19_,         p1_ir_reg_20_, p1_ir_reg_21_, p1_ir_reg_22_, p1_ir_reg_23_,         p1_ir_reg_24_, p1_ir_reg_25_, p1_ir_reg_26_, p1_ir_reg_27_,         p1_ir_reg_28_, p1_ir_reg_29_, p1_ir_reg_30_, p1_ir_reg_31_,         p1_d_reg_0_, p1_d_reg_1_, p1_d_reg_2_, p1_d_reg_3_, p1_d_reg_4_,         p1_d_reg_5_, p1_d_reg_6_, p1_d_reg_7_, p1_d_reg_8_, p1_d_reg_9_,         p1_d_reg_10_, p1_d_reg_11_, p1_d_reg_12_, p1_d_reg_13_, p1_d_reg_14_,         p1_d_reg_15_, p1_d_reg_16_, p1_d_reg_17_, p1_d_reg_18_, p1_d_reg_19_,         p1_d_reg_20_, p1_d_reg_21_, p1_d_reg_22_, p1_d_reg_23_, p1_d_reg_24_,         p1_d_reg_25_, p1_d_reg_26_, p1_d_reg_27_, p1_d_reg_28_, p1_d_reg_29_,         p1_d_reg_30_, p1_d_reg_31_, p1_reg0_reg_0_, p1_reg0_reg_1_,         p1_reg0_reg_2_, p1_reg0_reg_3_, p1_reg0_reg_4_, p1_reg0_reg_5_,         p1_reg0_reg_6_, p1_reg0_reg_7_, p1_reg0_reg_8_, p1_reg0_reg_9_,         p1_reg0_reg_10_, p1_reg0_reg_11_, p1_reg0_reg_12_, p1_reg0_reg_13_,         p1_reg0_reg_14_, p1_reg0_reg_15_, p1_reg0_reg_16_, p1_reg0_reg_17_,         p1_reg0_reg_18_, p1_reg0_reg_19_, p1_reg0_reg_20_, p1_reg0_reg_21_,         p1_reg0_reg_22_, p1_reg0_reg_23_, p1_reg0_reg_24_, p1_reg0_reg_25_,         p1_reg0_reg_26_, p1_reg0_reg_27_, p1_reg0_reg_28_, p1_reg0_reg_29_,         p1_reg0_reg_30_, p1_reg0_reg_31_, p1_reg1_reg_0_, p1_reg1_reg_1_,         p1_reg1_reg_2_, p1_reg1_reg_3_, p1_reg1_reg_4_, p1_reg1_reg_5_,         p1_reg1_reg_6_, p1_reg1_reg_7_, p1_reg1_reg_8_, p1_reg1_reg_9_,         p1_reg1_reg_10_, p1_reg1_reg_11_, p1_reg1_reg_12_, p1_reg1_reg_13_,         p1_reg1_reg_14_, p1_reg1_reg_15_, p1_reg1_reg_16_, p1_reg1_reg_17_,         p1_reg1_reg_18_, p1_reg1_reg_19_, p1_reg1_reg_20_, p1_reg1_reg_21_,         p1_reg1_reg_22_, p1_reg1_reg_23_, p1_reg1_reg_24_, p1_reg1_reg_25_,         p1_reg1_reg_26_, p1_reg1_reg_27_, p1_reg1_reg_28_, p1_reg1_reg_29_,         p1_reg1_reg_30_, p1_reg1_reg_31_, p1_reg2_reg_0_, p1_reg2_reg_1_,         p1_reg2_reg_2_, p1_reg2_reg_3_, p1_reg2_reg_4_, p1_reg2_reg_5_,         p1_reg2_reg_6_, p1_reg2_reg_7_, p1_reg2_reg_8_, p1_reg2_reg_9_,         p1_reg2_reg_10_, p1_reg2_reg_11_, p1_reg2_reg_12_, p1_reg2_reg_13_,         p1_reg2_reg_14_, p1_reg2_reg_15_, p1_reg2_reg_16_, p1_reg2_reg_17_,         p1_reg2_reg_18_, p1_reg2_reg_19_, p1_reg2_reg_20_, p1_reg2_reg_21_,         p1_reg2_reg_22_, p1_reg2_reg_23_, p1_reg2_reg_24_, p1_reg2_reg_25_,         p1_reg2_reg_26_, p1_reg2_reg_27_, p1_reg2_reg_28_, p1_reg2_reg_29_,         p1_reg2_reg_30_, p1_reg2_reg_31_, p1_addr_reg_19_, p1_addr_reg_18_,         p1_addr_reg_17_, p1_addr_reg_16_, p1_addr_reg_15_, p1_addr_reg_14_,         p1_addr_reg_13_, p1_addr_reg_12_, p1_addr_reg_11_, p1_addr_reg_10_,         p1_addr_reg_9_, p1_addr_reg_8_, p1_addr_reg_7_, p1_addr_reg_6_,         p1_addr_reg_5_, p1_addr_reg_4_, p1_addr_reg_3_, p1_addr_reg_2_,         p1_addr_reg_1_, p1_addr_reg_0_, p1_datao_reg_0_, p1_datao_reg_1_,         p1_datao_reg_2_, p1_datao_reg_3_, p1_datao_reg_4_, p1_datao_reg_5_,         p1_datao_reg_6_, p1_datao_reg_7_, p1_datao_reg_8_, p1_datao_reg_9_,         p1_datao_reg_10_, p1_datao_reg_11_, p1_datao_reg_12_, p1_datao_reg_13_,         p1_datao_reg_14_, p1_datao_reg_15_, p1_datao_reg_16_, p1_datao_reg_17_,         p1_datao_reg_18_, p1_datao_reg_19_, p1_datao_reg_20_, p1_datao_reg_21_,         p1_datao_reg_22_, p1_datao_reg_23_, p1_datao_reg_24_, p1_datao_reg_25_,         p1_datao_reg_26_, p1_datao_reg_27_, p1_datao_reg_28_, p1_datao_reg_29_,         p1_datao_reg_30_, p1_datao_reg_31_, p1_b_reg, p1_reg3_reg_15_,         p1_reg3_reg_26_, p1_reg3_reg_6_, p1_reg3_reg_18_, p1_reg3_reg_2_,         p1_reg3_reg_11_, p1_reg3_reg_22_, p1_reg3_reg_13_, p1_reg3_reg_20_,         p1_reg3_reg_0_, p1_reg3_reg_9_, p1_reg3_reg_4_, p1_reg3_reg_24_,         p1_reg3_reg_17_, p1_reg3_reg_5_, p1_reg3_reg_16_, p1_reg3_reg_25_,         p1_reg3_reg_12_, p1_reg3_reg_21_, p1_reg3_reg_1_, p1_reg3_reg_8_,         p1_reg3_reg_28_, p1_reg3_reg_19_, p1_reg3_reg_3_, p1_reg3_reg_10_,         p1_reg3_reg_23_, p1_reg3_reg_14_, p1_reg3_reg_27_, p1_reg3_reg_7_,         p1_state_reg, p1_rd_reg, p1_wr_reg, p2_ir_reg_0_, p2_ir_reg_1_,         p2_ir_reg_2_, p2_ir_reg_3_, p2_ir_reg_4_, p2_ir_reg_5_, p2_ir_reg_6_,         p2_ir_reg_7_, p2_ir_reg_8_, p2_ir_reg_9_, p2_ir_reg_10_, p2_ir_reg_11_,         p2_ir_reg_12_, p2_ir_reg_13_, p2_ir_reg_14_, p2_ir_reg_15_,         p2_ir_reg_16_, p2_ir_reg_17_, p2_ir_reg_18_, p2_ir_reg_19_,         p2_ir_reg_20_, p2_ir_reg_21_, p2_ir_reg_22_, p2_ir_reg_23_,         p2_ir_reg_24_, p2_ir_reg_25_, p2_ir_reg_26_, p2_ir_reg_27_,         p2_ir_reg_28_, p2_ir_reg_29_, p2_ir_reg_30_, p2_ir_reg_31_,         p2_d_reg_0_, p2_d_reg_1_, p2_d_reg_2_, p2_d_reg_3_, p2_d_reg_4_,         p2_d_reg_5_, p2_d_reg_6_, p2_d_reg_7_, p2_d_reg_8_, p2_d_reg_9_,         p2_d_reg_10_, p2_d_reg_11_, p2_d_reg_12_, p2_d_reg_13_, p2_d_reg_14_,         p2_d_reg_15_, p2_d_reg_16_, p2_d_reg_17_, p2_d_reg_18_, p2_d_reg_19_,         p2_d_reg_20_, p2_d_reg_21_, p2_d_reg_22_, p2_d_reg_23_, p2_d_reg_24_,         p2_d_reg_25_, p2_d_reg_26_, p2_d_reg_27_, p2_d_reg_28_, p2_d_reg_29_,         p2_d_reg_30_, p2_d_reg_31_, p2_reg0_reg_0_, p2_reg0_reg_1_,         p2_reg0_reg_2_, p2_reg0_reg_3_, p2_reg0_reg_4_, p2_reg0_reg_5_,         p2_reg0_reg_6_, p2_reg0_reg_7_, p2_reg0_reg_8_, p2_reg0_reg_9_,         p2_reg0_reg_10_, p2_reg0_reg_11_, p2_reg0_reg_12_, p2_reg0_reg_13_,         p2_reg0_reg_14_, p2_reg0_reg_15_, p2_reg0_reg_16_, p2_reg0_reg_17_,         p2_reg0_reg_18_, p2_reg0_reg_19_, p2_reg0_reg_20_, p2_reg0_reg_21_,         p2_reg0_reg_22_, p2_reg0_reg_23_, p2_reg0_reg_24_, p2_reg0_reg_25_,         p2_reg0_reg_26_, p2_reg0_reg_27_, p2_reg0_reg_28_, p2_reg0_reg_29_,         p2_reg0_reg_30_, p2_reg0_reg_31_, p2_reg1_reg_0_, p2_reg1_reg_1_,         p2_reg1_reg_2_, p2_reg1_reg_3_, p2_reg1_reg_4_, p2_reg1_reg_5_,         p2_reg1_reg_6_, p2_reg1_reg_7_, p2_reg1_reg_8_, p2_reg1_reg_9_,         p2_reg1_reg_10_, p2_reg1_reg_11_, p2_reg1_reg_12_, p2_reg1_reg_13_,         p2_reg1_reg_14_, p2_reg1_reg_15_, p2_reg1_reg_16_, p2_reg1_reg_17_,         p2_reg1_reg_18_, p2_reg1_reg_19_, p2_reg1_reg_20_, p2_reg1_reg_21_,         p2_reg1_reg_22_, p2_reg1_reg_23_, p2_reg1_reg_24_, p2_reg1_reg_25_,         p2_reg1_reg_26_, p2_reg1_reg_27_, p2_reg1_reg_28_, p2_reg1_reg_29_,         p2_reg1_reg_30_, p2_reg1_reg_31_, p2_reg2_reg_0_, p2_reg2_reg_1_,         p2_reg2_reg_2_, p2_reg2_reg_3_, p2_reg2_reg_4_, p2_reg2_reg_5_,         p2_reg2_reg_6_, p2_reg2_reg_7_, p2_reg2_reg_8_, p2_reg2_reg_9_,         p2_reg2_reg_10_, p2_reg2_reg_11_, p2_reg2_reg_12_, p2_reg2_reg_13_,         p2_reg2_reg_14_, p2_reg2_reg_15_, p2_reg2_reg_16_, p2_reg2_reg_17_,         p2_reg2_reg_18_, p2_reg2_reg_19_, p2_reg2_reg_20_, p2_reg2_reg_21_,         p2_reg2_reg_22_, p2_reg2_reg_23_, p2_reg2_reg_24_, p2_reg2_reg_25_,         p2_reg2_reg_26_, p2_reg2_reg_27_, p2_reg2_reg_28_, p2_reg2_reg_29_,         p2_reg2_reg_30_, p2_reg2_reg_31_, p2_addr_reg_19_, p2_addr_reg_18_,         p2_addr_reg_17_, p2_addr_reg_16_, p2_addr_reg_15_, p2_addr_reg_14_,         p2_addr_reg_13_, p2_addr_reg_12_, p2_addr_reg_11_, p2_addr_reg_10_,         p2_addr_reg_9_, p2_addr_reg_8_, p2_addr_reg_7_, p2_addr_reg_6_,         p2_addr_reg_5_, p2_addr_reg_4_, p2_addr_reg_3_, p2_addr_reg_2_,         p2_addr_reg_1_, p2_addr_reg_0_, p2_datao_reg_0_, p2_datao_reg_1_,         p2_datao_reg_2_, p2_datao_reg_3_, p2_datao_reg_4_, p2_datao_reg_5_,         p2_datao_reg_6_, p2_datao_reg_7_, p2_datao_reg_8_, p2_datao_reg_9_,         p2_datao_reg_10_, p2_datao_reg_11_, p2_datao_reg_12_, p2_datao_reg_13_,         p2_datao_reg_14_, p2_datao_reg_15_, p2_datao_reg_16_, p2_datao_reg_17_,         p2_datao_reg_18_, p2_datao_reg_19_, p2_datao_reg_20_, p2_datao_reg_21_,         p2_datao_reg_22_, p2_datao_reg_23_, p2_datao_reg_24_, p2_datao_reg_25_,         p2_datao_reg_26_, p2_datao_reg_27_, p2_datao_reg_28_, p2_datao_reg_29_,         p2_datao_reg_30_, p2_datao_reg_31_, p2_b_reg, p2_reg3_reg_15_,         p2_reg3_reg_26_, p2_reg3_reg_6_, p2_reg3_reg_18_, p2_reg3_reg_2_,         p2_reg3_reg_11_, p2_reg3_reg_22_, p2_reg3_reg_13_, p2_reg3_reg_20_,         p2_reg3_reg_0_, p2_reg3_reg_9_, p2_reg3_reg_4_, p2_reg3_reg_24_,         p2_reg3_reg_17_, p2_reg3_reg_5_, p2_reg3_reg_16_, p2_reg3_reg_25_,         p2_reg3_reg_12_, p2_reg3_reg_21_, p2_reg3_reg_1_, p2_reg3_reg_8_,         p2_reg3_reg_28_, p2_reg3_reg_19_, p2_reg3_reg_3_, p2_reg3_reg_10_,         p2_reg3_reg_23_, p2_reg3_reg_14_, p2_reg3_reg_27_, p2_reg3_reg_7_,         p2_state_reg, p2_rd_reg, p2_wr_reg, p3_ir_reg_0_, p3_ir_reg_1_,         p3_ir_reg_2_, p3_ir_reg_3_, p3_ir_reg_4_, p3_ir_reg_5_, p3_ir_reg_6_,         p3_ir_reg_7_, p3_ir_reg_8_, p3_ir_reg_9_, p3_ir_reg_10_, p3_ir_reg_11_,         p3_ir_reg_12_, p3_ir_reg_13_, p3_ir_reg_14_, p3_ir_reg_15_,         p3_ir_reg_16_, p3_ir_reg_17_, p3_ir_reg_18_, p3_ir_reg_19_,         p3_ir_reg_20_, p3_ir_reg_21_, p3_ir_reg_22_, p3_ir_reg_23_,         p3_ir_reg_24_, p3_ir_reg_25_, p3_ir_reg_26_, p3_ir_reg_27_,         p3_ir_reg_28_, p3_ir_reg_29_, p3_ir_reg_30_, p3_ir_reg_31_,         p3_d_reg_0_, p3_d_reg_1_, p3_d_reg_2_, p3_d_reg_3_, p3_d_reg_4_,         p3_d_reg_5_, p3_d_reg_6_, p3_d_reg_7_, p3_d_reg_8_, p3_d_reg_9_,         p3_d_reg_10_, p3_d_reg_11_, p3_d_reg_12_, p3_d_reg_13_, p3_d_reg_14_,         p3_d_reg_15_, p3_d_reg_16_, p3_d_reg_17_, p3_d_reg_18_, p3_d_reg_19_,         p3_d_reg_20_, p3_d_reg_21_, p3_d_reg_22_, p3_d_reg_23_, p3_d_reg_24_,         p3_d_reg_25_, p3_d_reg_26_, p3_d_reg_27_, p3_d_reg_28_, p3_d_reg_29_,         p3_d_reg_30_, p3_d_reg_31_, p3_reg0_reg_0_, p3_reg0_reg_1_,         p3_reg0_reg_2_, p3_reg0_reg_3_, p3_reg0_reg_4_, p3_reg0_reg_5_,         p3_reg0_reg_6_, p3_reg0_reg_7_, p3_reg0_reg_8_, p3_reg0_reg_9_,         p3_reg0_reg_10_, p3_reg0_reg_11_, p3_reg0_reg_12_, p3_reg0_reg_13_,         p3_reg0_reg_14_, p3_reg0_reg_15_, p3_reg0_reg_16_, p3_reg0_reg_17_,         p3_reg0_reg_18_, p3_reg0_reg_19_, p3_reg0_reg_20_, p3_reg0_reg_21_,         p3_reg0_reg_22_, p3_reg0_reg_23_, p3_reg0_reg_24_, p3_reg0_reg_25_,         p3_reg0_reg_26_, p3_reg0_reg_27_, p3_reg0_reg_28_, p3_reg0_reg_29_,         p3_reg0_reg_30_, p3_reg0_reg_31_, p3_reg1_reg_0_, p3_reg1_reg_1_,         p3_reg1_reg_2_, p3_reg1_reg_3_, p3_reg1_reg_4_, p3_reg1_reg_5_,         p3_reg1_reg_6_, p3_reg1_reg_7_, p3_reg1_reg_8_, p3_reg1_reg_9_,         p3_reg1_reg_10_, p3_reg1_reg_11_, p3_reg1_reg_12_, p3_reg1_reg_13_,         p3_reg1_reg_14_, p3_reg1_reg_15_, p3_reg1_reg_16_, p3_reg1_reg_17_,         p3_reg1_reg_18_, p3_reg1_reg_19_, p3_reg1_reg_20_, p3_reg1_reg_21_,         p3_reg1_reg_22_, p3_reg1_reg_23_, p3_reg1_reg_24_, p3_reg1_reg_25_,         p3_reg1_reg_26_, p3_reg1_reg_27_, p3_reg1_reg_28_, p3_reg1_reg_29_,         p3_reg1_reg_30_, p3_reg1_reg_31_, p3_reg2_reg_0_, p3_reg2_reg_1_,         p3_reg2_reg_2_, p3_reg2_reg_3_, p3_reg2_reg_4_, p3_reg2_reg_5_,         p3_reg2_reg_6_, p3_reg2_reg_7_, p3_reg2_reg_8_, p3_reg2_reg_9_,         p3_reg2_reg_10_, p3_reg2_reg_11_, p3_reg2_reg_12_, p3_reg2_reg_13_,         p3_reg2_reg_14_, p3_reg2_reg_15_, p3_reg2_reg_16_, p3_reg2_reg_17_,         p3_reg2_reg_18_, p3_reg2_reg_19_, p3_reg2_reg_20_, p3_reg2_reg_21_,         p3_reg2_reg_22_, p3_reg2_reg_23_, p3_reg2_reg_24_, p3_reg2_reg_25_,         p3_reg2_reg_26_, p3_reg2_reg_27_, p3_reg2_reg_28_, p3_reg2_reg_29_,         p3_reg2_reg_30_, p3_reg2_reg_31_, p3_addr_reg_19_, p3_addr_reg_18_,         p3_addr_reg_17_, p3_addr_reg_16_, p3_addr_reg_15_, p3_addr_reg_14_,         p3_addr_reg_13_, p3_addr_reg_12_, p3_addr_reg_11_, p3_addr_reg_10_,         p3_addr_reg_9_, p3_addr_reg_8_, p3_addr_reg_7_, p3_addr_reg_6_,         p3_addr_reg_5_, p3_addr_reg_4_, p3_addr_reg_3_, p3_addr_reg_2_,         p3_addr_reg_1_, p3_addr_reg_0_, p3_datao_reg_0_, p3_datao_reg_1_,         p3_datao_reg_2_, p3_datao_reg_3_, p3_datao_reg_4_, p3_datao_reg_5_,         p3_datao_reg_6_, p3_datao_reg_7_, p3_datao_reg_8_, p3_datao_reg_9_,         p3_datao_reg_10_, p3_datao_reg_11_, p3_datao_reg_12_, p3_datao_reg_13_,         p3_datao_reg_14_, p3_datao_reg_15_, p3_datao_reg_16_, p3_datao_reg_17_,         p3_datao_reg_18_, p3_datao_reg_19_, p3_datao_reg_20_, p3_datao_reg_21_,         p3_datao_reg_22_, p3_datao_reg_23_, p3_datao_reg_24_, p3_datao_reg_25_,         p3_datao_reg_26_, p3_datao_reg_27_, p3_datao_reg_28_, p3_datao_reg_29_,         p3_datao_reg_30_, p3_datao_reg_31_, p3_b_reg, p3_reg3_reg_15_,         p3_reg3_reg_26_, p3_reg3_reg_6_, p3_reg3_reg_18_, p3_reg3_reg_2_,         p3_reg3_reg_11_, p3_reg3_reg_22_, p3_reg3_reg_13_, p3_reg3_reg_20_,         p3_reg3_reg_0_, p3_reg3_reg_9_, p3_reg3_reg_4_, p3_reg3_reg_24_,         p3_reg3_reg_17_, p3_reg3_reg_5_, p3_reg3_reg_16_, p3_reg3_reg_25_,         p3_reg3_reg_12_, p3_reg3_reg_21_, p3_reg3_reg_1_, p3_reg3_reg_8_,         p3_reg3_reg_28_, p3_reg3_reg_19_, p3_reg3_reg_3_, p3_reg3_reg_10_,         p3_reg3_reg_23_, p3_reg3_reg_14_, p3_reg3_reg_27_, p3_reg3_reg_7_,         p3_state_reg, p3_rd_reg, p3_wr_reg, sub_1596_u4, sub_1596_u62,         sub_1596_u63, sub_1596_u64, sub_1596_u65, sub_1596_u66, sub_1596_u67,         sub_1596_u68, sub_1596_u69, sub_1596_u70, sub_1596_u54, sub_1596_u55,         sub_1596_u56, sub_1596_u57, sub_1596_u58, sub_1596_u59, sub_1596_u60,         sub_1596_u61, sub_1596_u5, sub_1596_u53, u29, u28, p1_u3355, p1_u3354,         p1_u3353, p1_u3352, p1_u3351, p1_u3350, p1_u3349, p1_u3348, p1_u3347,         p1_u3346, p1_u3345, p1_u3344, p1_u3343, p1_u3342, p1_u3341, p1_u3340,         p1_u3339, p1_u3338, p1_u3337, p1_u3336, p1_u3335, p1_u3334, p1_u3333,         p1_u3332, p1_u3331, p1_u3330, p1_u3329, p1_u3328, p1_u3327, p1_u3326,         p1_u3325, p1_u3324, p1_u3445, p1_u3446, p1_u3323, p1_u3322, p1_u3321,         p1_u3320, p1_u3319, p1_u3318, p1_u3317, p1_u3316, p1_u3315, p1_u3314,         p1_u3313, p1_u3312, p1_u3311, p1_u3310, p1_u3309, p1_u3308, p1_u3307,         p1_u3306, p1_u3305, p1_u3304, p1_u3303, p1_u3302, p1_u3301, p1_u3300,         p1_u3299, p1_u3298, p1_u3297, p1_u3296, p1_u3295, p1_u3294, p1_u3459,         p1_u3462, p1_u3465, p1_u3468, p1_u3471, p1_u3474, p1_u3477, p1_u3480,         p1_u3483, p1_u3486, p1_u3489, p1_u3492, p1_u3495, p1_u3498, p1_u3501,         p1_u3504, p1_u3507, p1_u3510, p1_u3513, p1_u3515, p1_u3516, p1_u3517,         p1_u3518, p1_u3519, p1_u3520, p1_u3521, p1_u3522, p1_u3523, p1_u3524,         p1_u3525, p1_u3526, p1_u3527, p1_u3528, p1_u3529, p1_u3530, p1_u3531,         p1_u3532, p1_u3533, p1_u3534, p1_u3535, p1_u3536, p1_u3537, p1_u3538,         p1_u3539, p1_u3540, p1_u3541, p1_u3542, p1_u3543, p1_u3544, p1_u3545,         p1_u3546, p1_u3547, p1_u3548, p1_u3549, p1_u3550, p1_u3551, p1_u3552,         p1_u3553, p1_u3554, p1_u3555, p1_u3556, p1_u3557, p1_u3558, p1_u3559,         p1_u3293, p1_u3292, p1_u3291, p1_u3290, p1_u3289, p1_u3288, p1_u3287,         p1_u3286, p1_u3285, p1_u3284, p1_u3283, p1_u3282, p1_u3281, p1_u3280,         p1_u3279, p1_u3278, p1_u3277, p1_u3276, p1_u3275, p1_u3274, p1_u3273,         p1_u3272, p1_u3271, p1_u3270, p1_u3269, p1_u3268, p1_u3267, p1_u3266,         p1_u3265, p1_u3356, p1_u3264, p1_u3263, p1_u3262, p1_u3261, p1_u3260,         p1_u3259, p1_u3258, p1_u3257, p1_u3256, p1_u3255, p1_u3254, p1_u3253,         p1_u3252, p1_u3251, p1_u3250, p1_u3249, p1_u3248, p1_u3247, p1_u3246,         p1_u3245, p1_u3244, p1_u3243, p1_u3560, p1_u3561, p1_u3562, p1_u3563,         p1_u3564, p1_u3565, p1_u3566, p1_u3567, p1_u3568, p1_u3569, p1_u3570,         p1_u3571, p1_u3572, p1_u3573, p1_u3574, p1_u3575, p1_u3576, p1_u3577,         p1_u3578, p1_u3579, p1_u3580, p1_u3581, p1_u3582, p1_u3583, p1_u3584,         p1_u3585, p1_u3586, p1_u3587, p1_u3588, p1_u3589, p1_u3590, p1_u3591,         p1_u3242, p1_u3241, p1_u3240, p1_u3239, p1_u3238, p1_u3237, p1_u3236,         p1_u3235, p1_u3234, p1_u3233, p1_u3232, p1_u3231, p1_u3230, p1_u3229,         p1_u3228, p1_u3227, p1_u3226, p1_u3225, p1_u3224, p1_u3223, p1_u3222,         p1_u3221, p1_u3220, p1_u3219, p1_u3218, p1_u3217, p1_u3216, p1_u3215,         p1_u3214, p1_u3213, p1_u3086, p1_u3085, p1_u4016, p2_u3327, p2_u3326,         p2_u3325, p2_u3324, p2_u3323, p2_u3322, p2_u3321, p2_u3320, p2_u3319,         p2_u3318, p2_u3317, p2_u3316, p2_u3315, p2_u3314, p2_u3313, p2_u3312,         p2_u3311, p2_u3310, p2_u3309, p2_u3308, p2_u3307, p2_u3306, p2_u3305,         p2_u3304, p2_u3303, p2_u3302, p2_u3301, p2_u3300, p2_u3299, p2_u3298,         p2_u3297, p2_u3296, p2_u3416, p2_u3417, p2_u3295, p2_u3294, p2_u3293,         p2_u3292, p2_u3291, p2_u3290, p2_u3289, p2_u3288, p2_u3287, p2_u3286,         p2_u3285, p2_u3284, p2_u3283, p2_u3282, p2_u3281, p2_u3280, p2_u3279,         p2_u3278, p2_u3277, p2_u3276, p2_u3275, p2_u3274, p2_u3273, p2_u3272,         p2_u3271, p2_u3270, p2_u3269, p2_u3268, p2_u3267, p2_u3266, p2_u3430,         p2_u3433, p2_u3436, p2_u3439, p2_u3442, p2_u3445, p2_u3448, p2_u3451,         p2_u3454, p2_u3457, p2_u3460, p2_u3463, p2_u3466, p2_u3469, p2_u3472,         p2_u3475, p2_u3478, p2_u3481, p2_u3484, p2_u3486, p2_u3487, p2_u3488,         p2_u3489, p2_u3490, p2_u3491, p2_u3492, p2_u3493, p2_u3494, p2_u3495,         p2_u3496, p2_u3497, p2_u3498, p2_u3499, p2_u3500, p2_u3501, p2_u3502,         p2_u3503, p2_u3504, p2_u3505, p2_u3506, p2_u3507, p2_u3508, p2_u3509,         p2_u3510, p2_u3511, p2_u3512, p2_u3513, p2_u3514, p2_u3515, p2_u3516,         p2_u3517, p2_u3518, p2_u3519, p2_u3520, p2_u3521, p2_u3522, p2_u3523,         p2_u3524, p2_u3525, p2_u3526, p2_u3527, p2_u3528, p2_u3529, p2_u3530,         p2_u3265, p2_u3264, p2_u3263, p2_u3262, p2_u3261, p2_u3260, p2_u3259,         p2_u3258, p2_u3257, p2_u3256, p2_u3255, p2_u3254, p2_u3253, p2_u3252,         p2_u3251, p2_u3250, p2_u3249, p2_u3248, p2_u3247, p2_u3246, p2_u3245,         p2_u3244, p2_u3243, p2_u3242, p2_u3241, p2_u3240, p2_u3239, p2_u3238,         p2_u3237, p2_u3236, p2_u3235, p2_u3234, p2_u3233, p2_u3232, p2_u3231,         p2_u3230, p2_u3229, p2_u3228, p2_u3227, p2_u3226, p2_u3225, p2_u3224,         p2_u3223, p2_u3222, p2_u3221, p2_u3220, p2_u3219, p2_u3218, p2_u3217,         p2_u3216, p2_u3215, p2_u3214, p2_u3531, p2_u3532, p2_u3533, p2_u3534,         p2_u3535, p2_u3536, p2_u3537, p2_u3538, p2_u3539, p2_u3540, p2_u3541,         p2_u3542, p2_u3543, p2_u3544, p2_u3545, p2_u3546, p2_u3547, p2_u3548,         p2_u3549, p2_u3550, p2_u3551, p2_u3552, p2_u3553, p2_u3554, p2_u3555,         p2_u3556, p2_u3557, p2_u3558, p2_u3559, p2_u3560, p2_u3561, p2_u3562,         p2_u3328, p2_u3213, p2_u3212, p2_u3211, p2_u3210, p2_u3209, p2_u3208,         p2_u3207, p2_u3206, p2_u3205, p2_u3204, p2_u3203, p2_u3202, p2_u3201,         p2_u3200, p2_u3199, p2_u3198, p2_u3197, p2_u3196, p2_u3195, p2_u3194,         p2_u3193, p2_u3192, p2_u3191, p2_u3190, p2_u3189, p2_u3188, p2_u3187,         p2_u3186, p2_u3185, p2_u3088, p2_u3087, p2_u3947, p3_u3295, p3_u3294,         p3_u3293, p3_u3292, p3_u3291, p3_u3290, p3_u3289, p3_u3288, p3_u3287,         p3_u3286, p3_u3285, p3_u3284, p3_u3283, p3_u3282, p3_u3281, p3_u3280,         p3_u3279, p3_u3278, p3_u3277, p3_u3276, p3_u3275, p3_u3274, p3_u3273,         p3_u3272, p3_u3271, p3_u3270, p3_u3269, p3_u3268, p3_u3267, p3_u3266,         p3_u3265, p3_u3264, p3_u3376, p3_u3377, p3_u3263, p3_u3262, p3_u3261,         p3_u3260, p3_u3259, p3_u3258, p3_u3257, p3_u3256, p3_u3255, p3_u3254,         p3_u3253, p3_u3252, p3_u3251, p3_u3250, p3_u3249, p3_u3248, p3_u3247,         p3_u3246, p3_u3245, p3_u3244, p3_u3243, p3_u3242, p3_u3241, p3_u3240,         p3_u3239, p3_u3238, p3_u3237, p3_u3236, p3_u3235, p3_u3234, p3_u3390,         p3_u3393, p3_u3396, p3_u3399, p3_u3402, p3_u3405, p3_u3408, p3_u3411,         p3_u3414, p3_u3417, p3_u3420, p3_u3423, p3_u3426, p3_u3429, p3_u3432,         p3_u3435, p3_u3438, p3_u3441, p3_u3444, p3_u3446, p3_u3447, p3_u3448,         p3_u3449, p3_u3450, p3_u3451, p3_u3452, p3_u3453, p3_u3454, p3_u3455,         p3_u3456, p3_u3457, p3_u3458, p3_u3459, p3_u3460, p3_u3461, p3_u3462,         p3_u3463, p3_u3464, p3_u3465, p3_u3466, p3_u3467, p3_u3468, p3_u3469,         p3_u3470, p3_u3471, p3_u3472, p3_u3473, p3_u3474, p3_u3475, p3_u3476,         p3_u3477, p3_u3478, p3_u3479, p3_u3480, p3_u3481, p3_u3482, p3_u3483,         p3_u3484, p3_u3485, p3_u3486, p3_u3487, p3_u3488, p3_u3489, p3_u3490,         p3_u3233, p3_u3232, p3_u3231, p3_u3230, p3_u3229, p3_u3228, p3_u3227,         p3_u3226, p3_u3225, p3_u3224, p3_u3223, p3_u3222, p3_u3221, p3_u3220,         p3_u3219, p3_u3218, p3_u3217, p3_u3216, p3_u3215, p3_u3214, p3_u3213,         p3_u3212, p3_u3211, p3_u3210, p3_u3209, p3_u3208, p3_u3207, p3_u3206,         p3_u3205, p3_u3204, p3_u3203, p3_u3202, p3_u3201, p3_u3200, p3_u3199,         p3_u3198, p3_u3197, p3_u3196, p3_u3195, p3_u3194, p3_u3193, p3_u3192,         p3_u3191, p3_u3190, p3_u3189, p3_u3188, p3_u3187, p3_u3186, p3_u3185,         p3_u3184, p3_u3183, p3_u3182, p3_u3491, p3_u3492, p3_u3493, p3_u3494,         p3_u3495, p3_u3496, p3_u3497, p3_u3498, p3_u3499, p3_u3500, p3_u3501,         p3_u3502, p3_u3503, p3_u3504, p3_u3505, p3_u3506, p3_u3507, p3_u3508,         p3_u3509, p3_u3510, p3_u3511, p3_u3512, p3_u3513, p3_u3514, p3_u3515,         p3_u3516, p3_u3517, p3_u3518, p3_u3519, p3_u3520, p3_u3521, p3_u3522,         p3_u3296, p3_u3181, p3_u3180, p3_u3179, p3_u3178, p3_u3177, p3_u3176,         p3_u3175, p3_u3174, p3_u3173, p3_u3172, p3_u3171, p3_u3170, p3_u3169,         p3_u3168, p3_u3167, p3_u3166, p3_u3165, p3_u3164, p3_u3163, p3_u3162,         p3_u3161, p3_u3160, p3_u3159, p3_u3158, p3_u3157, p3_u3156, p3_u3155,         p3_u3154, p3_u3153, p3_u3151, p3_u3150, p3_u3897 );
input si_31_, si_30_, si_29_, si_28_, si_27_, si_26_, si_25_, si_24_, si_23_,         si_22_, si_21_, si_20_, si_19_, si_18_, si_17_, si_16_, si_15_,         si_14_, si_13_, si_12_, si_11_, si_10_, si_9_, si_8_, si_7_, si_6_,         si_5_, si_4_, si_3_, si_2_, si_1_, si_0_, p1_ir_reg_0_, p1_ir_reg_1_,         p1_ir_reg_2_, p1_ir_reg_3_, p1_ir_reg_4_, p1_ir_reg_5_, p1_ir_reg_6_,         p1_ir_reg_7_, p1_ir_reg_8_, p1_ir_reg_9_, p1_ir_reg_10_,         p1_ir_reg_11_, p1_ir_reg_12_, p1_ir_reg_13_, p1_ir_reg_14_,         p1_ir_reg_15_, p1_ir_reg_16_, p1_ir_reg_17_, p1_ir_reg_18_,         p1_ir_reg_19_, p1_ir_reg_20_, p1_ir_reg_21_, p1_ir_reg_22_,         p1_ir_reg_23_, p1_ir_reg_24_, p1_ir_reg_25_, p1_ir_reg_26_,         p1_ir_reg_27_, p1_ir_reg_28_, p1_ir_reg_29_, p1_ir_reg_30_,         p1_ir_reg_31_, p1_d_reg_0_, p1_d_reg_1_, p1_d_reg_2_, p1_d_reg_3_,         p1_d_reg_4_, p1_d_reg_5_, p1_d_reg_6_, p1_d_reg_7_, p1_d_reg_8_,         p1_d_reg_9_, p1_d_reg_10_, p1_d_reg_11_, p1_d_reg_12_, p1_d_reg_13_,         p1_d_reg_14_, p1_d_reg_15_, p1_d_reg_16_, p1_d_reg_17_, p1_d_reg_18_,         p1_d_reg_19_, p1_d_reg_20_, p1_d_reg_21_, p1_d_reg_22_, p1_d_reg_23_,         p1_d_reg_24_, p1_d_reg_25_, p1_d_reg_26_, p1_d_reg_27_, p1_d_reg_28_,         p1_d_reg_29_, p1_d_reg_30_, p1_d_reg_31_, p1_reg0_reg_0_,         p1_reg0_reg_1_, p1_reg0_reg_2_, p1_reg0_reg_3_, p1_reg0_reg_4_,         p1_reg0_reg_5_, p1_reg0_reg_6_, p1_reg0_reg_7_, p1_reg0_reg_8_,         p1_reg0_reg_9_, p1_reg0_reg_10_, p1_reg0_reg_11_, p1_reg0_reg_12_,         p1_reg0_reg_13_, p1_reg0_reg_14_, p1_reg0_reg_15_, p1_reg0_reg_16_,         p1_reg0_reg_17_, p1_reg0_reg_18_, p1_reg0_reg_19_, p1_reg0_reg_20_,         p1_reg0_reg_21_, p1_reg0_reg_22_, p1_reg0_reg_23_, p1_reg0_reg_24_,         p1_reg0_reg_25_, p1_reg0_reg_26_, p1_reg0_reg_27_, p1_reg0_reg_28_,         p1_reg0_reg_29_, p1_reg0_reg_30_, p1_reg0_reg_31_, p1_reg1_reg_0_,         p1_reg1_reg_1_, p1_reg1_reg_2_, p1_reg1_reg_3_, p1_reg1_reg_4_,         p1_reg1_reg_5_, p1_reg1_reg_6_, p1_reg1_reg_7_, p1_reg1_reg_8_,         p1_reg1_reg_9_, p1_reg1_reg_10_, p1_reg1_reg_11_, p1_reg1_reg_12_,         p1_reg1_reg_13_, p1_reg1_reg_14_, p1_reg1_reg_15_, p1_reg1_reg_16_,         p1_reg1_reg_17_, p1_reg1_reg_18_, p1_reg1_reg_19_, p1_reg1_reg_20_,         p1_reg1_reg_21_, p1_reg1_reg_22_, p1_reg1_reg_23_, p1_reg1_reg_24_,         p1_reg1_reg_25_, p1_reg1_reg_26_, p1_reg1_reg_27_, p1_reg1_reg_28_,         p1_reg1_reg_29_, p1_reg1_reg_30_, p1_reg1_reg_31_, p1_reg2_reg_0_,         p1_reg2_reg_1_, p1_reg2_reg_2_, p1_reg2_reg_3_, p1_reg2_reg_4_,         p1_reg2_reg_5_, p1_reg2_reg_6_, p1_reg2_reg_7_, p1_reg2_reg_8_,         p1_reg2_reg_9_, p1_reg2_reg_10_, p1_reg2_reg_11_, p1_reg2_reg_12_,         p1_reg2_reg_13_, p1_reg2_reg_14_, p1_reg2_reg_15_, p1_reg2_reg_16_,         p1_reg2_reg_17_, p1_reg2_reg_18_, p1_reg2_reg_19_, p1_reg2_reg_20_,         p1_reg2_reg_21_, p1_reg2_reg_22_, p1_reg2_reg_23_, p1_reg2_reg_24_,         p1_reg2_reg_25_, p1_reg2_reg_26_, p1_reg2_reg_27_, p1_reg2_reg_28_,         p1_reg2_reg_29_, p1_reg2_reg_30_, p1_reg2_reg_31_, p1_addr_reg_19_,         p1_addr_reg_18_, p1_addr_reg_17_, p1_addr_reg_16_, p1_addr_reg_15_,         p1_addr_reg_14_, p1_addr_reg_13_, p1_addr_reg_12_, p1_addr_reg_11_,         p1_addr_reg_10_, p1_addr_reg_9_, p1_addr_reg_8_, p1_addr_reg_7_,         p1_addr_reg_6_, p1_addr_reg_5_, p1_addr_reg_4_, p1_addr_reg_3_,         p1_addr_reg_2_, p1_addr_reg_1_, p1_addr_reg_0_, p1_datao_reg_0_,         p1_datao_reg_1_, p1_datao_reg_2_, p1_datao_reg_3_, p1_datao_reg_4_,         p1_datao_reg_5_, p1_datao_reg_6_, p1_datao_reg_7_, p1_datao_reg_8_,         p1_datao_reg_9_, p1_datao_reg_10_, p1_datao_reg_11_, p1_datao_reg_12_,         p1_datao_reg_13_, p1_datao_reg_14_, p1_datao_reg_15_,         p1_datao_reg_16_, p1_datao_reg_17_, p1_datao_reg_18_,         p1_datao_reg_19_, p1_datao_reg_20_, p1_datao_reg_21_,         p1_datao_reg_22_, p1_datao_reg_23_, p1_datao_reg_24_,         p1_datao_reg_25_, p1_datao_reg_26_, p1_datao_reg_27_,         p1_datao_reg_28_, p1_datao_reg_29_, p1_datao_reg_30_,         p1_datao_reg_31_, p1_b_reg, p1_reg3_reg_15_, p1_reg3_reg_26_,         p1_reg3_reg_6_, p1_reg3_reg_18_, p1_reg3_reg_2_, p1_reg3_reg_11_,         p1_reg3_reg_22_, p1_reg3_reg_13_, p1_reg3_reg_20_, p1_reg3_reg_0_,         p1_reg3_reg_9_, p1_reg3_reg_4_, p1_reg3_reg_24_, p1_reg3_reg_17_,         p1_reg3_reg_5_, p1_reg3_reg_16_, p1_reg3_reg_25_, p1_reg3_reg_12_,         p1_reg3_reg_21_, p1_reg3_reg_1_, p1_reg3_reg_8_, p1_reg3_reg_28_,         p1_reg3_reg_19_, p1_reg3_reg_3_, p1_reg3_reg_10_, p1_reg3_reg_23_,         p1_reg3_reg_14_, p1_reg3_reg_27_, p1_reg3_reg_7_, p1_state_reg,         p1_rd_reg, p1_wr_reg, p2_ir_reg_0_, p2_ir_reg_1_, p2_ir_reg_2_,         p2_ir_reg_3_, p2_ir_reg_4_, p2_ir_reg_5_, p2_ir_reg_6_, p2_ir_reg_7_,         p2_ir_reg_8_, p2_ir_reg_9_, p2_ir_reg_10_, p2_ir_reg_11_,         p2_ir_reg_12_, p2_ir_reg_13_, p2_ir_reg_14_, p2_ir_reg_15_,         p2_ir_reg_16_, p2_ir_reg_17_, p2_ir_reg_18_, p2_ir_reg_19_,         p2_ir_reg_20_, p2_ir_reg_21_, p2_ir_reg_22_, p2_ir_reg_23_,         p2_ir_reg_24_, p2_ir_reg_25_, p2_ir_reg_26_, p2_ir_reg_27_,         p2_ir_reg_28_, p2_ir_reg_29_, p2_ir_reg_30_, p2_ir_reg_31_,         p2_d_reg_0_, p2_d_reg_1_, p2_d_reg_2_, p2_d_reg_3_, p2_d_reg_4_,         p2_d_reg_5_, p2_d_reg_6_, p2_d_reg_7_, p2_d_reg_8_, p2_d_reg_9_,         p2_d_reg_10_, p2_d_reg_11_, p2_d_reg_12_, p2_d_reg_13_, p2_d_reg_14_,         p2_d_reg_15_, p2_d_reg_16_, p2_d_reg_17_, p2_d_reg_18_, p2_d_reg_19_,         p2_d_reg_20_, p2_d_reg_21_, p2_d_reg_22_, p2_d_reg_23_, p2_d_reg_24_,         p2_d_reg_25_, p2_d_reg_26_, p2_d_reg_27_, p2_d_reg_28_, p2_d_reg_29_,         p2_d_reg_30_, p2_d_reg_31_, p2_reg0_reg_0_, p2_reg0_reg_1_,         p2_reg0_reg_2_, p2_reg0_reg_3_, p2_reg0_reg_4_, p2_reg0_reg_5_,         p2_reg0_reg_6_, p2_reg0_reg_7_, p2_reg0_reg_8_, p2_reg0_reg_9_,         p2_reg0_reg_10_, p2_reg0_reg_11_, p2_reg0_reg_12_, p2_reg0_reg_13_,         p2_reg0_reg_14_, p2_reg0_reg_15_, p2_reg0_reg_16_, p2_reg0_reg_17_,         p2_reg0_reg_18_, p2_reg0_reg_19_, p2_reg0_reg_20_, p2_reg0_reg_21_,         p2_reg0_reg_22_, p2_reg0_reg_23_, p2_reg0_reg_24_, p2_reg0_reg_25_,         p2_reg0_reg_26_, p2_reg0_reg_27_, p2_reg0_reg_28_, p2_reg0_reg_29_,         p2_reg0_reg_30_, p2_reg0_reg_31_, p2_reg1_reg_0_, p2_reg1_reg_1_,         p2_reg1_reg_2_, p2_reg1_reg_3_, p2_reg1_reg_4_, p2_reg1_reg_5_,         p2_reg1_reg_6_, p2_reg1_reg_7_, p2_reg1_reg_8_, p2_reg1_reg_9_,         p2_reg1_reg_10_, p2_reg1_reg_11_, p2_reg1_reg_12_, p2_reg1_reg_13_,         p2_reg1_reg_14_, p2_reg1_reg_15_, p2_reg1_reg_16_, p2_reg1_reg_17_,         p2_reg1_reg_18_, p2_reg1_reg_19_, p2_reg1_reg_20_, p2_reg1_reg_21_,         p2_reg1_reg_22_, p2_reg1_reg_23_, p2_reg1_reg_24_, p2_reg1_reg_25_,         p2_reg1_reg_26_, p2_reg1_reg_27_, p2_reg1_reg_28_, p2_reg1_reg_29_,         p2_reg1_reg_30_, p2_reg1_reg_31_, p2_reg2_reg_0_, p2_reg2_reg_1_,         p2_reg2_reg_2_, p2_reg2_reg_3_, p2_reg2_reg_4_, p2_reg2_reg_5_,         p2_reg2_reg_6_, p2_reg2_reg_7_, p2_reg2_reg_8_, p2_reg2_reg_9_,         p2_reg2_reg_10_, p2_reg2_reg_11_, p2_reg2_reg_12_, p2_reg2_reg_13_,         p2_reg2_reg_14_, p2_reg2_reg_15_, p2_reg2_reg_16_, p2_reg2_reg_17_,         p2_reg2_reg_18_, p2_reg2_reg_19_, p2_reg2_reg_20_, p2_reg2_reg_21_,         p2_reg2_reg_22_, p2_reg2_reg_23_, p2_reg2_reg_24_, p2_reg2_reg_25_,         p2_reg2_reg_26_, p2_reg2_reg_27_, p2_reg2_reg_28_, p2_reg2_reg_29_,         p2_reg2_reg_30_, p2_reg2_reg_31_, p2_addr_reg_19_, p2_addr_reg_18_,         p2_addr_reg_17_, p2_addr_reg_16_, p2_addr_reg_15_, p2_addr_reg_14_,         p2_addr_reg_13_, p2_addr_reg_12_, p2_addr_reg_11_, p2_addr_reg_10_,         p2_addr_reg_9_, p2_addr_reg_8_, p2_addr_reg_7_, p2_addr_reg_6_,         p2_addr_reg_5_, p2_addr_reg_4_, p2_addr_reg_3_, p2_addr_reg_2_,         p2_addr_reg_1_, p2_addr_reg_0_, p2_datao_reg_0_, p2_datao_reg_1_,         p2_datao_reg_2_, p2_datao_reg_3_, p2_datao_reg_4_, p2_datao_reg_5_,         p2_datao_reg_6_, p2_datao_reg_7_, p2_datao_reg_8_, p2_datao_reg_9_,         p2_datao_reg_10_, p2_datao_reg_11_, p2_datao_reg_12_,         p2_datao_reg_13_, p2_datao_reg_14_, p2_datao_reg_15_,         p2_datao_reg_16_, p2_datao_reg_17_, p2_datao_reg_18_,         p2_datao_reg_19_, p2_datao_reg_20_, p2_datao_reg_21_,         p2_datao_reg_22_, p2_datao_reg_23_, p2_datao_reg_24_,         p2_datao_reg_25_, p2_datao_reg_26_, p2_datao_reg_27_,         p2_datao_reg_28_, p2_datao_reg_29_, p2_datao_reg_30_,         p2_datao_reg_31_, p2_b_reg, p2_reg3_reg_15_, p2_reg3_reg_26_,         p2_reg3_reg_6_, p2_reg3_reg_18_, p2_reg3_reg_2_, p2_reg3_reg_11_,         p2_reg3_reg_22_, p2_reg3_reg_13_, p2_reg3_reg_20_, p2_reg3_reg_0_,         p2_reg3_reg_9_, p2_reg3_reg_4_, p2_reg3_reg_24_, p2_reg3_reg_17_,         p2_reg3_reg_5_, p2_reg3_reg_16_, p2_reg3_reg_25_, p2_reg3_reg_12_,         p2_reg3_reg_21_, p2_reg3_reg_1_, p2_reg3_reg_8_, p2_reg3_reg_28_,         p2_reg3_reg_19_, p2_reg3_reg_3_, p2_reg3_reg_10_, p2_reg3_reg_23_,         p2_reg3_reg_14_, p2_reg3_reg_27_, p2_reg3_reg_7_, p2_state_reg,         p2_rd_reg, p2_wr_reg, p3_ir_reg_0_, p3_ir_reg_1_, p3_ir_reg_2_,         p3_ir_reg_3_, p3_ir_reg_4_, p3_ir_reg_5_, p3_ir_reg_6_, p3_ir_reg_7_,         p3_ir_reg_8_, p3_ir_reg_9_, p3_ir_reg_10_, p3_ir_reg_11_,         p3_ir_reg_12_, p3_ir_reg_13_, p3_ir_reg_14_, p3_ir_reg_15_,         p3_ir_reg_16_, p3_ir_reg_17_, p3_ir_reg_18_, p3_ir_reg_19_,         p3_ir_reg_20_, p3_ir_reg_21_, p3_ir_reg_22_, p3_ir_reg_23_,         p3_ir_reg_24_, p3_ir_reg_25_, p3_ir_reg_26_, p3_ir_reg_27_,         p3_ir_reg_28_, p3_ir_reg_29_, p3_ir_reg_30_, p3_ir_reg_31_,         p3_d_reg_0_, p3_d_reg_1_, p3_d_reg_2_, p3_d_reg_3_, p3_d_reg_4_,         p3_d_reg_5_, p3_d_reg_6_, p3_d_reg_7_, p3_d_reg_8_, p3_d_reg_9_,         p3_d_reg_10_, p3_d_reg_11_, p3_d_reg_12_, p3_d_reg_13_, p3_d_reg_14_,         p3_d_reg_15_, p3_d_reg_16_, p3_d_reg_17_, p3_d_reg_18_, p3_d_reg_19_,         p3_d_reg_20_, p3_d_reg_21_, p3_d_reg_22_, p3_d_reg_23_, p3_d_reg_24_,         p3_d_reg_25_, p3_d_reg_26_, p3_d_reg_27_, p3_d_reg_28_, p3_d_reg_29_,         p3_d_reg_30_, p3_d_reg_31_, p3_reg0_reg_0_, p3_reg0_reg_1_,         p3_reg0_reg_2_, p3_reg0_reg_3_, p3_reg0_reg_4_, p3_reg0_reg_5_,         p3_reg0_reg_6_, p3_reg0_reg_7_, p3_reg0_reg_8_, p3_reg0_reg_9_,         p3_reg0_reg_10_, p3_reg0_reg_11_, p3_reg0_reg_12_, p3_reg0_reg_13_,         p3_reg0_reg_14_, p3_reg0_reg_15_, p3_reg0_reg_16_, p3_reg0_reg_17_,         p3_reg0_reg_18_, p3_reg0_reg_19_, p3_reg0_reg_20_, p3_reg0_reg_21_,         p3_reg0_reg_22_, p3_reg0_reg_23_, p3_reg0_reg_24_, p3_reg0_reg_25_,         p3_reg0_reg_26_, p3_reg0_reg_27_, p3_reg0_reg_28_, p3_reg0_reg_29_,         p3_reg0_reg_30_, p3_reg0_reg_31_, p3_reg1_reg_0_, p3_reg1_reg_1_,         p3_reg1_reg_2_, p3_reg1_reg_3_, p3_reg1_reg_4_, p3_reg1_reg_5_,         p3_reg1_reg_6_, p3_reg1_reg_7_, p3_reg1_reg_8_, p3_reg1_reg_9_,         p3_reg1_reg_10_, p3_reg1_reg_11_, p3_reg1_reg_12_, p3_reg1_reg_13_,         p3_reg1_reg_14_, p3_reg1_reg_15_, p3_reg1_reg_16_, p3_reg1_reg_17_,         p3_reg1_reg_18_, p3_reg1_reg_19_, p3_reg1_reg_20_, p3_reg1_reg_21_,         p3_reg1_reg_22_, p3_reg1_reg_23_, p3_reg1_reg_24_, p3_reg1_reg_25_,         p3_reg1_reg_26_, p3_reg1_reg_27_, p3_reg1_reg_28_, p3_reg1_reg_29_,         p3_reg1_reg_30_, p3_reg1_reg_31_, p3_reg2_reg_0_, p3_reg2_reg_1_,         p3_reg2_reg_2_, p3_reg2_reg_3_, p3_reg2_reg_4_, p3_reg2_reg_5_,         p3_reg2_reg_6_, p3_reg2_reg_7_, p3_reg2_reg_8_, p3_reg2_reg_9_,         p3_reg2_reg_10_, p3_reg2_reg_11_, p3_reg2_reg_12_, p3_reg2_reg_13_,         p3_reg2_reg_14_, p3_reg2_reg_15_, p3_reg2_reg_16_, p3_reg2_reg_17_,         p3_reg2_reg_18_, p3_reg2_reg_19_, p3_reg2_reg_20_, p3_reg2_reg_21_,         p3_reg2_reg_22_, p3_reg2_reg_23_, p3_reg2_reg_24_, p3_reg2_reg_25_,         p3_reg2_reg_26_, p3_reg2_reg_27_, p3_reg2_reg_28_, p3_reg2_reg_29_,         p3_reg2_reg_30_, p3_reg2_reg_31_, p3_addr_reg_19_, p3_addr_reg_18_,         p3_addr_reg_17_, p3_addr_reg_16_, p3_addr_reg_15_, p3_addr_reg_14_,         p3_addr_reg_13_, p3_addr_reg_12_, p3_addr_reg_11_, p3_addr_reg_10_,         p3_addr_reg_9_, p3_addr_reg_8_, p3_addr_reg_7_, p3_addr_reg_6_,         p3_addr_reg_5_, p3_addr_reg_4_, p3_addr_reg_3_, p3_addr_reg_2_,         p3_addr_reg_1_, p3_addr_reg_0_, p3_datao_reg_0_, p3_datao_reg_1_,         p3_datao_reg_2_, p3_datao_reg_3_, p3_datao_reg_4_, p3_datao_reg_5_,         p3_datao_reg_6_, p3_datao_reg_7_, p3_datao_reg_8_, p3_datao_reg_9_,         p3_datao_reg_10_, p3_datao_reg_11_, p3_datao_reg_12_,         p3_datao_reg_13_, p3_datao_reg_14_, p3_datao_reg_15_,         p3_datao_reg_16_, p3_datao_reg_17_, p3_datao_reg_18_,         p3_datao_reg_19_, p3_datao_reg_20_, p3_datao_reg_21_,         p3_datao_reg_22_, p3_datao_reg_23_, p3_datao_reg_24_,         p3_datao_reg_25_, p3_datao_reg_26_, p3_datao_reg_27_,         p3_datao_reg_28_, p3_datao_reg_29_, p3_datao_reg_30_,         p3_datao_reg_31_, p3_b_reg, p3_reg3_reg_15_, p3_reg3_reg_26_,         p3_reg3_reg_6_, p3_reg3_reg_18_, p3_reg3_reg_2_, p3_reg3_reg_11_,         p3_reg3_reg_22_, p3_reg3_reg_13_, p3_reg3_reg_20_, p3_reg3_reg_0_,         p3_reg3_reg_9_, p3_reg3_reg_4_, p3_reg3_reg_24_, p3_reg3_reg_17_,         p3_reg3_reg_5_, p3_reg3_reg_16_, p3_reg3_reg_25_, p3_reg3_reg_12_,         p3_reg3_reg_21_, p3_reg3_reg_1_, p3_reg3_reg_8_, p3_reg3_reg_28_,         p3_reg3_reg_19_, p3_reg3_reg_3_, p3_reg3_reg_10_, p3_reg3_reg_23_,         p3_reg3_reg_14_, p3_reg3_reg_27_, p3_reg3_reg_7_, p3_state_reg,         p3_rd_reg, p3_wr_reg;
output sub_1596_u4, sub_1596_u62, sub_1596_u63, sub_1596_u64, sub_1596_u65,         sub_1596_u66, sub_1596_u67, sub_1596_u68, sub_1596_u69, sub_1596_u70,         sub_1596_u54, sub_1596_u55, sub_1596_u56, sub_1596_u57, sub_1596_u58,         sub_1596_u59, sub_1596_u60, sub_1596_u61, sub_1596_u5, sub_1596_u53,         u29, u28, p1_u3355, p1_u3354, p1_u3353, p1_u3352, p1_u3351, p1_u3350,         p1_u3349, p1_u3348, p1_u3347, p1_u3346, p1_u3345, p1_u3344, p1_u3343,         p1_u3342, p1_u3341, p1_u3340, p1_u3339, p1_u3338, p1_u3337, p1_u3336,         p1_u3335, p1_u3334, p1_u3333, p1_u3332, p1_u3331, p1_u3330, p1_u3329,         p1_u3328, p1_u3327, p1_u3326, p1_u3325, p1_u3324, p1_u3445, p1_u3446,         p1_u3323, p1_u3322, p1_u3321, p1_u3320, p1_u3319, p1_u3318, p1_u3317,         p1_u3316, p1_u3315, p1_u3314, p1_u3313, p1_u3312, p1_u3311, p1_u3310,         p1_u3309, p1_u3308, p1_u3307, p1_u3306, p1_u3305, p1_u3304, p1_u3303,         p1_u3302, p1_u3301, p1_u3300, p1_u3299, p1_u3298, p1_u3297, p1_u3296,         p1_u3295, p1_u3294, p1_u3459, p1_u3462, p1_u3465, p1_u3468, p1_u3471,         p1_u3474, p1_u3477, p1_u3480, p1_u3483, p1_u3486, p1_u3489, p1_u3492,         p1_u3495, p1_u3498, p1_u3501, p1_u3504, p1_u3507, p1_u3510, p1_u3513,         p1_u3515, p1_u3516, p1_u3517, p1_u3518, p1_u3519, p1_u3520, p1_u3521,         p1_u3522, p1_u3523, p1_u3524, p1_u3525, p1_u3526, p1_u3527, p1_u3528,         p1_u3529, p1_u3530, p1_u3531, p1_u3532, p1_u3533, p1_u3534, p1_u3535,         p1_u3536, p1_u3537, p1_u3538, p1_u3539, p1_u3540, p1_u3541, p1_u3542,         p1_u3543, p1_u3544, p1_u3545, p1_u3546, p1_u3547, p1_u3548, p1_u3549,         p1_u3550, p1_u3551, p1_u3552, p1_u3553, p1_u3554, p1_u3555, p1_u3556,         p1_u3557, p1_u3558, p1_u3559, p1_u3293, p1_u3292, p1_u3291, p1_u3290,         p1_u3289, p1_u3288, p1_u3287, p1_u3286, p1_u3285, p1_u3284, p1_u3283,         p1_u3282, p1_u3281, p1_u3280, p1_u3279, p1_u3278, p1_u3277, p1_u3276,         p1_u3275, p1_u3274, p1_u3273, p1_u3272, p1_u3271, p1_u3270, p1_u3269,         p1_u3268, p1_u3267, p1_u3266, p1_u3265, p1_u3356, p1_u3264, p1_u3263,         p1_u3262, p1_u3261, p1_u3260, p1_u3259, p1_u3258, p1_u3257, p1_u3256,         p1_u3255, p1_u3254, p1_u3253, p1_u3252, p1_u3251, p1_u3250, p1_u3249,         p1_u3248, p1_u3247, p1_u3246, p1_u3245, p1_u3244, p1_u3243, p1_u3560,         p1_u3561, p1_u3562, p1_u3563, p1_u3564, p1_u3565, p1_u3566, p1_u3567,         p1_u3568, p1_u3569, p1_u3570, p1_u3571, p1_u3572, p1_u3573, p1_u3574,         p1_u3575, p1_u3576, p1_u3577, p1_u3578, p1_u3579, p1_u3580, p1_u3581,         p1_u3582, p1_u3583, p1_u3584, p1_u3585, p1_u3586, p1_u3587, p1_u3588,         p1_u3589, p1_u3590, p1_u3591, p1_u3242, p1_u3241, p1_u3240, p1_u3239,         p1_u3238, p1_u3237, p1_u3236, p1_u3235, p1_u3234, p1_u3233, p1_u3232,         p1_u3231, p1_u3230, p1_u3229, p1_u3228, p1_u3227, p1_u3226, p1_u3225,         p1_u3224, p1_u3223, p1_u3222, p1_u3221, p1_u3220, p1_u3219, p1_u3218,         p1_u3217, p1_u3216, p1_u3215, p1_u3214, p1_u3213, p1_u3086, p1_u3085,         p1_u4016, p2_u3327, p2_u3326, p2_u3325, p2_u3324, p2_u3323, p2_u3322,         p2_u3321, p2_u3320, p2_u3319, p2_u3318, p2_u3317, p2_u3316, p2_u3315,         p2_u3314, p2_u3313, p2_u3312, p2_u3311, p2_u3310, p2_u3309, p2_u3308,         p2_u3307, p2_u3306, p2_u3305, p2_u3304, p2_u3303, p2_u3302, p2_u3301,         p2_u3300, p2_u3299, p2_u3298, p2_u3297, p2_u3296, p2_u3416, p2_u3417,         p2_u3295, p2_u3294, p2_u3293, p2_u3292, p2_u3291, p2_u3290, p2_u3289,         p2_u3288, p2_u3287, p2_u3286, p2_u3285, p2_u3284, p2_u3283, p2_u3282,         p2_u3281, p2_u3280, p2_u3279, p2_u3278, p2_u3277, p2_u3276, p2_u3275,         p2_u3274, p2_u3273, p2_u3272, p2_u3271, p2_u3270, p2_u3269, p2_u3268,         p2_u3267, p2_u3266, p2_u3430, p2_u3433, p2_u3436, p2_u3439, p2_u3442,         p2_u3445, p2_u3448, p2_u3451, p2_u3454, p2_u3457, p2_u3460, p2_u3463,         p2_u3466, p2_u3469, p2_u3472, p2_u3475, p2_u3478, p2_u3481, p2_u3484,         p2_u3486, p2_u3487, p2_u3488, p2_u3489, p2_u3490, p2_u3491, p2_u3492,         p2_u3493, p2_u3494, p2_u3495, p2_u3496, p2_u3497, p2_u3498, p2_u3499,         p2_u3500, p2_u3501, p2_u3502, p2_u3503, p2_u3504, p2_u3505, p2_u3506,         p2_u3507, p2_u3508, p2_u3509, p2_u3510, p2_u3511, p2_u3512, p2_u3513,         p2_u3514, p2_u3515, p2_u3516, p2_u3517, p2_u3518, p2_u3519, p2_u3520,         p2_u3521, p2_u3522, p2_u3523, p2_u3524, p2_u3525, p2_u3526, p2_u3527,         p2_u3528, p2_u3529, p2_u3530, p2_u3265, p2_u3264, p2_u3263, p2_u3262,         p2_u3261, p2_u3260, p2_u3259, p2_u3258, p2_u3257, p2_u3256, p2_u3255,         p2_u3254, p2_u3253, p2_u3252, p2_u3251, p2_u3250, p2_u3249, p2_u3248,         p2_u3247, p2_u3246, p2_u3245, p2_u3244, p2_u3243, p2_u3242, p2_u3241,         p2_u3240, p2_u3239, p2_u3238, p2_u3237, p2_u3236, p2_u3235, p2_u3234,         p2_u3233, p2_u3232, p2_u3231, p2_u3230, p2_u3229, p2_u3228, p2_u3227,         p2_u3226, p2_u3225, p2_u3224, p2_u3223, p2_u3222, p2_u3221, p2_u3220,         p2_u3219, p2_u3218, p2_u3217, p2_u3216, p2_u3215, p2_u3214, p2_u3531,         p2_u3532, p2_u3533, p2_u3534, p2_u3535, p2_u3536, p2_u3537, p2_u3538,         p2_u3539, p2_u3540, p2_u3541, p2_u3542, p2_u3543, p2_u3544, p2_u3545,         p2_u3546, p2_u3547, p2_u3548, p2_u3549, p2_u3550, p2_u3551, p2_u3552,         p2_u3553, p2_u3554, p2_u3555, p2_u3556, p2_u3557, p2_u3558, p2_u3559,         p2_u3560, p2_u3561, p2_u3562, p2_u3328, p2_u3213, p2_u3212, p2_u3211,         p2_u3210, p2_u3209, p2_u3208, p2_u3207, p2_u3206, p2_u3205, p2_u3204,         p2_u3203, p2_u3202, p2_u3201, p2_u3200, p2_u3199, p2_u3198, p2_u3197,         p2_u3196, p2_u3195, p2_u3194, p2_u3193, p2_u3192, p2_u3191, p2_u3190,         p2_u3189, p2_u3188, p2_u3187, p2_u3186, p2_u3185, p2_u3088, p2_u3087,         p2_u3947, p3_u3295, p3_u3294, p3_u3293, p3_u3292, p3_u3291, p3_u3290,         p3_u3289, p3_u3288, p3_u3287, p3_u3286, p3_u3285, p3_u3284, p3_u3283,         p3_u3282, p3_u3281, p3_u3280, p3_u3279, p3_u3278, p3_u3277, p3_u3276,         p3_u3275, p3_u3274, p3_u3273, p3_u3272, p3_u3271, p3_u3270, p3_u3269,         p3_u3268, p3_u3267, p3_u3266, p3_u3265, p3_u3264, p3_u3376, p3_u3377,         p3_u3263, p3_u3262, p3_u3261, p3_u3260, p3_u3259, p3_u3258, p3_u3257,         p3_u3256, p3_u3255, p3_u3254, p3_u3253, p3_u3252, p3_u3251, p3_u3250,         p3_u3249, p3_u3248, p3_u3247, p3_u3246, p3_u3245, p3_u3244, p3_u3243,         p3_u3242, p3_u3241, p3_u3240, p3_u3239, p3_u3238, p3_u3237, p3_u3236,         p3_u3235, p3_u3234, p3_u3390, p3_u3393, p3_u3396, p3_u3399, p3_u3402,         p3_u3405, p3_u3408, p3_u3411, p3_u3414, p3_u3417, p3_u3420, p3_u3423,         p3_u3426, p3_u3429, p3_u3432, p3_u3435, p3_u3438, p3_u3441, p3_u3444,         p3_u3446, p3_u3447, p3_u3448, p3_u3449, p3_u3450, p3_u3451, p3_u3452,         p3_u3453, p3_u3454, p3_u3455, p3_u3456, p3_u3457, p3_u3458, p3_u3459,         p3_u3460, p3_u3461, p3_u3462, p3_u3463, p3_u3464, p3_u3465, p3_u3466,         p3_u3467, p3_u3468, p3_u3469, p3_u3470, p3_u3471, p3_u3472, p3_u3473,         p3_u3474, p3_u3475, p3_u3476, p3_u3477, p3_u3478, p3_u3479, p3_u3480,         p3_u3481, p3_u3482, p3_u3483, p3_u3484, p3_u3485, p3_u3486, p3_u3487,         p3_u3488, p3_u3489, p3_u3490, p3_u3233, p3_u3232, p3_u3231, p3_u3230,         p3_u3229, p3_u3228, p3_u3227, p3_u3226, p3_u3225, p3_u3224, p3_u3223,         p3_u3222, p3_u3221, p3_u3220, p3_u3219, p3_u3218, p3_u3217, p3_u3216,         p3_u3215, p3_u3214, p3_u3213, p3_u3212, p3_u3211, p3_u3210, p3_u3209,         p3_u3208, p3_u3207, p3_u3206, p3_u3205, p3_u3204, p3_u3203, p3_u3202,         p3_u3201, p3_u3200, p3_u3199, p3_u3198, p3_u3197, p3_u3196, p3_u3195,         p3_u3194, p3_u3193, p3_u3192, p3_u3191, p3_u3190, p3_u3189, p3_u3188,         p3_u3187, p3_u3186, p3_u3185, p3_u3184, p3_u3183, p3_u3182, p3_u3491,         p3_u3492, p3_u3493, p3_u3494, p3_u3495, p3_u3496, p3_u3497, p3_u3498,         p3_u3499, p3_u3500, p3_u3501, p3_u3502, p3_u3503, p3_u3504, p3_u3505,         p3_u3506, p3_u3507, p3_u3508, p3_u3509, p3_u3510, p3_u3511, p3_u3512,         p3_u3513, p3_u3514, p3_u3515, p3_u3516, p3_u3517, p3_u3518, p3_u3519,         p3_u3520, p3_u3521, p3_u3522, p3_u3296, p3_u3181, p3_u3180, p3_u3179,         p3_u3178, p3_u3177, p3_u3176, p3_u3175, p3_u3174, p3_u3173, p3_u3172,         p3_u3171, p3_u3170, p3_u3169, p3_u3168, p3_u3167, p3_u3166, p3_u3165,         p3_u3164, p3_u3163, p3_u3162, p3_u3161, p3_u3160, p3_u3159, p3_u3158,         p3_u3157, p3_u3156, p3_u3155, p3_u3154, p3_u3153, p3_u3151, p3_u3150,         p3_u3897;
wire   n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,         n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,         n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928,         n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936,         n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944,         n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952,         n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,         n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968,         n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976,         n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984,         n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,         n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000,         n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008,         n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016,         n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,         n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032,         n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040,         n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048,         n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056,         n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,         n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072,         n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080,         n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,         n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096,         n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104,         n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112,         n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120,         n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128,         n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136,         n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144,         n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152,         n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160,         n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168,         n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176,         n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184,         n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192,         n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200,         n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208,         n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216,         n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224,         n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232,         n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240,         n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248,         n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256,         n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264,         n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272,         n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280,         n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288,         n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296,         n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304,         n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312,         n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320,         n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328,         n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336,         n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344,         n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352,         n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360,         n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368,         n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376,         n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384,         n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392,         n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400,         n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408,         n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416,         n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424,         n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432,         n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440,         n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448,         n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456,         n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464,         n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472,         n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480,         n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488,         n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496,         n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504,         n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512,         n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520,         n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528,         n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536,         n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544,         n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552,         n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560,         n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568,         n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576,         n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584,         n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592,         n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600,         n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608,         n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616,         n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624,         n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632,         n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640,         n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648,         n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656,         n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664,         n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672,         n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680,         n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688,         n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696,         n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704,         n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712,         n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720,         n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728,         n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736,         n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744,         n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752,         n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760,         n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768,         n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776,         n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784,         n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792,         n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800,         n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808,         n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816,         n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824,         n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832,         n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840,         n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848,         n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856,         n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864,         n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872,         n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880,         n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888,         n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896,         n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904,         n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912,         n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920,         n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928,         n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936,         n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944,         n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952,         n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960,         n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968,         n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976,         n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984,         n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992,         n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000,         n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008,         n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016,         n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024,         n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032,         n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040,         n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048,         n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056,         n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064,         n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072,         n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080,         n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088,         n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096,         n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104,         n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112,         n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120,         n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128,         n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136,         n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144,         n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152,         n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160,         n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168,         n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176,         n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184,         n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192,         n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200,         n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208,         n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216,         n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224,         n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232,         n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240,         n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248,         n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256,         n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264,         n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272,         n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280,         n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288,         n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296,         n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304,         n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312,         n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320,         n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328,         n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336,         n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344,         n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352,         n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360,         n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368,         n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376,         n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384,         n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392,         n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400,         n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408,         n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416,         n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424,         n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432,         n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440,         n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448,         n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456,         n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464,         n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472,         n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480,         n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488,         n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496,         n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504,         n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512,         n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520,         n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528,         n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536,         n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544,         n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552,         n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560,         n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568,         n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576,         n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584,         n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592,         n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600,         n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608,         n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616,         n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624,         n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632,         n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640,         n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648,         n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656,         n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664,         n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672,         n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680,         n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688,         n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696,         n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704,         n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712,         n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720,         n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728,         n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736,         n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744,         n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752,         n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760,         n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768,         n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776,         n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784,         n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792,         n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800,         n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808,         n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816,         n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824,         n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832,         n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840,         n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848,         n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856,         n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864,         n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872,         n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880,         n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888,         n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896,         n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904,         n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912,         n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920,         n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928,         n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936,         n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944,         n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952,         n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960,         n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968,         n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976,         n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984,         n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992,         n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000,         n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008,         n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016,         n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024,         n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032,         n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040,         n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048,         n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056,         n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064,         n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072,         n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080,         n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088,         n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096,         n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104,         n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112,         n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120,         n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128,         n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136,         n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144,         n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152,         n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160,         n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168,         n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176,         n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184,         n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192,         n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200,         n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208,         n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216,         n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224,         n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232,         n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240,         n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248,         n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256,         n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264,         n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272,         n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280,         n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288,         n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296,         n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304,         n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312,         n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320,         n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328,         n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336,         n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344,         n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352,         n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360,         n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368,         n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376,         n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384,         n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392,         n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400,         n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408,         n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416,         n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424,         n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432,         n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440,         n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448,         n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456,         n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464,         n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472,         n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480,         n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488,         n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496,         n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504,         n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512,         n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520,         n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528,         n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536,         n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544,         n23545, n23546, n23547, n23548, n23549, n23550, n23551, n23552,         n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560,         n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568,         n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576,         n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584,         n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592,         n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600,         n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608,         n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616,         n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624,         n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632,         n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640,         n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648,         n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656,         n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664,         n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672,         n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680,         n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688,         n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696,         n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704,         n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712,         n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720,         n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728,         n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736,         n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744,         n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752,         n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760,         n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768,         n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776,         n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784,         n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792,         n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800,         n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808,         n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816,         n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824,         n23825, n23826, n23827, n23828, n23829, n23830, n23831, n23832,         n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840,         n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848,         n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856,         n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864,         n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872,         n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880,         n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888,         n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896,         n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904,         n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23912,         n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920,         n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928,         n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936,         n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944,         n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952,         n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960,         n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968,         n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976,         n23977, n23978, n23979, n23980, n23981, n23982, n23983, n23984,         n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992,         n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000,         n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008,         n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016,         n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024,         n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032,         n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040,         n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048,         n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056,         n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064,         n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072,         n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080,         n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088,         n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096,         n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104,         n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112,         n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120,         n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128,         n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136,         n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144,         n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152,         n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160,         n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168,         n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176,         n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184,         n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192,         n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200,         n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208,         n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216,         n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224,         n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232,         n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240,         n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248,         n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256,         n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264,         n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272,         n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280,         n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288,         n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296,         n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304,         n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312,         n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24320,         n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328,         n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336,         n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344,         n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352,         n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360,         n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368,         n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376,         n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384,         n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392,         n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400,         n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408,         n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416,         n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424,         n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432,         n24433, n24434, n24435, n24436, n24437, n24438, n24439, n24440,         n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448,         n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456,         n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464,         n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24472,         n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480,         n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488,         n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496,         n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504,         n24505, n24506, n24507, n24508, n24509, n24510, n24511, n24512,         n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520,         n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528,         n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536,         n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544,         n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552,         n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560,         n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568,         n24569, n24570, n24571, n24572, n24573, n24574, n24575, n24576,         n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584,         n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592,         n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600,         n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608,         n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616,         n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624,         n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632,         n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640,         n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648,         n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656,         n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664,         n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672,         n24673, n24674, n24675, n24676, n24677, n24678, n24679, n24680,         n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688,         n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696,         n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704,         n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712,         n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720,         n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24728,         n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736,         n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744,         n24745, n24746, n24747, n24748, n24749, n24750, n24751, n24752,         n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760,         n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768,         n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776,         n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784,         n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792,         n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800,         n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808,         n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816,         n24817, n24818, n24819, n24820, n24821, n24822, n24823, n24824,         n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832,         n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840,         n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848,         n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856,         n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864,         n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872,         n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880,         n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888,         n24889, n24890, n24891, n24892, n24893, n24894, n24895, n24896,         n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904,         n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912,         n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920,         n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928,         n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936,         n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944,         n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952,         n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960,         n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968,         n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976,         n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984,         n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992,         n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000,         n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008,         n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016,         n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024,         n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032,         n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040,         n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048,         n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056,         n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064,         n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072,         n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080,         n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088,         n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096,         n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104,         n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112,         n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120,         n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128,         n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136,         n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144,         n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152,         n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160,         n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168,         n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176,         n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184,         n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192,         n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200,         n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208,         n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216,         n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224,         n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232,         n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240,         n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248,         n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256,         n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264,         n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272,         n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280,         n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288,         n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296,         n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304,         n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312,         n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320,         n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328,         n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336,         n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344,         n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352,         n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360,         n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368,         n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376,         n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384,         n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392,         n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400,         n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408,         n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416,         n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424,         n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432,         n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440,         n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448,         n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456,         n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464,         n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472,         n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480,         n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488,         n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496,         n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504,         n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512,         n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520,         n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528,         n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536,         n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544,         n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552,         n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560,         n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568,         n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576,         n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584,         n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592,         n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600,         n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608,         n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616,         n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624,         n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632,         n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640,         n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648,         n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656,         n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664,         n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672,         n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680,         n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688,         n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696,         n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704,         n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712,         n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720,         n25721, n25722, n25723, n25724, n25725, n25726, n25727, n25728,         n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736,         n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744,         n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752,         n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760,         n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768,         n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776,         n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784,         n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792,         n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800,         n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808,         n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816,         n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824,         n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832,         n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840,         n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848,         n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856,         n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864,         n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872,         n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880,         n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888,         n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896,         n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904,         n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912,         n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920,         n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928,         n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936,         n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944,         n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952,         n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960,         n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968,         n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976,         n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984,         n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992,         n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26000,         n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008,         n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016,         n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024,         n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032,         n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040,         n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048,         n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056,         n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064,         n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072,         n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080,         n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088,         n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096,         n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104,         n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112,         n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120,         n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128,         n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136,         n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144,         n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152,         n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160,         n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168,         n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176,         n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184,         n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192,         n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200,         n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208,         n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216,         n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224,         n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232,         n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240,         n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248,         n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256,         n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26264,         n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272,         n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280,         n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288,         n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296,         n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304,         n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312,         n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320,         n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328,         n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336,         n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344,         n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352,         n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360,         n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368,         n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376,         n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384,         n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392,         n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400,         n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408,         n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416,         n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424,         n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432,         n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440,         n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448,         n26449, n26450, n26451, n26452, n26453, n26454, n26455, n26456,         n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464,         n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472,         n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480,         n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488,         n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496,         n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504,         n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512,         n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520,         n26521, n26522, n26523, n26524, n26525, n26526, n26527, n26528,         n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536,         n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544,         n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552,         n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560,         n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568,         n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576,         n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584,         n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592,         n26593, n26594, n26595, n26596, n26597, n26598, n26599, n26600,         n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608,         n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616,         n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624,         n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632,         n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640,         n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648,         n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656,         n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664,         n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672,         n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680,         n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688,         n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696,         n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704,         n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712,         n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720,         n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728,         n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736,         n26737, n26738, n26739, n26740, n26741, n26742, n26743, n26744,         n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752,         n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760,         n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768,         n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776,         n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784,         n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792,         n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800,         n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808,         n26809, n26810, n26811, n26812, n26813, n26814, n26815, n26816,         n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824,         n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832,         n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840,         n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848,         n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856,         n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864,         n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872,         n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880,         n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888,         n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896,         n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904,         n26905, n26906, n26907, n26908, n26909, n26910, n26911, n26912,         n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920,         n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928,         n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936,         n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944,         n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952,         n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960,         n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968,         n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976,         n26977, n26978, n26979, n26980, n26981, n26982, n26983, n26984,         n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992,         n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000,         n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008,         n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016,         n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024,         n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032,         n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040,         n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048,         n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056,         n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064,         n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072,         n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080,         n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088,         n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096,         n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104,         n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112,         n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120,         n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128,         n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136,         n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144,         n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152,         n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160,         n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168,         n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176,         n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184,         n27185, n27186, n27187, n27188, n27189, n27190, n27191, n27192,         n27193, n27194, n27195, n27196, n27197, n27198, n27199, n27200,         n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208,         n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216,         n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224,         n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232,         n27233, n27234, n27235, n27236, n27237, n27238, n27239, n27240,         n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248,         n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256,         n27257, n27258, n27259, n27260, n27261, n27262, n27263, n27264,         n27265, n27266, n27267, n27268, n27269, n27270, n27271, n27272,         n27273, n27274, n27275, n27276, n27277, n27278, n27279, n27280,         n27281, n27282, n27283, n27284, n27285, n27286, n27287, n27288,         n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296,         n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304,         n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312,         n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320,         n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328,         n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336,         n27337, n27338, n27339, n27340, n27341, n27342, n27343, n27344,         n27345, n27346, n27347, n27348, n27349, n27350, n27351, n27352,         n27353, n27354, n27355, n27356, n27357, n27358, n27359, n27360,         n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368,         n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376,         n27377, n27378, n27379, n27380, n27381, n27382, n27383, n27384,         n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392,         n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400,         n27401, n27402, n27403, n27404, n27405, n27406, n27407, n27408,         n27409, n27410, n27411, n27412, n27413, n27414, n27415, n27416,         n27417, n27418, n27419, n27420, n27421, n27422, n27423, n27424,         n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432,         n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440,         n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448,         n27449, n27450, n27451, n27452, n27453, n27454, n27455, n27456,         n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464,         n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472,         n27473, n27474, n27475, n27476, n27477, n27478, n27479, n27480,         n27481, n27482, n27483, n27484, n27485, n27486, n27487, n27488,         n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496,         n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504,         n27505, n27506, n27507, n27508, n27509, n27510, n27511, n27512,         n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520,         n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528,         n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536,         n27537, n27538, n27539, n27540, n27541, n27542, n27543, n27544,         n27545, n27546, n27547, n27548, n27549, n27550, n27551, n27552,         n27553, n27554, n27555, n27556;

   nand U14304 ( n15991,n16257,n16172 );
   nand U14305 ( n15992,n16258,n16259 );
   not U14306 ( n20291,n20314 );
   not U14307 ( n24254,p1_ir_reg_31_ );
   nand U14308 ( n16692,n17520,n15559 );
   nor U14309 ( n15567,n18437,p3_u3151,n15944 );
   nand U14310 ( n16630,n16260,n16264 );
   nand U14311 ( n24400,n26133,n25806 );
   not U14312 ( n18499,n18453 );
   nor U14313 ( n18830,n17554,n18453 );
   nor U14314 ( n18674,n15340,n18453 );
   nor U14315 ( n18703,n17536,n18453 );
   nor U14316 ( n18842,n17440,n18453 );
   nor U14317 ( n18633,n15873,n18453 );
   nand U14318 ( n16628,n16264,n17480,n15943 );
   nor U14319 ( n17591,n19438,n19439 );
   nor U14320 ( n26179,n27446,n27447 );
   nor U14321 ( n21827,n23302,n23303 );
   nand U14322 ( n23606,n25105,n25264 );
   nand U14323 ( n16598,n15559,n15560,n16604 );
   nand U14324 ( n18470,n15805,n17520,n15810 );
   nand U14325 ( n24395,n26133,n25787 );
   nand U14326 ( n21040,n23307,n20139 );
   nand U14327 ( n15828,n16264,n16257,n15577 );
   not U14328 ( n15310,n15398 );
   nor U14329 ( n17592,n19438,n19437 );
   nor U14330 ( n26178,n27446,n27445 );
   nor U14331 ( n21826,n23302,n23301 );
   not U14332 ( n19777,n19739 );
   nor U14333 ( n19739,n20145,n20228 );
   not U14334 ( n22488,n22451 );
   not U14335 ( n18921,n17657 );
   nand U14336 ( n21222,n20910,n21760 );
   not U14337 ( n17734,n17825 );
   nand U14338 ( n17825,n15937,n18430 );
   nand U14339 ( n24449,n25104,n24012 );
   not U14340 ( n21939,n21969 );
   not U14341 ( n26222,n26299 );
   nor U14342 ( n22954,n16576,n21918 );
   not U14343 ( n21918,n21921 );
   not U14344 ( n21957,n22413 );
   nand U14345 ( n23621,n23978,n23979 );
   nand U14346 ( n15831,n17480,n16257,n16264 );
   not U14347 ( n17708,n17823 );
   nand U14348 ( n17823,n17659,n18430 );
   and U14349 ( n18456,n15567,n19295 );
   and U14350 ( n21825,n23303,n23302 );
   and U14351 ( n17590,n19439,n19438 );
   and U14352 ( n26177,n27447,n27446 );
   nand U14353 ( n24265,n27529,n27530,n27531 );
   or U14354 ( n16590,n19501,n19504 );
   not U14355 ( p2_u3088,p2_state_reg );
   nand U14356 ( n19776,n21828,n20148 );
   nor U14357 ( n16641,n17662,n16603 );
   nand U14358 ( n24302,n25112,n24012 );
   nand U14359 ( n26547,n27435,n27436 );
   nand U14360 ( n23608,n25105,n25106 );
   not U14361 ( n15290,n15341 );
   nand U14362 ( n19759,n20149,n20137 );
   nand U14363 ( n20915,n20910,n19739 );
   nand U14364 ( n25861,n26171,n24395,n26127,n26211 );
   nand U14365 ( n22605,n22432,n21040,n23306,n21042 );
   nor U14366 ( n16316,n16315,p3_u3151 );
   not U14367 ( n23994,n23993 );
   nand U14368 ( n23993,n23566,n24265 );
   not U14369 ( n15814,n15813 );
   nand U14370 ( n15813,n15567,n16590 );
   nand U14371 ( n24394,n25785,n23990 );
   not U14372 ( n16602,n16640 );
   nand U14373 ( n16640,n17685,n16604 );
   not U14374 ( n22469,n22452 );
   nand U14375 ( n16631,n15943,n17480,n15946 );
   not U14376 ( n25265,n27492 );
   not U14377 ( n21958,n22429 );
   nor U14378 ( n22956,n16572,n21918 );
   nand U14379 ( n20608,n20167,n21948,n22434 );
   not U14380 ( n16642,n16599 );
   not U14381 ( n22449,n22557 );
   nand U14382 ( n16634,n15578,n16260 );
   not U14383 ( n15602,n15618 );
   nand U14384 ( n21949,n20217,n22424 );
   nand U14385 ( n18452,n15805,n15560,n15810 );
   nand U14386 ( n19760,n20137,n20138,n20139 );
   not U14387 ( n26225,n26298 );
   not U14388 ( n26240,n26223 );
   nor U14389 ( n17640,n16572,n18921 );
   not U14390 ( n25283,n25567 );
   not U14391 ( n17719,n17763 );
   nand U14392 ( n17763,p3_u3897,n18431 );
   nor U14393 ( n17643,n16576,n18921 );
   not U14394 ( n17731,n15937 );
   nand U14395 ( n15937,n19532,n19533,n16553 );
   nand U14396 ( n20294,n20566,n20591 );
   nor U14397 ( n20617,n16576,p2_state_reg );
   not U14398 ( n25298,n25684 );
   and U14399 ( n22798,n23301,n23302 );
   and U14400 ( n26563,n27445,n27446 );
   not U14401 ( n24009,n24282 );
   nor U14402 ( n16317,n16572,p3_state_reg );
   not U14403 ( n20290,n20315 );
   not U14404 ( n20153,n20152 );
   not U14405 ( n26543,n27435 );
   not U14406 ( n23575,n23742 );
   nand U14407 ( n24281,n24012,n25267 );
   and U14408 ( n18768,n19437,n19438 );
   nand U14409 ( n25856,n26127,n24395,n26128 );
   nand U14410 ( n25860,n26131,n24347,n26132 );
   not U14411 ( n23624,n23573 );
   not U14412 ( n15295,n15289 );
   nand U14413 ( n15289,n15566,n15567,n15568,n15569 );
   nor U14414 ( n20613,n16572,p2_state_reg );
   not U14415 ( n23569,n23577 );
   nand U14416 ( n23577,n23564,n23980,n23566 );
   not U14417 ( n23468,n23470 );
   nand U14418 ( n23470,n23564,n23565,n23566 );
   not U14419 ( n19735,n19743 );
   nand U14420 ( n19743,n19732,n20140 );
   not U14421 ( n19635,n19637 );
   nand U14422 ( n19637,n19731,n19732 );
   nor U14423 ( n24041,n16572,p1_state_reg );
   nor U14424 ( n24045,n16576,p1_state_reg );
   nor U14425 ( n16313,n16576,p3_state_reg );
   and U14426 ( n15589,n15592,n15562 );
   nor U14427 ( n26136,n16572,n25265 );
   nor U14428 ( n26140,n16576,n25265 );
   nand U14429 ( n19774,n20148,n20216 );
   not U14430 ( n26652,n26364 );
   nand U14431 ( n26364,n27436,n27437,n27438 );
   not U14432 ( p2_u3947,n19538 );
   nand U14433 ( n19538,n22436,p2_state_reg,n22437 );
   not U14434 ( p1_u4016,n23371 );
   nand U14435 ( n23371,n25791,p1_state_reg,n25790 );
   not U14436 ( p3_u3897,n15191 );
   nand U14437 ( n15191,n15824,p3_state_reg,n18437 );
   not U14438 ( n20916,n20932 );
   not U14439 ( p3_u3151,p3_state_reg );
   nand U14440 ( n25857,n26185,n24347,n26186 );
   nand U14441 ( n24347,n26188,n25787 );
   nor U14442 ( n24044,n24043,p1_u3086 );
   not U14443 ( n24043,n24073 );
   not U14444 ( n24012,n24011 );
   nand U14445 ( n24011,n23566,n25268 );
   not U14446 ( n16604,n16603 );
   nand U14447 ( n16603,n15567,n17686 );
   not U14448 ( n18859,n18755 );
   nand U14449 ( n18755,n17522,n15942,n19442 );
   not U14450 ( n15588,n15592 );
   nand U14451 ( n15592,n15798,n15799 );
   not U14452 ( n20910,n20902 );
   nand U14453 ( n20902,n20141,n21928 );
   not U14454 ( n16572,n16576 );
   nand U14455 ( n16576,n27493,n27494 );
   nor U14456 ( n20616,n20615,p2_u3088 );
   not U14457 ( n14937,n22788 );
   not U14458 ( n22788,n22785 );
   nor U14459 ( n22785,n20168,n20149,n23307 );
   nor U14460 ( n26542,n25783,n25790 );
   or U14461 ( u29,p3_rd_reg,n14938 );
   xor U14462 ( n14938,n14939,p1_rd_reg );
   nand U14463 ( u28,n14940,n14941 );
   not U14464 ( n14941,p3_wr_reg );
   xor U14465 ( n14940,p2_wr_reg,p1_wr_reg );
   xor U14466 ( sub_1596_u70,n14942,n14943 );
   xor U14467 ( n14943,p2_addr_reg_10_,n14944 );
   xor U14468 ( sub_1596_u69,n14945,n14946 );
   xor U14469 ( n14946,p2_addr_reg_11_,n14947 );
   xor U14470 ( sub_1596_u68,n14948,n14949 );
   xor U14471 ( n14949,p2_addr_reg_12_,n14950 );
   xor U14472 ( sub_1596_u67,n14951,n14952 );
   xor U14473 ( n14952,p2_addr_reg_13_,n14953 );
   xor U14474 ( sub_1596_u66,n14954,n14955 );
   xor U14475 ( n14955,p2_addr_reg_14_,n14956 );
   xor U14476 ( sub_1596_u65,n14957,n14958 );
   xor U14477 ( n14958,p2_addr_reg_15_,n14959 );
   xor U14478 ( sub_1596_u64,n14960,n14961 );
   xor U14479 ( n14961,p2_addr_reg_16_,n14962 );
   xor U14480 ( sub_1596_u63,n14963,n14964 );
   xor U14481 ( n14964,p2_addr_reg_17_,n14965 );
   xor U14482 ( sub_1596_u62,n14966,n14967 );
   xor U14483 ( n14967,p2_addr_reg_18_,n14968 );
   xor U14484 ( sub_1596_u61,n14969,n14970 );
   xor U14485 ( n14970,n14971,p2_addr_reg_2_ );
   xor U14486 ( sub_1596_u60,n14972,n14973 );
   xor U14487 ( n14973,n14974,n14975 );
   not U14488 ( n14972,n14976 );
   xor U14489 ( sub_1596_u59,n14977,n14978 );
   xor U14490 ( n14977,n14979,p2_addr_reg_4_ );
   xor U14491 ( sub_1596_u58,n14980,n14981 );
   xor U14492 ( n14980,n14982,p2_addr_reg_5_ );
   xor U14493 ( sub_1596_u57,n14983,n14984 );
   xor U14494 ( n14983,n14985,p2_addr_reg_6_ );
   xor U14495 ( sub_1596_u56,n14986,n14987 );
   xor U14496 ( n14987,p2_addr_reg_7_,n14988 );
   xor U14497 ( sub_1596_u55,n14989,n14990 );
   xor U14498 ( n14990,p2_addr_reg_8_,n14991 );
   xor U14499 ( sub_1596_u54,n14992,n14993 );
   xor U14500 ( n14993,p2_addr_reg_9_,n14994 );
   xor U14501 ( sub_1596_u53,p2_addr_reg_0_,n14995 );
   xor U14502 ( sub_1596_u5,n14996,n14997 );
   xor U14503 ( n14996,p2_addr_reg_1_,n14998 );
   xor U14504 ( sub_1596_u4,n14999,n15000 );
   nand U14505 ( n15000,n15001,n15002 );
   nand U14506 ( n15002,p2_addr_reg_18_,n15003 );
   nand U14507 ( n15003,n14966,n14968 );
   or U14508 ( n15001,n14966,n14968 );
   nand U14509 ( n14968,n15004,n15005 );
   nand U14510 ( n15005,n15006,n15007 );
   not U14511 ( n15007,p2_addr_reg_17_ );
   or U14512 ( n15006,n14963,n14965 );
   nand U14513 ( n15004,n14963,n14965 );
   nand U14514 ( n14965,n15008,n15009 );
   nand U14515 ( n15009,n15010,n15011 );
   not U14516 ( n15011,p2_addr_reg_16_ );
   or U14517 ( n15010,n14960,n14962 );
   nand U14518 ( n15008,n14960,n14962 );
   nand U14519 ( n14962,n15012,n15013 );
   nand U14520 ( n15013,n15014,n15015 );
   not U14521 ( n15015,p2_addr_reg_15_ );
   or U14522 ( n15014,n14957,n14959 );
   nand U14523 ( n15012,n14957,n14959 );
   nand U14524 ( n14959,n15016,n15017 );
   nand U14525 ( n15017,n15018,n15019 );
   not U14526 ( n15019,p2_addr_reg_14_ );
   or U14527 ( n15018,n14954,n14956 );
   nand U14528 ( n15016,n14954,n14956 );
   nand U14529 ( n14956,n15020,n15021 );
   nand U14530 ( n15021,n15022,n15023 );
   not U14531 ( n15023,p2_addr_reg_13_ );
   or U14532 ( n15022,n14951,n14953 );
   nand U14533 ( n15020,n14951,n14953 );
   nand U14534 ( n14953,n15024,n15025 );
   nand U14535 ( n15025,n15026,n15027 );
   not U14536 ( n15027,p2_addr_reg_12_ );
   or U14537 ( n15026,n14948,n14950 );
   nand U14538 ( n15024,n14948,n14950 );
   nand U14539 ( n14950,n15028,n15029 );
   nand U14540 ( n15029,n15030,n15031 );
   not U14541 ( n15031,p2_addr_reg_11_ );
   or U14542 ( n15030,n14945,n14947 );
   nand U14543 ( n15028,n14945,n14947 );
   nand U14544 ( n14947,n15032,n15033 );
   nand U14545 ( n15033,n15034,n15035 );
   not U14546 ( n15035,p2_addr_reg_10_ );
   or U14547 ( n15034,n14942,n14944 );
   nand U14548 ( n15032,n14942,n14944 );
   nand U14549 ( n14944,n15036,n15037 );
   nand U14550 ( n15037,n15038,n15039 );
   not U14551 ( n15039,p2_addr_reg_9_ );
   or U14552 ( n15038,n14994,n14992 );
   nand U14553 ( n15036,n14992,n14994 );
   nand U14554 ( n14994,n15040,n15041 );
   nand U14555 ( n15041,n15042,n15043 );
   not U14556 ( n15043,p2_addr_reg_8_ );
   or U14557 ( n15042,n14991,n14989 );
   nand U14558 ( n15040,n14989,n14991 );
   nand U14559 ( n14991,n15044,n15045 );
   nand U14560 ( n15045,n15046,n15047 );
   not U14561 ( n15047,p2_addr_reg_7_ );
   or U14562 ( n15046,n14988,n14986 );
   nand U14563 ( n15044,n14986,n14988 );
   nand U14564 ( n14988,n15048,n15049 );
   nand U14565 ( n15049,n15050,n15051 );
   not U14566 ( n15051,p2_addr_reg_6_ );
   nand U14567 ( n15050,n14985,n14984 );
   or U14568 ( n15048,n14984,n14985 );
   and U14569 ( n14985,n15052,n15053 );
   nand U14570 ( n15053,n15054,n15055 );
   not U14571 ( n15055,p2_addr_reg_5_ );
   nand U14572 ( n15054,n14982,n14981 );
   or U14573 ( n15052,n14981,n14982 );
   and U14574 ( n14982,n15056,n15057 );
   nand U14575 ( n15057,n15058,n15059 );
   not U14576 ( n15059,p2_addr_reg_4_ );
   or U14577 ( n15058,n14979,n14978 );
   nand U14578 ( n15056,n14978,n14979 );
   nand U14579 ( n14979,n15060,n15061 );
   nand U14580 ( n15061,n15062,n14975 );
   not U14581 ( n14975,p2_addr_reg_3_ );
   nand U14582 ( n15062,n14976,n14974 );
   or U14583 ( n15060,n14974,n14976 );
   xor U14584 ( n14976,n15063,n15064 );
   xor U14585 ( n15063,p3_addr_reg_3_,p1_addr_reg_3_ );
   nand U14586 ( n14974,n15065,n15066 );
   nand U14587 ( n15066,p2_addr_reg_2_,n15067 );
   nand U14588 ( n15067,n14969,n14971 );
   or U14589 ( n15065,n14971,n14969 );
   xor U14590 ( n14969,n15068,n15069 );
   xor U14591 ( n15068,p3_addr_reg_2_,p1_addr_reg_2_ );
   nand U14592 ( n14971,n15070,n15071 );
   nand U14593 ( n15071,n15072,n15073 );
   not U14594 ( n15073,p2_addr_reg_1_ );
   or U14595 ( n15072,n14998,n14997 );
   nand U14596 ( n15070,n14997,n14998 );
   nand U14597 ( n14998,p2_addr_reg_0_,n14995 );
   nand U14598 ( n14995,n15074,n15075 );
   nand U14599 ( n15075,p1_addr_reg_0_,n15076 );
   xor U14600 ( n14997,n15077,n15074 );
   xor U14601 ( n15077,p3_addr_reg_1_,p1_addr_reg_1_ );
   xor U14602 ( n14978,n15078,n15079 );
   xor U14603 ( n15078,p3_addr_reg_4_,p1_addr_reg_4_ );
   xor U14604 ( n14981,n15080,n15081 );
   xor U14605 ( n15080,p3_addr_reg_5_,p1_addr_reg_5_ );
   xor U14606 ( n14984,n15082,n15083 );
   xor U14607 ( n15082,p3_addr_reg_6_,p1_addr_reg_6_ );
   xor U14608 ( n14986,n15084,n15085 );
   xor U14609 ( n15084,p3_addr_reg_7_,n15086 );
   xor U14610 ( n14989,n15087,n15088 );
   xor U14611 ( n15087,p3_addr_reg_8_,n15089 );
   xor U14612 ( n14992,n15090,n15091 );
   xor U14613 ( n15090,p3_addr_reg_9_,n15092 );
   xor U14614 ( n14942,n15093,n15094 );
   xor U14615 ( n15093,p3_addr_reg_10_,p1_addr_reg_10_ );
   xor U14616 ( n14945,n15095,n15096 );
   xor U14617 ( n15095,p3_addr_reg_11_,p1_addr_reg_11_ );
   xor U14618 ( n14948,n15097,n15098 );
   xor U14619 ( n15097,p3_addr_reg_12_,p1_addr_reg_12_ );
   xor U14620 ( n14951,n15099,n15100 );
   xor U14621 ( n15099,p3_addr_reg_13_,p1_addr_reg_13_ );
   xor U14622 ( n14954,n15101,n15102 );
   xor U14623 ( n15101,p3_addr_reg_14_,p1_addr_reg_14_ );
   xor U14624 ( n14957,n15103,n15104 );
   xor U14625 ( n15103,p3_addr_reg_15_,p1_addr_reg_15_ );
   xor U14626 ( n14960,n15105,n15106 );
   xor U14627 ( n15105,p3_addr_reg_16_,p1_addr_reg_16_ );
   xor U14628 ( n14963,n15107,n15108 );
   xor U14629 ( n15107,p3_addr_reg_17_,p1_addr_reg_17_ );
   xor U14630 ( n14966,n15109,n15110 );
   xor U14631 ( n15109,p3_addr_reg_18_,p1_addr_reg_18_ );
   xor U14632 ( n14999,p2_addr_reg_19_,n15111 );
   nand U14633 ( n15111,n15112,n15113 );
   nand U14634 ( n15113,n15114,n15115,n15116 );
   xor U14635 ( n15116,p3_addr_reg_19_,n15117 );
   nand U14636 ( n15115,n15118,n15119 );
   not U14637 ( n15119,p3_addr_reg_18_ );
   nand U14638 ( n15112,n15118,n15120,n15121 );
   xor U14639 ( n15121,p3_addr_reg_19_,p1_addr_reg_19_ );
   nand U14640 ( n15120,p3_addr_reg_18_,n15114 );
   nand U14641 ( n15114,n15110,p1_addr_reg_18_ );
   not U14642 ( n15110,n15122 );
   nand U14643 ( n15118,n15123,n15122 );
   nand U14644 ( n15122,n15124,n15125 );
   nand U14645 ( n15125,p3_addr_reg_17_,n15126 );
   nand U14646 ( n15126,n15108,p1_addr_reg_17_ );
   not U14647 ( n15108,n15127 );
   nand U14648 ( n15124,n15127,n15128 );
   nand U14649 ( n15127,n15129,n15130 );
   nand U14650 ( n15130,p3_addr_reg_16_,n15131 );
   nand U14651 ( n15131,n15106,p1_addr_reg_16_ );
   or U14652 ( n15129,n15106,p1_addr_reg_16_ );
   and U14653 ( n15106,n15132,n15133 );
   nand U14654 ( n15133,p3_addr_reg_15_,n15134 );
   nand U14655 ( n15134,n15104,p1_addr_reg_15_ );
   or U14656 ( n15132,n15104,p1_addr_reg_15_ );
   and U14657 ( n15104,n15135,n15136 );
   nand U14658 ( n15136,p3_addr_reg_14_,n15137 );
   nand U14659 ( n15137,n15102,p1_addr_reg_14_ );
   or U14660 ( n15135,n15102,p1_addr_reg_14_ );
   and U14661 ( n15102,n15138,n15139 );
   nand U14662 ( n15139,p3_addr_reg_13_,n15140 );
   nand U14663 ( n15140,n15100,p1_addr_reg_13_ );
   not U14664 ( n15100,n15141 );
   nand U14665 ( n15138,n15141,n15142 );
   nand U14666 ( n15141,n15143,n15144 );
   nand U14667 ( n15144,p3_addr_reg_12_,n15145 );
   nand U14668 ( n15145,n15098,p1_addr_reg_12_ );
   not U14669 ( n15098,n15146 );
   nand U14670 ( n15143,n15146,n15147 );
   nand U14671 ( n15146,n15148,n15149 );
   nand U14672 ( n15149,p3_addr_reg_11_,n15150 );
   nand U14673 ( n15150,n15096,p1_addr_reg_11_ );
   or U14674 ( n15148,n15096,p1_addr_reg_11_ );
   and U14675 ( n15096,n15151,n15152 );
   nand U14676 ( n15152,p3_addr_reg_10_,n15153 );
   nand U14677 ( n15153,n15094,p1_addr_reg_10_ );
   not U14678 ( n15094,n15154 );
   nand U14679 ( n15151,n15154,n15155 );
   nand U14680 ( n15154,n15156,n15157 );
   nand U14681 ( n15157,p3_addr_reg_9_,n15158 );
   or U14682 ( n15158,n15092,n15091 );
   nand U14683 ( n15156,n15091,n15092 );
   nand U14684 ( n15091,n15159,n15160 );
   nand U14685 ( n15160,p3_addr_reg_8_,n15161 );
   or U14686 ( n15161,n15089,n15088 );
   nand U14687 ( n15159,n15088,n15089 );
   nand U14688 ( n15088,n15162,n15163 );
   nand U14689 ( n15163,p3_addr_reg_7_,n15164 );
   or U14690 ( n15164,n15086,n15085 );
   nand U14691 ( n15162,n15085,n15086 );
   nand U14692 ( n15085,n15165,n15166 );
   nand U14693 ( n15166,p3_addr_reg_6_,n15167 );
   or U14694 ( n15167,n15168,n15083 );
   nand U14695 ( n15165,n15083,n15168 );
   nand U14696 ( n15083,n15169,n15170 );
   nand U14697 ( n15170,p3_addr_reg_5_,n15171 );
   or U14698 ( n15171,n15172,n15081 );
   nand U14699 ( n15169,n15081,n15172 );
   nand U14700 ( n15081,n15173,n15174 );
   nand U14701 ( n15174,p3_addr_reg_4_,n15175 );
   nand U14702 ( n15175,p1_addr_reg_4_,n15079 );
   or U14703 ( n15173,n15079,p1_addr_reg_4_ );
   and U14704 ( n15079,n15176,n15177 );
   nand U14705 ( n15177,p3_addr_reg_3_,n15178 );
   or U14706 ( n15178,n15179,n15064 );
   nand U14707 ( n15176,n15064,n15179 );
   nand U14708 ( n15064,n15180,n15181 );
   nand U14709 ( n15181,p3_addr_reg_2_,n15182 );
   nand U14710 ( n15182,p1_addr_reg_2_,n15069 );
   or U14711 ( n15180,n15069,p1_addr_reg_2_ );
   nand U14712 ( n15069,n15183,n15184 );
   nand U14713 ( n15184,n15185,n15186 );
   not U14714 ( n15186,p3_addr_reg_1_ );
   nand U14715 ( n15185,n15187,n15188 );
   nand U14716 ( n15183,p1_addr_reg_1_,n15074 );
   not U14717 ( n15074,n15187 );
   nor U14718 ( n15187,n15076,p1_addr_reg_0_ );
   not U14719 ( n15123,p1_addr_reg_18_ );
   nand U14720 ( p3_u3522,n15189,n15190 );
   nand U14721 ( n15190,p3_datao_reg_31_,n15191 );
   nand U14722 ( n15189,p3_u3897,n15192 );
   nand U14723 ( p3_u3521,n15193,n15194 );
   nand U14724 ( n15194,p3_datao_reg_30_,n15191 );
   nand U14725 ( n15193,p3_u3897,n15195 );
   nand U14726 ( p3_u3520,n15196,n15197 );
   nand U14727 ( n15197,p3_datao_reg_29_,n15191 );
   nand U14728 ( n15196,p3_u3897,n15198 );
   nand U14729 ( p3_u3519,n15199,n15200 );
   nand U14730 ( n15200,p3_datao_reg_28_,n15191 );
   nand U14731 ( n15199,p3_u3897,n15201 );
   nand U14732 ( p3_u3518,n15202,n15203 );
   nand U14733 ( n15203,p3_datao_reg_27_,n15191 );
   nand U14734 ( n15202,p3_u3897,n15204 );
   nand U14735 ( p3_u3517,n15205,n15206 );
   nand U14736 ( n15206,p3_datao_reg_26_,n15191 );
   nand U14737 ( n15205,p3_u3897,n15207 );
   nand U14738 ( p3_u3516,n15208,n15209 );
   nand U14739 ( n15209,p3_datao_reg_25_,n15191 );
   nand U14740 ( n15208,p3_u3897,n15210 );
   nand U14741 ( p3_u3515,n15211,n15212 );
   nand U14742 ( n15212,p3_datao_reg_24_,n15191 );
   nand U14743 ( n15211,p3_u3897,n15213 );
   nand U14744 ( p3_u3514,n15214,n15215 );
   nand U14745 ( n15215,p3_datao_reg_23_,n15191 );
   nand U14746 ( n15214,p3_u3897,n15216 );
   nand U14747 ( p3_u3513,n15217,n15218 );
   nand U14748 ( n15218,p3_datao_reg_22_,n15191 );
   nand U14749 ( n15217,p3_u3897,n15219 );
   nand U14750 ( p3_u3512,n15220,n15221 );
   nand U14751 ( n15221,p3_datao_reg_21_,n15191 );
   nand U14752 ( n15220,p3_u3897,n15222 );
   nand U14753 ( p3_u3511,n15223,n15224 );
   nand U14754 ( n15224,p3_datao_reg_20_,n15191 );
   nand U14755 ( n15223,p3_u3897,n15225 );
   nand U14756 ( p3_u3510,n15226,n15227 );
   nand U14757 ( n15227,p3_datao_reg_19_,n15191 );
   nand U14758 ( n15226,p3_u3897,n15228 );
   nand U14759 ( p3_u3509,n15229,n15230 );
   nand U14760 ( n15230,p3_datao_reg_18_,n15191 );
   nand U14761 ( n15229,p3_u3897,n15231 );
   nand U14762 ( p3_u3508,n15232,n15233 );
   nand U14763 ( n15233,p3_datao_reg_17_,n15191 );
   nand U14764 ( n15232,p3_u3897,n15234 );
   nand U14765 ( p3_u3507,n15235,n15236 );
   nand U14766 ( n15236,p3_datao_reg_16_,n15191 );
   nand U14767 ( n15235,p3_u3897,n15237 );
   nand U14768 ( p3_u3506,n15238,n15239 );
   nand U14769 ( n15239,p3_datao_reg_15_,n15191 );
   nand U14770 ( n15238,p3_u3897,n15240 );
   nand U14771 ( p3_u3505,n15241,n15242 );
   nand U14772 ( n15242,p3_datao_reg_14_,n15191 );
   nand U14773 ( n15241,p3_u3897,n15243 );
   nand U14774 ( p3_u3504,n15244,n15245 );
   nand U14775 ( n15245,p3_datao_reg_13_,n15191 );
   nand U14776 ( n15244,p3_u3897,n15246 );
   nand U14777 ( p3_u3503,n15247,n15248 );
   nand U14778 ( n15248,p3_datao_reg_12_,n15191 );
   nand U14779 ( n15247,p3_u3897,n15249 );
   nand U14780 ( p3_u3502,n15250,n15251 );
   nand U14781 ( n15251,p3_datao_reg_11_,n15191 );
   nand U14782 ( n15250,p3_u3897,n15252 );
   nand U14783 ( p3_u3501,n15253,n15254 );
   nand U14784 ( n15254,p3_datao_reg_10_,n15191 );
   nand U14785 ( n15253,p3_u3897,n15255 );
   nand U14786 ( p3_u3500,n15256,n15257 );
   nand U14787 ( n15257,p3_datao_reg_9_,n15191 );
   nand U14788 ( n15256,p3_u3897,n15258 );
   nand U14789 ( p3_u3499,n15259,n15260 );
   nand U14790 ( n15260,p3_datao_reg_8_,n15191 );
   nand U14791 ( n15259,p3_u3897,n15261 );
   nand U14792 ( p3_u3498,n15262,n15263 );
   nand U14793 ( n15263,p3_datao_reg_7_,n15191 );
   nand U14794 ( n15262,p3_u3897,n15264 );
   nand U14795 ( p3_u3497,n15265,n15266 );
   nand U14796 ( n15266,p3_datao_reg_6_,n15191 );
   nand U14797 ( n15265,p3_u3897,n15267 );
   nand U14798 ( p3_u3496,n15268,n15269 );
   nand U14799 ( n15269,p3_datao_reg_5_,n15191 );
   nand U14800 ( n15268,p3_u3897,n15270 );
   nand U14801 ( p3_u3495,n15271,n15272 );
   nand U14802 ( n15272,p3_datao_reg_4_,n15191 );
   nand U14803 ( n15271,p3_u3897,n15273 );
   nand U14804 ( p3_u3494,n15274,n15275 );
   nand U14805 ( n15275,p3_datao_reg_3_,n15191 );
   nand U14806 ( n15274,p3_u3897,n15276 );
   nand U14807 ( p3_u3493,n15277,n15278 );
   nand U14808 ( n15278,p3_datao_reg_2_,n15191 );
   nand U14809 ( n15277,p3_u3897,n15279 );
   nand U14810 ( p3_u3492,n15280,n15281 );
   nand U14811 ( n15281,p3_datao_reg_1_,n15191 );
   nand U14812 ( n15280,p3_u3897,n15282 );
   nand U14813 ( p3_u3491,n15283,n15284 );
   nand U14814 ( n15284,p3_datao_reg_0_,n15191 );
   nand U14815 ( n15283,p3_u3897,n15285 );
   nand U14816 ( p3_u3490,n15286,n15287,n15288 );
   nand U14817 ( n15288,p3_reg1_reg_31_,n15289 );
   nand U14818 ( n15286,n15290,n15291 );
   nand U14819 ( p3_u3489,n15292,n15287,n15293 );
   nand U14820 ( n15293,p3_reg1_reg_30_,n15289 );
   nand U14821 ( n15287,n15294,n15295 );
   nand U14822 ( n15292,n15290,n15296 );
   nand U14823 ( p3_u3488,n15297,n15298,n15299,n15300 );
   nand U14824 ( n15300,p3_reg1_reg_29_,n15289 );
   nand U14825 ( n15299,n15295,n15301 );
   nand U14826 ( n15298,n15302,n15303 );
   nand U14827 ( n15297,n15290,n15304 );
   nand U14828 ( p3_u3487,n15305,n15306,n15307,n15308 );
   nand U14829 ( n15308,n15302,n15309 );
   nand U14830 ( n15307,n15310,n15198 );
   nand U14831 ( n15306,n15290,n15311 );
   nor U14832 ( n15305,n15312,n15313 );
   and U14833 ( n15313,n15289,p3_reg1_reg_28_ );
   nor U14834 ( n15312,n15314,n15289 );
   nand U14835 ( p3_u3486,n15315,n15316,n15317,n15318 );
   nand U14836 ( n15318,n15302,n15319 );
   nand U14837 ( n15317,n15310,n15201 );
   nand U14838 ( n15316,n15290,n15320 );
   nor U14839 ( n15315,n15321,n15322 );
   and U14840 ( n15322,n15289,p3_reg1_reg_27_ );
   nor U14841 ( n15321,n15323,n15289 );
   nand U14842 ( p3_u3485,n15324,n15325,n15326,n15327 );
   nand U14843 ( n15327,n15328,n15302 );
   nand U14844 ( n15326,n15310,n15204 );
   nand U14845 ( n15325,n15290,n15329 );
   nor U14846 ( n15324,n15330,n15331 );
   and U14847 ( n15331,n15289,p3_reg1_reg_26_ );
   and U14848 ( n15330,n15332,n15295 );
   nand U14849 ( p3_u3484,n15333,n15334,n15335 );
   nor U14850 ( n15335,n15336,n15337,n15338 );
   and U14851 ( n15338,n15289,p3_reg1_reg_25_ );
   nor U14852 ( n15337,n15339,n15289 );
   nor U14853 ( n15336,n15340,n15341 );
   nand U14854 ( n15334,n15342,n15302 );
   nand U14855 ( n15333,n15310,n15207 );
   nand U14856 ( p3_u3483,n15343,n15344,n15345 );
   nor U14857 ( n15345,n15346,n15347,n15348 );
   and U14858 ( n15348,n15289,p3_reg1_reg_24_ );
   nor U14859 ( n15347,n15349,n15289 );
   nor U14860 ( n15346,n15350,n15341 );
   nand U14861 ( n15344,n15351,n15302 );
   nand U14862 ( n15343,n15310,n15210 );
   nand U14863 ( p3_u3482,n15352,n15353,n15354,n15355 );
   nand U14864 ( n15355,n15302,n15356 );
   nand U14865 ( n15354,n15310,n15213 );
   nand U14866 ( n15353,n15290,n15357 );
   nor U14867 ( n15352,n15358,n15359 );
   and U14868 ( n15359,n15289,p3_reg1_reg_23_ );
   nor U14869 ( n15358,n15360,n15289 );
   nand U14870 ( p3_u3481,n15361,n15362,n15363,n15364 );
   nand U14871 ( n15364,p3_reg1_reg_22_,n15289 );
   nand U14872 ( n15363,n15295,n15365 );
   nand U14873 ( n15362,n15310,n15216 );
   nand U14874 ( n15361,n15290,n15366 );
   nand U14875 ( p3_u3480,n15367,n15368,n15369,n15370 );
   nand U14876 ( n15370,p3_reg1_reg_21_,n15289 );
   nand U14877 ( n15369,n15295,n15371 );
   nand U14878 ( n15368,n15310,n15219 );
   nand U14879 ( n15367,n15290,n15372 );
   nand U14880 ( p3_u3479,n15373,n15374,n15375 );
   nor U14881 ( n15375,n15376,n15377,n15378 );
   and U14882 ( n15378,n15289,p3_reg1_reg_20_ );
   nor U14883 ( n15377,n15379,n15289 );
   nor U14884 ( n15376,n15380,n15341 );
   nand U14885 ( n15374,n15381,n15302 );
   nand U14886 ( n15373,n15310,n15222 );
   nand U14887 ( p3_u3478,n15382,n15383,n15384,n15385 );
   nand U14888 ( n15385,n15386,n15302 );
   nand U14889 ( n15384,n15310,n15225 );
   nand U14890 ( n15383,n15290,n15387 );
   nor U14891 ( n15382,n15388,n15389 );
   and U14892 ( n15389,n15289,p3_reg1_reg_19_ );
   nor U14893 ( n15388,n15390,n15289 );
   nand U14894 ( p3_u3477,n15391,n15392,n15393,n15394 );
   nor U14895 ( n15394,n15395,n15396 );
   nor U14896 ( n15396,n15397,n15398 );
   nor U14897 ( n15395,n15399,n15400 );
   nand U14898 ( n15393,n15290,n15401 );
   nand U14899 ( n15392,n15295,n15402 );
   nand U14900 ( n15391,p3_reg1_reg_18_,n15289 );
   nand U14901 ( p3_u3476,n15403,n15404,n15405,n15406 );
   nor U14902 ( n15406,n15407,n15408 );
   nor U14903 ( n15408,n15409,n15398 );
   nor U14904 ( n15407,n15410,n15399 );
   nand U14905 ( n15405,n15290,n15411 );
   nand U14906 ( n15404,p3_reg1_reg_17_,n15289 );
   nand U14907 ( n15403,n15295,n15412 );
   nand U14908 ( p3_u3475,n15413,n15414,n15415,n15416 );
   nand U14909 ( n15416,n15302,n15417 );
   nand U14910 ( n15415,n15310,n15234 );
   nand U14911 ( n15414,n15290,n15418 );
   nor U14912 ( n15413,n15419,n15420 );
   nor U14913 ( n15420,n15295,n15421 );
   nor U14914 ( n15419,n15422,n15289 );
   nand U14915 ( p3_u3474,n15423,n15424,n15425,n15426 );
   nand U14916 ( n15426,p3_reg1_reg_15_,n15289 );
   nand U14917 ( n15425,n15295,n15427 );
   nand U14918 ( n15424,n15310,n15237 );
   nand U14919 ( n15423,n15290,n15428 );
   nand U14920 ( p3_u3473,n15429,n15430,n15431,n15432 );
   nor U14921 ( n15432,n15433,n15434 );
   nor U14922 ( n15434,n15435,n15398 );
   nor U14923 ( n15433,n15436,n15399 );
   nand U14924 ( n15431,n15290,n15437 );
   nand U14925 ( n15430,p3_reg1_reg_14_,n15289 );
   nand U14926 ( n15429,n15295,n15438 );
   nand U14927 ( p3_u3472,n15439,n15440,n15441,n15442 );
   nand U14928 ( n15442,n15443,n15302 );
   nand U14929 ( n15441,n15310,n15243 );
   nand U14930 ( n15440,n15290,n15444 );
   nor U14931 ( n15439,n15445,n15446 );
   nor U14932 ( n15446,n15295,n15447 );
   nor U14933 ( n15445,n15448,n15289 );
   nand U14934 ( p3_u3471,n15449,n15450,n15451,n15452 );
   nand U14935 ( n15452,n15302,n15453 );
   nand U14936 ( n15451,n15310,n15246 );
   nand U14937 ( n15450,n15290,n15454 );
   nor U14938 ( n15449,n15455,n15456 );
   nor U14939 ( n15456,n15295,n15457 );
   nor U14940 ( n15455,n15458,n15289 );
   nand U14941 ( p3_u3470,n15459,n15460,n15461,n15462 );
   nand U14942 ( n15462,n15302,n15463 );
   nand U14943 ( n15461,n15310,n15249 );
   nand U14944 ( n15460,n15290,n15464 );
   nor U14945 ( n15459,n15465,n15466 );
   nor U14946 ( n15466,n15295,n15467 );
   nor U14947 ( n15465,n15468,n15289 );
   nand U14948 ( p3_u3469,n15469,n15470,n15471,n15472 );
   nand U14949 ( n15472,p3_reg1_reg_10_,n15289 );
   nand U14950 ( n15471,n15295,n15473 );
   nand U14951 ( n15470,n15310,n15252 );
   nand U14952 ( n15469,n15290,n15474 );
   nand U14953 ( p3_u3468,n15475,n15476,n15477,n15478 );
   nand U14954 ( n15478,p3_reg1_reg_9_,n15289 );
   nand U14955 ( n15477,n15295,n15479 );
   nand U14956 ( n15476,n15310,n15255 );
   nand U14957 ( n15475,n15290,n15480 );
   nand U14958 ( p3_u3467,n15481,n15482,n15483,n15484 );
   nor U14959 ( n15484,n15485,n15486 );
   nor U14960 ( n15486,n15487,n15398 );
   nor U14961 ( n15485,n15488,n15399 );
   nand U14962 ( n15483,n15290,n15489 );
   nand U14963 ( n15482,p3_reg1_reg_8_,n15289 );
   nand U14964 ( n15481,n15295,n15490 );
   nand U14965 ( p3_u3466,n15491,n15492,n15493,n15494 );
   nand U14966 ( n15494,n15495,n15302 );
   nand U14967 ( n15493,n15310,n15261 );
   nand U14968 ( n15492,n15290,n15496 );
   nor U14969 ( n15491,n15497,n15498 );
   nor U14970 ( n15498,n15295,n15499 );
   nor U14971 ( n15497,n15500,n15289 );
   nand U14972 ( p3_u3465,n15501,n15502,n15503,n15504 );
   nor U14973 ( n15504,n15505,n15506 );
   nor U14974 ( n15506,n15507,n15398 );
   nor U14975 ( n15505,n15508,n15399 );
   nand U14976 ( n15503,n15290,n15509 );
   nand U14977 ( n15502,n15295,n15510 );
   nand U14978 ( n15501,p3_reg1_reg_6_,n15289 );
   nand U14979 ( p3_u3464,n15511,n15512,n15513,n15514 );
   nand U14980 ( n15514,p3_reg1_reg_5_,n15289 );
   nand U14981 ( n15513,n15295,n15515 );
   nand U14982 ( n15512,n15310,n15267 );
   nand U14983 ( n15511,n15290,n15516 );
   nand U14984 ( p3_u3463,n15517,n15518,n15519,n15520 );
   nand U14985 ( n15520,p3_reg1_reg_4_,n15289 );
   nand U14986 ( n15519,n15295,n15521 );
   nand U14987 ( n15518,n15310,n15270 );
   nand U14988 ( n15517,n15290,n15522 );
   nand U14989 ( p3_u3462,n15523,n15524,n15525,n15526 );
   nand U14990 ( n15526,n15302,n15527 );
   nand U14991 ( n15525,n15310,n15273 );
   nand U14992 ( n15524,n15290,n15528 );
   nor U14993 ( n15523,n15529,n15530 );
   nor U14994 ( n15530,n15295,n15531 );
   nor U14995 ( n15529,n15532,n15289 );
   nand U14996 ( p3_u3461,n15533,n15534,n15535,n15536 );
   or U14997 ( n15536,n15537,n15399 );
   nand U14998 ( n15535,n15310,n15276 );
   nand U14999 ( n15534,n15290,n15538 );
   nor U15000 ( n15533,n15539,n15540 );
   and U15001 ( n15540,n15541,n15295 );
   nor U15002 ( n15539,n15295,n15542 );
   nand U15003 ( p3_u3460,n15543,n15544,n15545,n15546 );
   nand U15004 ( n15546,n15302,n15547 );
   nand U15005 ( n15545,n15310,n15279 );
   nand U15006 ( n15544,n15290,n15548 );
   nor U15007 ( n15543,n15549,n15550 );
   nor U15008 ( n15550,n15295,n15551 );
   nor U15009 ( n15549,n15552,n15289 );
   nand U15010 ( p3_u3459,n15553,n15554,n15555,n15556 );
   nand U15011 ( n15556,n15302,n15557 );
   not U15012 ( n15302,n15399 );
   nand U15013 ( n15399,n15558,n15295 );
   nand U15014 ( n15555,n15310,n15282 );
   nand U15015 ( n15398,n15559,n15560,n15295 );
   nand U15016 ( n15554,n15290,n15561 );
   nand U15017 ( n15341,n15295,n15562 );
   nor U15018 ( n15553,n15563,n15564 );
   and U15019 ( n15564,n15565,n15295 );
   and U15020 ( n15563,n15289,p3_reg1_reg_0_ );
   nand U15021 ( n15569,n15570,n15571 );
   nand U15022 ( n15571,n15572,n15573 );
   nand U15023 ( n15573,n15574,n15575,n15576 );
   nand U15024 ( n15575,n15577,n15578 );
   nand U15025 ( n15574,n15579,n15580 );
   nand U15026 ( n15568,n15581,n15582 );
   nand U15027 ( n15581,n15583,n15584 );
   nand U15028 ( p3_u3458,n15585,n15586,n15587 );
   nand U15029 ( n15587,n15588,p3_reg0_reg_31_ );
   nand U15030 ( n15585,n15589,n15291 );
   nand U15031 ( p3_u3457,n15590,n15586,n15591 );
   nand U15032 ( n15591,n15588,p3_reg0_reg_30_ );
   nand U15033 ( n15586,n15294,n15592 );
   nand U15034 ( n15590,n15589,n15296 );
   nand U15035 ( p3_u3456,n15593,n15594,n15595,n15596 );
   nand U15036 ( n15596,n15588,p3_reg0_reg_29_ );
   nand U15037 ( n15595,n15592,n15301 );
   nand U15038 ( n15594,n15597,n15303 );
   nand U15039 ( n15593,n15589,n15304 );
   nand U15040 ( p3_u3455,n15598,n15599,n15600,n15601 );
   nand U15041 ( n15601,n15597,n15309 );
   nand U15042 ( n15600,n15602,n15198 );
   nand U15043 ( n15599,n15589,n15311 );
   nor U15044 ( n15598,n15603,n15604 );
   nor U15045 ( n15604,n15314,n15588 );
   and U15046 ( n15603,p3_reg0_reg_28_,n15588 );
   nand U15047 ( p3_u3454,n15605,n15606,n15607,n15608 );
   nand U15048 ( n15608,n15597,n15319 );
   nand U15049 ( n15607,n15602,n15201 );
   nand U15050 ( n15606,n15589,n15320 );
   nor U15051 ( n15605,n15609,n15610 );
   nor U15052 ( n15610,n15323,n15588 );
   and U15053 ( n15609,p3_reg0_reg_27_,n15588 );
   nand U15054 ( p3_u3453,n15611,n15612,n15613,n15614 );
   nor U15055 ( n15614,n15615,n15616 );
   nor U15056 ( n15616,n15617,n15618 );
   nor U15057 ( n15615,n15619,n15620 );
   nand U15058 ( n15613,n15589,n15329 );
   nand U15059 ( n15612,n15588,p3_reg0_reg_26_ );
   nand U15060 ( n15611,n15592,n15332 );
   nand U15061 ( p3_u3452,n15621,n15622,n15623,n15624 );
   nand U15062 ( n15624,n15597,n15342 );
   nand U15063 ( n15623,n15602,n15207 );
   nand U15064 ( n15622,n15589,n15625 );
   nor U15065 ( n15621,n15626,n15627 );
   nor U15066 ( n15627,n15339,n15588 );
   and U15067 ( n15626,p3_reg0_reg_25_,n15588 );
   nand U15068 ( p3_u3451,n15628,n15629,n15630,n15631 );
   nand U15069 ( n15631,n15597,n15351 );
   nand U15070 ( n15630,n15602,n15210 );
   nand U15071 ( n15629,n15589,n15632 );
   nor U15072 ( n15628,n15633,n15634 );
   nor U15073 ( n15634,n15349,n15588 );
   and U15074 ( n15633,p3_reg0_reg_24_,n15588 );
   nand U15075 ( p3_u3450,n15635,n15636,n15637,n15638 );
   nand U15076 ( n15638,n15597,n15356 );
   nand U15077 ( n15637,n15602,n15213 );
   nand U15078 ( n15636,n15589,n15357 );
   nor U15079 ( n15635,n15639,n15640 );
   nor U15080 ( n15640,n15360,n15588 );
   and U15081 ( n15639,p3_reg0_reg_23_,n15588 );
   nand U15082 ( p3_u3449,n15641,n15642,n15643,n15644 );
   nand U15083 ( n15644,n15588,p3_reg0_reg_22_ );
   nand U15084 ( n15643,n15592,n15365 );
   nand U15085 ( n15365,n15645,n15646 );
   nand U15086 ( n15646,n15558,n15647 );
   not U15087 ( n15645,n15648 );
   nand U15088 ( n15642,n15602,n15216 );
   nand U15089 ( n15641,n15589,n15366 );
   nand U15090 ( p3_u3448,n15649,n15650,n15651,n15652 );
   nand U15091 ( n15652,n15588,p3_reg0_reg_21_ );
   nand U15092 ( n15651,n15592,n15371 );
   nand U15093 ( n15371,n15653,n15654 );
   nand U15094 ( n15654,n15558,n15655 );
   not U15095 ( n15653,n15656 );
   nand U15096 ( n15650,n15602,n15219 );
   nand U15097 ( n15649,n15589,n15372 );
   nand U15098 ( p3_u3447,n15657,n15658,n15659,n15660 );
   nand U15099 ( n15660,n15597,n15381 );
   nand U15100 ( n15659,n15602,n15222 );
   nand U15101 ( n15658,n15589,n15661 );
   nor U15102 ( n15657,n15662,n15663 );
   nor U15103 ( n15663,n15379,n15588 );
   and U15104 ( n15662,p3_reg0_reg_20_,n15588 );
   nand U15105 ( p3_u3446,n15664,n15665,n15666,n15667 );
   nand U15106 ( n15667,n15597,n15386 );
   nand U15107 ( n15666,n15602,n15225 );
   nand U15108 ( n15665,n15589,n15387 );
   nor U15109 ( n15664,n15668,n15669 );
   nor U15110 ( n15669,n15390,n15588 );
   and U15111 ( n15668,p3_reg0_reg_19_,n15588 );
   nand U15112 ( p3_u3444,n15670,n15671,n15672,n15673 );
   nor U15113 ( n15673,n15674,n15675 );
   nor U15114 ( n15675,n15397,n15618 );
   nor U15115 ( n15674,n15400,n15620 );
   nand U15116 ( n15672,n15589,n15401 );
   nand U15117 ( n15671,n15588,p3_reg0_reg_18_ );
   nand U15118 ( n15670,n15592,n15402 );
   nand U15119 ( p3_u3441,n15676,n15677,n15678,n15679 );
   nor U15120 ( n15679,n15680,n15681 );
   nor U15121 ( n15681,n15409,n15618 );
   nor U15122 ( n15680,n15410,n15620 );
   nand U15123 ( n15678,n15589,n15411 );
   nand U15124 ( n15677,n15588,p3_reg0_reg_17_ );
   nand U15125 ( n15676,n15592,n15412 );
   nand U15126 ( p3_u3438,n15682,n15683,n15684,n15685 );
   nand U15127 ( n15685,n15597,n15417 );
   nand U15128 ( n15684,n15602,n15234 );
   nand U15129 ( n15683,n15589,n15418 );
   nor U15130 ( n15682,n15686,n15687 );
   nor U15131 ( n15687,n15422,n15588 );
   and U15132 ( n15686,p3_reg0_reg_16_,n15588 );
   nand U15133 ( p3_u3435,n15688,n15689,n15690,n15691 );
   nand U15134 ( n15691,n15588,p3_reg0_reg_15_ );
   nand U15135 ( n15690,n15592,n15427 );
   nand U15136 ( n15427,n15692,n15693 );
   nand U15137 ( n15693,n15558,n15694 );
   not U15138 ( n15692,n15695 );
   nand U15139 ( n15689,n15602,n15237 );
   nand U15140 ( n15688,n15589,n15428 );
   nand U15141 ( p3_u3432,n15696,n15697,n15698,n15699 );
   nor U15142 ( n15699,n15700,n15701 );
   nor U15143 ( n15701,n15435,n15618 );
   nor U15144 ( n15700,n15436,n15620 );
   nand U15145 ( n15698,n15589,n15437 );
   nand U15146 ( n15697,n15588,p3_reg0_reg_14_ );
   nand U15147 ( n15696,n15592,n15438 );
   nand U15148 ( p3_u3429,n15702,n15703,n15704,n15705 );
   nand U15149 ( n15705,n15597,n15443 );
   nand U15150 ( n15704,n15602,n15243 );
   nand U15151 ( n15703,n15589,n15444 );
   nor U15152 ( n15702,n15706,n15707 );
   nor U15153 ( n15707,n15448,n15588 );
   and U15154 ( n15706,p3_reg0_reg_13_,n15588 );
   nand U15155 ( p3_u3426,n15708,n15709,n15710,n15711 );
   nand U15156 ( n15711,n15597,n15453 );
   nand U15157 ( n15710,n15602,n15246 );
   nand U15158 ( n15709,n15589,n15454 );
   nor U15159 ( n15708,n15712,n15713 );
   nor U15160 ( n15713,n15458,n15588 );
   and U15161 ( n15712,p3_reg0_reg_12_,n15588 );
   nand U15162 ( p3_u3423,n15714,n15715,n15716,n15717 );
   nand U15163 ( n15717,n15597,n15463 );
   nand U15164 ( n15716,n15602,n15249 );
   nand U15165 ( n15715,n15589,n15464 );
   nor U15166 ( n15714,n15718,n15719 );
   nor U15167 ( n15719,n15468,n15588 );
   and U15168 ( n15718,p3_reg0_reg_11_,n15588 );
   nand U15169 ( p3_u3420,n15720,n15721,n15722,n15723 );
   nand U15170 ( n15723,n15588,p3_reg0_reg_10_ );
   nand U15171 ( n15722,n15592,n15473 );
   nand U15172 ( n15473,n15724,n15725 );
   nand U15173 ( n15725,n15558,n15726 );
   not U15174 ( n15724,n15727 );
   nand U15175 ( n15721,n15602,n15252 );
   nand U15176 ( n15720,n15589,n15474 );
   nand U15177 ( p3_u3417,n15728,n15729,n15730,n15731 );
   nand U15178 ( n15731,n15588,p3_reg0_reg_9_ );
   nand U15179 ( n15730,n15592,n15479 );
   nand U15180 ( n15479,n15732,n15733 );
   nand U15181 ( n15733,n15558,n15734 );
   not U15182 ( n15732,n15735 );
   nand U15183 ( n15729,n15602,n15255 );
   nand U15184 ( n15728,n15589,n15480 );
   nand U15185 ( p3_u3414,n15736,n15737,n15738,n15739 );
   nor U15186 ( n15739,n15740,n15741 );
   nor U15187 ( n15741,n15487,n15618 );
   nor U15188 ( n15740,n15488,n15620 );
   nand U15189 ( n15738,n15589,n15489 );
   nand U15190 ( n15737,n15588,p3_reg0_reg_8_ );
   nand U15191 ( n15736,n15592,n15490 );
   nand U15192 ( p3_u3411,n15742,n15743,n15744,n15745 );
   nand U15193 ( n15745,n15597,n15495 );
   nand U15194 ( n15744,n15602,n15261 );
   nand U15195 ( n15743,n15589,n15496 );
   nor U15196 ( n15742,n15746,n15747 );
   nor U15197 ( n15747,n15500,n15588 );
   not U15198 ( n15500,n15748 );
   and U15199 ( n15746,p3_reg0_reg_7_,n15588 );
   nand U15200 ( p3_u3408,n15749,n15750,n15751,n15752 );
   nor U15201 ( n15752,n15753,n15754 );
   nor U15202 ( n15754,n15507,n15618 );
   nor U15203 ( n15753,n15508,n15620 );
   nand U15204 ( n15751,n15589,n15509 );
   nand U15205 ( n15750,n15588,p3_reg0_reg_6_ );
   nand U15206 ( n15749,n15592,n15510 );
   nand U15207 ( p3_u3405,n15755,n15756,n15757,n15758 );
   nand U15208 ( n15758,n15588,p3_reg0_reg_5_ );
   nand U15209 ( n15757,n15592,n15515 );
   nand U15210 ( n15515,n15759,n15760 );
   nand U15211 ( n15760,n15558,n15761 );
   not U15212 ( n15759,n15762 );
   nand U15213 ( n15756,n15602,n15267 );
   nand U15214 ( n15755,n15589,n15516 );
   nand U15215 ( p3_u3402,n15763,n15764,n15765,n15766 );
   nand U15216 ( n15766,n15588,p3_reg0_reg_4_ );
   nand U15217 ( n15765,n15592,n15521 );
   nand U15218 ( n15521,n15767,n15768 );
   nand U15219 ( n15768,n15558,n15769 );
   not U15220 ( n15767,n15770 );
   nand U15221 ( n15764,n15602,n15270 );
   nand U15222 ( n15763,n15589,n15522 );
   nand U15223 ( p3_u3399,n15771,n15772,n15773,n15774 );
   nand U15224 ( n15774,n15597,n15527 );
   nand U15225 ( n15773,n15602,n15273 );
   nand U15226 ( n15772,n15589,n15528 );
   nor U15227 ( n15771,n15775,n15776 );
   nor U15228 ( n15776,n15532,n15588 );
   and U15229 ( n15775,p3_reg0_reg_3_,n15588 );
   nand U15230 ( p3_u3396,n15777,n15778,n15779,n15780 );
   nor U15231 ( n15780,n15781,n15782 );
   nor U15232 ( n15782,n15783,n15618 );
   nor U15233 ( n15781,n15537,n15620 );
   nand U15234 ( n15779,n15589,n15538 );
   nand U15235 ( n15778,n15588,p3_reg0_reg_2_ );
   nand U15236 ( n15777,n15592,n15541 );
   nand U15237 ( p3_u3393,n15784,n15785,n15786,n15787 );
   nand U15238 ( n15787,n15597,n15547 );
   not U15239 ( n15597,n15620 );
   nand U15240 ( n15786,n15602,n15279 );
   nand U15241 ( n15785,n15589,n15548 );
   nor U15242 ( n15784,n15788,n15789 );
   nor U15243 ( n15789,n15552,n15588 );
   and U15244 ( n15788,p3_reg0_reg_1_,n15588 );
   nand U15245 ( p3_u3390,n15790,n15791,n15792,n15793 );
   nor U15246 ( n15793,n15794,n15795 );
   nor U15247 ( n15795,n15796,n15618 );
   nand U15248 ( n15618,n15592,n15560,n15559 );
   nor U15249 ( n15794,n15797,n15620 );
   nand U15250 ( n15620,n15558,n15592 );
   nand U15251 ( n15792,n15589,n15561 );
   nand U15252 ( n15791,n15588,p3_reg0_reg_0_ );
   nand U15253 ( n15790,n15592,n15565 );
   nand U15254 ( n15799,n15567,n15800 );
   nand U15255 ( n15800,n15801,n15802 );
   nand U15256 ( n15802,n15803,n15804 );
   nand U15257 ( n15801,n15805,n15806 );
   nand U15258 ( n15806,n15807,n15808 );
   nand U15259 ( n15808,n15577,n15809 );
   xor U15260 ( n15807,n15579,n15580 );
   nand U15261 ( n15798,n15810,n15804 );
   nand U15262 ( p3_u3377,n15811,n15812 );
   nand U15263 ( n15812,p3_d_reg_1_,n15813 );
   nand U15264 ( n15811,n15814,n15815 );
   nand U15265 ( p3_u3376,n15816,n15817 );
   nand U15266 ( n15817,p3_d_reg_0_,n15813 );
   nand U15267 ( n15816,n15814,n15818 );
   nor U15268 ( p3_u3296,n15819,n15820 );
   nor U15269 ( n15820,n15821,n15822 );
   not U15270 ( n15822,n15823 );
   nor U15271 ( n15821,p3_u3151,n15824 );
   nor U15272 ( n15819,n15825,n15826,n15827 );
   nor U15273 ( n15827,n15828,n15829 );
   nor U15274 ( n15826,n15830,n15831 );
   not U15275 ( n15830,n15829 );
   nand U15276 ( n15829,n15832,n15833 );
   nand U15277 ( n15833,n15834,n15291 );
   nand U15278 ( n15834,n15192,n15835 );
   nand U15279 ( n15832,n15836,n15837,n15838 );
   nand U15280 ( n15837,n15839,n15296 );
   nand U15281 ( n15836,n15840,n15841 );
   nand U15282 ( n15841,n15842,n15843 );
   nand U15283 ( n15843,n15844,n15304 );
   nand U15284 ( n15842,n15845,n15846 );
   nand U15285 ( n15846,n15847,n15848,n15849 );
   nand U15286 ( n15849,n15850,n15851,n15852 );
   nand U15287 ( n15850,n15853,n15854,n15855,n15856 );
   nand U15288 ( n15854,n15857,n15858 );
   nand U15289 ( n15857,n15859,n15860 );
   nand U15290 ( n15860,n15861,n15862 );
   not U15291 ( n15861,n15863 );
   nand U15292 ( n15853,n15864,n15865,n15866 );
   and U15293 ( n15866,n15867,n15858,n15862 );
   or U15294 ( n15867,n15868,n15869,n15870,n15871 );
   nor U15295 ( n15871,n15380,n15225 );
   nor U15296 ( n15870,n15872,n15873,n15234 );
   nor U15297 ( n15869,n15874,n15228 );
   nand U15298 ( n15868,n15875,n15876,n15877,n15878 );
   nand U15299 ( n15876,n15879,n15880,n15881,n15882 );
   nand U15300 ( n15882,n15883,n15884 );
   nand U15301 ( n15884,n15885,n15886 );
   nand U15302 ( n15885,n15887,n15888 );
   nand U15303 ( n15888,n15889,n15890 );
   nand U15304 ( n15889,n15891,n15892,n15893,n15894 );
   nand U15305 ( n15893,n15895,n15896,n15897,n15898 );
   nand U15306 ( n15896,n15899,n15900,n15901 );
   nand U15307 ( n15901,n15902,n15903 );
   nand U15308 ( n15903,n15904,n15261 );
   nand U15309 ( n15902,n15905,n15906,n15907 );
   nand U15310 ( n15907,n15908,n15489 );
   nand U15311 ( n15905,n15909,n15910 );
   nand U15312 ( n15909,n15911,n15912,n15913 );
   nand U15313 ( n15913,n15914,n15915 );
   nand U15314 ( n15911,n15916,n15917 );
   not U15315 ( n15895,n15918 );
   nand U15316 ( n15892,n15919,n15897 );
   nand U15317 ( n15919,n15920,n15921 );
   nand U15318 ( n15921,n15922,n15898 );
   not U15319 ( n15922,n15923 );
   nand U15320 ( n15880,n15873,n15234 );
   not U15321 ( n15879,n15872 );
   nand U15322 ( n15872,n15924,n15925 );
   nand U15323 ( n15925,n15926,n15231 );
   nand U15324 ( n15875,n15924,n15401,n15409 );
   nand U15325 ( n15865,n15927,n15878 );
   nand U15326 ( n15927,n15928,n15929 );
   nand U15327 ( n15929,n15225,n15877,n15380 );
   nand U15328 ( n15840,n15930,n15198 );
   nand U15329 ( n15825,n15931,n15932,n15823 );
   nand U15330 ( n15823,p3_b_reg,n15933 );
   nand U15331 ( n15933,n15934,n15935,p3_state_reg );
   nand U15332 ( n15935,n15936,n15824 );
   nand U15333 ( n15936,n15937,n15938,n15939,n15940 );
   nor U15334 ( n15940,n15941,n15942 );
   nand U15335 ( n15934,n15943,n15944 );
   nand U15336 ( n15932,n15945,n15946 );
   xor U15337 ( n15945,n15947,n15948 );
   nand U15338 ( n15948,n15949,n15950,n15951 );
   nand U15339 ( n15951,n15952,n15953 );
   nand U15340 ( n15953,n15954,n15955,n15956,n15957 );
   nand U15341 ( n15957,n15958,n15959 );
   nand U15342 ( n15959,n15960,n15961 );
   nand U15343 ( n15961,n15962,n15963 );
   nand U15344 ( n15960,n15964,n15965 );
   not U15345 ( n15958,n15966 );
   nand U15346 ( n15956,n15967,n15968 );
   or U15347 ( n15967,n15969,n15970 );
   nand U15348 ( n15955,n15970,n15969 );
   nand U15349 ( n15969,n15971,n15972 );
   nand U15350 ( n15972,n15973,n15974,n15975 );
   nand U15351 ( n15971,n15976,n15977 );
   nand U15352 ( n15954,n15978,n15979 );
   not U15353 ( n15952,n15980 );
   nand U15354 ( n15950,n15981,n15982,n15983,n15984 );
   nor U15355 ( n15984,n15980,n15985,n15966 );
   nand U15356 ( n15966,n15986,n15987,n15988,n15974 );
   or U15357 ( n15974,n15977,n15976 );
   and U15358 ( n15976,n15989,n15990 );
   nand U15359 ( n15990,n15991,n15311 );
   nand U15360 ( n15989,n15992,n15201 );
   nand U15361 ( n15977,n15993,n15994 );
   nand U15362 ( n15994,n15311,n15992 );
   nand U15363 ( n15993,n15201,n15991 );
   or U15364 ( n15988,n15965,n15964 );
   and U15365 ( n15964,n15995,n15996 );
   nand U15366 ( n15996,n15991,n15329 );
   nand U15367 ( n15995,n15992,n15207 );
   nand U15368 ( n15965,n15997,n15998 );
   nand U15369 ( n15998,n15329,n15992 );
   nand U15370 ( n15997,n15207,n15991 );
   or U15371 ( n15987,n15973,n15975 );
   and U15372 ( n15975,n15999,n16000 );
   nand U15373 ( n16000,n15991,n15320 );
   nand U15374 ( n15999,n15992,n15204 );
   nand U15375 ( n15973,n16001,n16002 );
   nand U15376 ( n16002,n15991,n15204 );
   nand U15377 ( n16001,n15992,n15320 );
   or U15378 ( n15986,n15968,n15970 );
   and U15379 ( n15970,n16003,n16004 );
   nand U15380 ( n16004,n15991,n15304 );
   nand U15381 ( n16003,n15992,n15198 );
   nand U15382 ( n15968,n16005,n16006 );
   nand U15383 ( n16006,n15991,n15198 );
   nand U15384 ( n16005,n15992,n15304 );
   nor U15385 ( n15985,n15962,n15963 );
   nand U15386 ( n15963,n16007,n16008 );
   nand U15387 ( n16008,n15991,n15210 );
   nand U15388 ( n16007,n15992,n15625 );
   and U15389 ( n15962,n16009,n16010 );
   nand U15390 ( n16010,n15991,n15625 );
   nand U15391 ( n16009,n15992,n15210 );
   nand U15392 ( n15980,n16011,n16012 );
   or U15393 ( n16012,n15979,n15978 );
   and U15394 ( n15978,n16013,n16014 );
   nand U15395 ( n16014,n15991,n15296 );
   nand U15396 ( n16013,n15992,n15195 );
   nand U15397 ( n15979,n16015,n16016 );
   nand U15398 ( n16016,n15991,n15195 );
   nand U15399 ( n16015,n15992,n15296 );
   nand U15400 ( n16011,n16017,n16018 );
   nand U15401 ( n15983,n16019,n16020 );
   nand U15402 ( n15982,n16021,n16022,n16023 );
   not U15403 ( n16022,n16024 );
   nand U15404 ( n16021,n16025,n16026 );
   nand U15405 ( n16026,n16027,n16028 );
   or U15406 ( n16025,n16029,n16030 );
   nand U15407 ( n15981,n16023,n16031,n16032,n16033 );
   nor U15408 ( n16033,n16034,n16035,n16024 );
   nor U15409 ( n16024,n16020,n16019 );
   and U15410 ( n16019,n16036,n16037 );
   nand U15411 ( n16037,n15991,n15213 );
   nand U15412 ( n16036,n15992,n15632 );
   nand U15413 ( n16020,n16038,n16039 );
   nand U15414 ( n16039,n15991,n15632 );
   nand U15415 ( n16038,n15992,n15213 );
   nor U15416 ( n16035,n16040,n16041 );
   nor U15417 ( n16034,n16042,n16043 );
   nor U15418 ( n16043,n16044,n16045 );
   nor U15419 ( n16045,n16046,n16047 );
   nor U15420 ( n16044,n16048,n16049,n16050 );
   not U15421 ( n16049,n16051 );
   not U15422 ( n16042,n16052 );
   nand U15423 ( n16032,n16051,n16052,n16053,n16054 );
   nor U15424 ( n16054,n16055,n16056 );
   nor U15425 ( n16056,n16057,n16058 );
   and U15426 ( n16055,n16048,n16050 );
   and U15427 ( n16050,n16059,n16060 );
   nand U15428 ( n16060,n15991,n15228 );
   nand U15429 ( n16059,n15992,n15387 );
   nand U15430 ( n16048,n16061,n16062 );
   nand U15431 ( n16062,n15991,n15387 );
   nand U15432 ( n16061,n15992,n15228 );
   nand U15433 ( n16053,n16063,n16064 );
   nand U15434 ( n16064,n16058,n16057 );
   nand U15435 ( n16057,n16065,n16066 );
   nand U15436 ( n16066,n16067,n16068,n16069 );
   not U15437 ( n16069,n16070 );
   nand U15438 ( n16065,n16071,n16072 );
   nand U15439 ( n16072,n16070,n16073 );
   nand U15440 ( n16073,n16067,n16068 );
   nand U15441 ( n16068,n16074,n16075,n16076 );
   nand U15442 ( n16076,n16077,n16078 );
   nand U15443 ( n16075,n16079,n16080,n16081 );
   or U15444 ( n16081,n16082,n16083 );
   nand U15445 ( n16080,n15991,n15428 );
   nand U15446 ( n16079,n15992,n15240 );
   nand U15447 ( n16074,n16083,n16082 );
   nand U15448 ( n16082,n16084,n16085 );
   nand U15449 ( n16085,n15991,n15240 );
   nand U15450 ( n16084,n15992,n15428 );
   nand U15451 ( n16083,n16086,n16087 );
   nand U15452 ( n16087,n16088,n16089 );
   nand U15453 ( n16089,n16090,n16091 );
   nand U15454 ( n16088,n16092,n16093 );
   nand U15455 ( n16093,n16094,n16095,n16096,n16097 );
   nand U15456 ( n16097,n16098,n16099 );
   nand U15457 ( n16096,n16100,n16101,n16102 );
   nand U15458 ( n16095,n16103,n16101,n16104 );
   or U15459 ( n16104,n16100,n16102 );
   and U15460 ( n16102,n16105,n16106 );
   nand U15461 ( n16106,n15991,n15252 );
   nand U15462 ( n16105,n15992,n15464 );
   nand U15463 ( n16100,n16107,n16108 );
   nand U15464 ( n16108,n15991,n15464 );
   nand U15465 ( n16107,n15992,n15252 );
   or U15466 ( n16101,n16099,n16098 );
   and U15467 ( n16098,n16109,n16110 );
   nand U15468 ( n16110,n15991,n15249 );
   nand U15469 ( n16109,n15992,n15454 );
   nand U15470 ( n16099,n16111,n16112 );
   nand U15471 ( n16112,n15991,n15454 );
   nand U15472 ( n16111,n15992,n15249 );
   nand U15473 ( n16103,n16113,n16114 );
   nand U15474 ( n16114,n16115,n16116,n16117 );
   nand U15475 ( n16117,n16118,n16119 );
   nand U15476 ( n16116,n16120,n16121,n16122 );
   not U15477 ( n16122,n16123 );
   nand U15478 ( n16115,n16124,n16125 );
   nand U15479 ( n16125,n16123,n16126 );
   nand U15480 ( n16126,n16120,n16121 );
   nand U15481 ( n16121,n16127,n16128,n16129 );
   nand U15482 ( n16129,n16130,n16131 );
   nand U15483 ( n16128,n16132,n16133,n16134,n16135 );
   nor U15484 ( n16135,n16136,n16137 );
   nor U15485 ( n16137,n16138,n16139 );
   nor U15486 ( n16136,n16130,n16131 );
   nand U15487 ( n16131,n16140,n16141 );
   nand U15488 ( n16141,n15991,n15264 );
   nand U15489 ( n16140,n15992,n15496 );
   and U15490 ( n16130,n16142,n16143 );
   nand U15491 ( n16143,n15991,n15496 );
   nand U15492 ( n16142,n15992,n15264 );
   nand U15493 ( n16134,n16144,n16145,n16146 );
   nand U15494 ( n16133,n16144,n16147,n16148,n16149 );
   nand U15495 ( n16149,n16150,n16151,n16152 );
   nand U15496 ( n16152,n16153,n16154 );
   nand U15497 ( n16151,n16155,n16156,n16157 );
   nand U15498 ( n16157,n16158,n16159 );
   nand U15499 ( n16156,n16160,n16161 );
   or U15500 ( n16161,n16159,n16158 );
   and U15501 ( n16158,n16162,n16163 );
   nand U15502 ( n16163,n15991,n15548 );
   nand U15503 ( n16162,n15992,n15282 );
   nand U15504 ( n16159,n16164,n16165 );
   nand U15505 ( n16165,n15991,n15282 );
   nand U15506 ( n16164,n15992,n15548 );
   nand U15507 ( n16160,n16166,n16167 );
   nand U15508 ( n16167,n16168,n16169,n16170 );
   nand U15509 ( n16169,n15285,n15992 );
   or U15510 ( n16168,n16171,n16172 );
   nand U15511 ( n16166,n16171,n16172 );
   nand U15512 ( n16171,n16173,n16174 );
   nand U15513 ( n16174,n15991,n15285 );
   nand U15514 ( n16173,n15992,n15561 );
   nand U15515 ( n16155,n16175,n16176 );
   or U15516 ( n16150,n16176,n16175 );
   and U15517 ( n16175,n16177,n16178 );
   nand U15518 ( n16178,n15991,n15538 );
   nand U15519 ( n16177,n15992,n15279 );
   nand U15520 ( n16176,n16179,n16180 );
   nand U15521 ( n16180,n15991,n15279 );
   nand U15522 ( n16179,n15992,n15538 );
   or U15523 ( n16148,n16154,n16153 );
   and U15524 ( n16153,n16181,n16182 );
   nand U15525 ( n16182,n15991,n15276 );
   nand U15526 ( n16181,n15992,n15528 );
   nand U15527 ( n16154,n16183,n16184 );
   nand U15528 ( n16184,n15991,n15528 );
   nand U15529 ( n16183,n15992,n15276 );
   or U15530 ( n16147,n16145,n16146 );
   and U15531 ( n16146,n16185,n16186 );
   nand U15532 ( n16186,n15991,n15273 );
   nand U15533 ( n16185,n15992,n15522 );
   nand U15534 ( n16145,n16187,n16188 );
   nand U15535 ( n16188,n15991,n15522 );
   nand U15536 ( n16187,n15992,n15273 );
   and U15537 ( n16144,n16189,n16190 );
   or U15538 ( n16190,n16191,n16192 );
   nand U15539 ( n16132,n16191,n16189,n16192 );
   and U15540 ( n16192,n16193,n16194 );
   nand U15541 ( n16194,n15991,n15270 );
   nand U15542 ( n16193,n15992,n15516 );
   nand U15543 ( n16189,n16138,n16139 );
   nand U15544 ( n16139,n16195,n16196 );
   nand U15545 ( n16196,n15991,n15267 );
   nand U15546 ( n16195,n15992,n15509 );
   and U15547 ( n16138,n16197,n16198 );
   nand U15548 ( n16198,n15991,n15509 );
   nand U15549 ( n16197,n15992,n15267 );
   nand U15550 ( n16191,n16199,n16200 );
   nand U15551 ( n16200,n15991,n15516 );
   nand U15552 ( n16199,n15992,n15270 );
   nand U15553 ( n16127,n16201,n16202 );
   or U15554 ( n16120,n16202,n16201 );
   and U15555 ( n16201,n16203,n16204 );
   nand U15556 ( n16204,n15991,n15489 );
   nand U15557 ( n16203,n15992,n15261 );
   nand U15558 ( n16202,n16205,n16206 );
   nand U15559 ( n16206,n15991,n15261 );
   nand U15560 ( n16205,n15992,n15489 );
   nand U15561 ( n16123,n16207,n16208 );
   nand U15562 ( n16208,n15991,n15480 );
   nand U15563 ( n16207,n15992,n15258 );
   nand U15564 ( n16124,n16209,n16210 );
   nand U15565 ( n16210,n15991,n15258 );
   nand U15566 ( n16209,n15992,n15480 );
   or U15567 ( n16113,n16119,n16118 );
   and U15568 ( n16118,n16211,n16212 );
   nand U15569 ( n16212,n15991,n15474 );
   nand U15570 ( n16211,n15992,n15255 );
   nand U15571 ( n16119,n16213,n16214 );
   nand U15572 ( n16214,n15991,n15255 );
   nand U15573 ( n16213,n15992,n15474 );
   nand U15574 ( n16094,n16215,n16216 );
   or U15575 ( n16092,n16216,n16215 );
   and U15576 ( n16215,n16217,n16218 );
   nand U15577 ( n16218,n15991,n15246 );
   nand U15578 ( n16217,n15992,n15444 );
   nand U15579 ( n16216,n16219,n16220 );
   nand U15580 ( n16220,n15991,n15444 );
   nand U15581 ( n16219,n15992,n15246 );
   or U15582 ( n16086,n16091,n16090 );
   and U15583 ( n16090,n16221,n16222 );
   nand U15584 ( n16222,n15991,n15243 );
   nand U15585 ( n16221,n15992,n15437 );
   nand U15586 ( n16091,n16223,n16224 );
   nand U15587 ( n16224,n15991,n15437 );
   nand U15588 ( n16223,n15992,n15243 );
   or U15589 ( n16067,n16078,n16077 );
   and U15590 ( n16077,n16225,n16226 );
   nand U15591 ( n16226,n15991,n15418 );
   nand U15592 ( n16225,n15992,n15237 );
   nand U15593 ( n16078,n16227,n16228 );
   nand U15594 ( n16228,n15991,n15237 );
   nand U15595 ( n16227,n15992,n15418 );
   nand U15596 ( n16070,n16229,n16230 );
   nand U15597 ( n16230,n15991,n15411 );
   nand U15598 ( n16229,n15992,n15234 );
   nand U15599 ( n16071,n16231,n16232 );
   nand U15600 ( n16232,n15991,n15234 );
   nand U15601 ( n16231,n15992,n15411 );
   nand U15602 ( n16058,n16233,n16234 );
   nand U15603 ( n16234,n15991,n15231 );
   nand U15604 ( n16233,n15992,n15401 );
   nand U15605 ( n16063,n16235,n16236 );
   nand U15606 ( n16236,n15991,n15401 );
   nand U15607 ( n16235,n15992,n15231 );
   nand U15608 ( n16052,n16040,n16041 );
   nand U15609 ( n16041,n16237,n16238 );
   nand U15610 ( n16238,n15991,n15372 );
   nand U15611 ( n16237,n15992,n15222 );
   and U15612 ( n16040,n16239,n16240 );
   nand U15613 ( n16240,n15991,n15222 );
   nand U15614 ( n16239,n15992,n15372 );
   nand U15615 ( n16051,n16046,n16047 );
   nand U15616 ( n16047,n16241,n16242 );
   nand U15617 ( n16242,n15991,n15661 );
   nand U15618 ( n16241,n15992,n15225 );
   and U15619 ( n16046,n16243,n16244 );
   nand U15620 ( n16244,n15991,n15225 );
   nand U15621 ( n16243,n15992,n15661 );
   or U15622 ( n16031,n16028,n16027 );
   and U15623 ( n16027,n16245,n16246 );
   nand U15624 ( n16246,n15991,n15219 );
   nand U15625 ( n16245,n15992,n15366 );
   nand U15626 ( n16028,n16247,n16248 );
   nand U15627 ( n16248,n15991,n15366 );
   nand U15628 ( n16247,n15992,n15219 );
   nand U15629 ( n16023,n16030,n16029 );
   nand U15630 ( n16029,n16249,n16250 );
   nand U15631 ( n16250,n15991,n15216 );
   nand U15632 ( n16249,n15992,n15357 );
   and U15633 ( n16030,n16251,n16252 );
   nand U15634 ( n16252,n15991,n15357 );
   nand U15635 ( n16251,n15992,n15216 );
   or U15636 ( n15949,n16018,n16017 );
   and U15637 ( n16017,n16253,n16254 );
   nand U15638 ( n16254,n15991,n15291 );
   nand U15639 ( n16253,n15992,n15192 );
   nand U15640 ( n16018,n16255,n16256 );
   nand U15641 ( n16256,n15991,n15192 );
   nand U15642 ( n16255,n15992,n15291 );
   nand U15643 ( n16259,n16260,n16257 );
   nand U15644 ( n15947,n16258,n16261 );
   nand U15645 ( n16261,n15577,n16262 );
   nand U15646 ( n15931,n16263,n15809,n16264 );
   xor U15647 ( n16263,n15577,n16265 );
   nand U15648 ( n16265,n16266,n16267,n16268,n16269 );
   nor U15649 ( n16269,n16270,n16271,n16272,n16273 );
   nand U15650 ( n16273,n16274,n15838,n16275,n16276 );
   and U15651 ( n15838,n16277,n16278 );
   or U15652 ( n16278,n15195,n16279 );
   or U15653 ( n16277,n15291,n15839 );
   nand U15654 ( n16272,n16280,n16281,n16282,n15835 );
   nand U15655 ( n15835,n16279,n15195 );
   not U15656 ( n16279,n15296 );
   nand U15657 ( n16282,n15839,n15291 );
   not U15658 ( n15839,n15192 );
   nand U15659 ( n16271,n16283,n16284,n16285,n16286 );
   nand U15660 ( n16270,n16287,n16288,n16289,n16290 );
   nor U15661 ( n16268,n16291,n16292,n16293,n16294 );
   or U15662 ( n16292,n16295,n16296,n16297 );
   nand U15663 ( n16291,n16298,n16299,n16300,n16301 );
   nor U15664 ( n16267,n16302,n16303,n16304,n16305 );
   and U15665 ( n16266,n16306,n16307,n16308,n16309 );
   nand U15666 ( p3_u3295,n16310,n16311,n16312 );
   nand U15667 ( n16312,n16313,si_0_ );
   nand U15668 ( n16311,p3_ir_reg_0_,n16314 );
   or U15669 ( n16314,n16315,n16316 );
   nand U15670 ( n16310,n16317,n16318 );
   nand U15671 ( p3_u3294,n16319,n16320,n16321,n16322 );
   nand U15672 ( n16322,p3_ir_reg_1_,n16323 );
   nand U15673 ( n16323,n16324,n16325 );
   nand U15674 ( n16325,n16316,n16326 );
   nand U15675 ( n16321,n16316,p3_ir_reg_0_,n16327 );
   nand U15676 ( n16320,n16317,n16328 );
   nand U15677 ( n16319,n16313,si_1_ );
   nand U15678 ( p3_u3293,n16329,n16330,n16331,n16332 );
   nand U15679 ( n16332,n16333,n16316 );
   not U15680 ( n16333,n16334 );
   nand U15681 ( n16331,n16317,n16335 );
   nand U15682 ( n16330,n16315,p3_ir_reg_2_ );
   nand U15683 ( n16329,n16313,si_2_ );
   nand U15684 ( p3_u3292,n16336,n16337,n16338,n16339 );
   nand U15685 ( n16339,p3_ir_reg_3_,n16340 );
   nand U15686 ( n16340,n16324,n16341 );
   nand U15687 ( n16341,n16316,n16342 );
   nand U15688 ( n16338,n16316,n16343,n16344 );
   nand U15689 ( n16337,n16317,n16345 );
   nand U15690 ( n16336,n16313,si_3_ );
   nand U15691 ( p3_u3291,n16346,n16347,n16348,n16349 );
   nand U15692 ( n16349,n16350,n16351,n16316 );
   nand U15693 ( n16348,n16317,n16352 );
   nand U15694 ( n16347,n16315,p3_ir_reg_4_ );
   nand U15695 ( n16346,n16313,si_4_ );
   nand U15696 ( p3_u3290,n16353,n16354,n16355,n16356 );
   nand U15697 ( n16356,p3_ir_reg_5_,n16357 );
   nand U15698 ( n16357,n16324,n16358 );
   nand U15699 ( n16358,n16316,n16359 );
   nand U15700 ( n16355,n16316,n16351,n16360 );
   nand U15701 ( n16354,n16317,n16361 );
   nand U15702 ( n16353,n16313,si_5_ );
   nand U15703 ( p3_u3289,n16362,n16363,n16364,n16365 );
   nand U15704 ( n16365,n16366,n16367,n16316 );
   nand U15705 ( n16364,n16317,n16368 );
   nand U15706 ( n16363,n16315,p3_ir_reg_6_ );
   nand U15707 ( n16362,n16313,si_6_ );
   nand U15708 ( p3_u3288,n16369,n16370,n16371,n16372 );
   nand U15709 ( n16372,p3_ir_reg_7_,n16373 );
   nand U15710 ( n16373,n16324,n16374 );
   nand U15711 ( n16374,n16316,n16375 );
   nand U15712 ( n16371,n16316,n16367,n16376 );
   nand U15713 ( n16370,n16317,n16377 );
   nand U15714 ( n16369,n16313,si_7_ );
   nand U15715 ( p3_u3287,n16378,n16379,n16380,n16381 );
   nand U15716 ( n16381,n16382,n16383,n16316 );
   nand U15717 ( n16380,n16315,p3_ir_reg_8_ );
   nand U15718 ( n16379,n16313,si_8_ );
   nand U15719 ( n16378,n16384,p3_u3151 );
   nand U15720 ( p3_u3286,n16385,n16386,n16387,n16388 );
   nand U15721 ( n16388,p3_ir_reg_9_,n16389 );
   nand U15722 ( n16389,n16324,n16390 );
   nand U15723 ( n16390,n16316,n16391 );
   nand U15724 ( n16387,n16316,n16383,n16392 );
   nand U15725 ( n16386,n16317,n16393 );
   nand U15726 ( n16385,n16313,si_9_ );
   nand U15727 ( p3_u3285,n16394,n16395,n16396,n16397 );
   nand U15728 ( n16397,n16398,n16316 );
   not U15729 ( n16398,n16399 );
   nand U15730 ( n16396,n16317,n16400 );
   nand U15731 ( n16395,n16315,p3_ir_reg_10_ );
   nand U15732 ( n16394,n16313,si_10_ );
   nand U15733 ( p3_u3284,n16401,n16402,n16403,n16404 );
   nand U15734 ( n16404,p3_ir_reg_11_,n16405 );
   nand U15735 ( n16405,n16324,n16406 );
   nand U15736 ( n16406,n16316,n16407 );
   nand U15737 ( n16403,n16316,n16408,n16409 );
   nand U15738 ( n16402,n16313,si_11_ );
   nand U15739 ( n16401,n16410,p3_u3151 );
   nand U15740 ( p3_u3283,n16411,n16412,n16413,n16414 );
   nand U15741 ( n16414,n16415,n16316 );
   not U15742 ( n16415,n16416 );
   nand U15743 ( n16413,n16315,p3_ir_reg_12_ );
   nand U15744 ( n16412,n16313,si_12_ );
   nand U15745 ( n16411,n16417,p3_u3151 );
   nand U15746 ( p3_u3282,n16418,n16419,n16420,n16421 );
   nand U15747 ( n16421,p3_ir_reg_13_,n16422 );
   nand U15748 ( n16422,n16324,n16423 );
   nand U15749 ( n16423,n16316,n16424 );
   nand U15750 ( n16420,n16316,n16425,n16426 );
   nand U15751 ( n16419,n16317,n16427 );
   nand U15752 ( n16418,n16313,si_13_ );
   nand U15753 ( p3_u3281,n16428,n16429,n16430,n16431 );
   nand U15754 ( n16431,n16432,n16316 );
   not U15755 ( n16432,n16433 );
   nand U15756 ( n16430,n16317,n16434 );
   nand U15757 ( n16429,n16315,p3_ir_reg_14_ );
   nand U15758 ( n16428,n16313,si_14_ );
   nand U15759 ( p3_u3280,n16435,n16436,n16437,n16438 );
   nand U15760 ( n16438,p3_ir_reg_15_,n16439 );
   nand U15761 ( n16439,n16324,n16440 );
   nand U15762 ( n16440,n16316,n16441 );
   nand U15763 ( n16437,n16316,n16442,n16443 );
   nand U15764 ( n16436,n16317,n16444 );
   nand U15765 ( n16435,n16313,si_15_ );
   nand U15766 ( p3_u3279,n16445,n16446,n16447,n16448 );
   nand U15767 ( n16448,n16449,n16316 );
   not U15768 ( n16449,n16450 );
   nand U15769 ( n16447,n16317,n16451 );
   nand U15770 ( n16446,n16315,p3_ir_reg_16_ );
   nand U15771 ( n16445,n16313,si_16_ );
   nand U15772 ( p3_u3278,n16452,n16453,n16454,n16455 );
   nand U15773 ( n16455,p3_ir_reg_17_,n16456 );
   nand U15774 ( n16456,n16324,n16457 );
   nand U15775 ( n16457,n16316,n16458 );
   nand U15776 ( n16454,n16316,n16459,n16460 );
   nand U15777 ( n16453,n16317,n16461 );
   nand U15778 ( n16452,n16313,si_17_ );
   nand U15779 ( p3_u3277,n16462,n16463,n16464,n16465 );
   nand U15780 ( n16465,p3_ir_reg_18_,n16466 );
   nand U15781 ( n16466,n16324,n16467 );
   nand U15782 ( n16467,n16316,n16468 );
   nand U15783 ( n16464,n16316,n16469,n16470 );
   nand U15784 ( n16463,n16317,n16471 );
   nand U15785 ( n16462,n16313,si_18_ );
   nand U15786 ( p3_u3276,n16472,n16473,n16474,n16475 );
   nand U15787 ( n16475,n16476,n16477,n16316 );
   nand U15788 ( n16474,n16317,n16478 );
   nand U15789 ( n16473,n16315,p3_ir_reg_19_ );
   nand U15790 ( n16472,n16313,si_19_ );
   nand U15791 ( p3_u3275,n16479,n16480,n16481,n16482 );
   nand U15792 ( n16482,n16483,n16484,n16316 );
   nand U15793 ( n16481,n16317,n16485 );
   nand U15794 ( n16480,n16315,p3_ir_reg_20_ );
   nand U15795 ( n16479,n16313,si_20_ );
   nand U15796 ( p3_u3274,n16486,n16487,n16488,n16489 );
   nand U15797 ( n16489,p3_ir_reg_21_,n16490 );
   nand U15798 ( n16490,n16324,n16491 );
   nand U15799 ( n16491,n16316,n16492 );
   nand U15800 ( n16488,n16316,n16484,n16493 );
   nand U15801 ( n16487,n16317,n16494 );
   nand U15802 ( n16486,n16313,si_21_ );
   nand U15803 ( p3_u3273,n16495,n16496,n16497,n16498 );
   nand U15804 ( n16498,n16499,n16316 );
   not U15805 ( n16499,n16500 );
   nand U15806 ( n16497,n16317,n16501 );
   nand U15807 ( n16496,n16315,p3_ir_reg_22_ );
   nand U15808 ( n16495,n16313,si_22_ );
   nand U15809 ( p3_u3272,n16502,n16503,n16504,n16505 );
   nand U15810 ( n16505,p3_ir_reg_23_,n16506 );
   nand U15811 ( n16506,n16324,n16507 );
   nand U15812 ( n16507,n16316,n16508 );
   nand U15813 ( n16504,n16316,n16509,n16510 );
   nand U15814 ( n16503,n16317,n16511 );
   nand U15815 ( n16502,n16313,si_23_ );
   nand U15816 ( p3_u3271,n16512,n16513,n16514,n16515 );
   nand U15817 ( n16515,n16516,n16316 );
   not U15818 ( n16516,n16517 );
   nand U15819 ( n16514,n16317,n16518 );
   nand U15820 ( n16513,n16315,p3_ir_reg_24_ );
   nand U15821 ( n16512,n16313,si_24_ );
   nand U15822 ( p3_u3270,n16519,n16520,n16521,n16522 );
   nand U15823 ( n16522,p3_ir_reg_25_,n16523 );
   nand U15824 ( n16523,n16324,n16524 );
   nand U15825 ( n16524,n16316,n16525 );
   nand U15826 ( n16521,n16316,n16526,n16527 );
   nand U15827 ( n16520,n16317,n16528 );
   nand U15828 ( n16519,n16313,si_25_ );
   nand U15829 ( p3_u3269,n16529,n16530,n16531,n16532 );
   nand U15830 ( n16532,n16533,n16316 );
   not U15831 ( n16533,n16534 );
   nand U15832 ( n16531,n16317,n16535 );
   nand U15833 ( n16530,n16315,p3_ir_reg_26_ );
   nand U15834 ( n16529,n16313,si_26_ );
   nand U15835 ( p3_u3268,n16536,n16537,n16538,n16539 );
   nand U15836 ( n16539,p3_ir_reg_27_,n16540 );
   nand U15837 ( n16540,n16324,n16541 );
   nand U15838 ( n16541,n16316,n16542 );
   nand U15839 ( n16538,n16316,n16543,n16544 );
   nand U15840 ( n16537,n16317,n16545 );
   nand U15841 ( n16536,n16313,si_27_ );
   nand U15842 ( p3_u3267,n16546,n16547,n16548,n16549 );
   nand U15843 ( n16549,p3_ir_reg_28_,n16550 );
   nand U15844 ( n16550,n16324,n16551 );
   nand U15845 ( n16551,n16316,n16552 );
   nand U15846 ( n16548,n16316,n16553,n16554 );
   nand U15847 ( n16547,n16317,n16555 );
   nand U15848 ( n16546,n16313,si_28_ );
   nand U15849 ( p3_u3266,n16556,n16557,n16558,n16559 );
   nand U15850 ( n16559,n16560,n16561,n16316 );
   nand U15851 ( n16558,n16317,n16562 );
   nand U15852 ( n16557,n16315,p3_ir_reg_29_ );
   nand U15853 ( n16556,n16313,si_29_ );
   nand U15854 ( p3_u3265,n16563,n16564,n16565,n16566 );
   nand U15855 ( n16566,p3_ir_reg_30_,n16567 );
   nand U15856 ( n16567,n16324,n16568 );
   nand U15857 ( n16568,n16569,n16316 );
   nand U15858 ( n16565,n16316,n16561,n16570 );
   not U15859 ( n16561,n16569 );
   nand U15860 ( n16564,n16317,n16571 );
   nand U15861 ( n16563,n16313,si_30_ );
   nand U15862 ( p3_u3264,n16573,n16574,n16575 );
   nand U15863 ( n16575,n16313,si_31_ );
   nand U15864 ( n16574,n16316,n16570,n16569 );
   nor U15865 ( n16569,n16577,p3_ir_reg_29_ );
   not U15866 ( n16315,n16324 );
   nand U15867 ( n16324,p3_state_reg,n16578 );
   nand U15868 ( n16573,n16579,p3_u3151 );
   nor U15869 ( p3_u3263,n15814,n16580 );
   and U15870 ( p3_u3262,n15813,p3_d_reg_3_ );
   and U15871 ( p3_u3261,n15813,p3_d_reg_4_ );
   and U15872 ( p3_u3260,n15813,p3_d_reg_5_ );
   nor U15873 ( p3_u3259,n15814,n16581 );
   and U15874 ( p3_u3258,n15813,p3_d_reg_7_ );
   and U15875 ( p3_u3257,n15813,p3_d_reg_8_ );
   and U15876 ( p3_u3256,n15813,p3_d_reg_9_ );
   nor U15877 ( p3_u3255,n15814,n16582 );
   and U15878 ( p3_u3254,n15813,p3_d_reg_11_ );
   and U15879 ( p3_u3253,n15813,p3_d_reg_12_ );
   nor U15880 ( p3_u3252,n15814,n16583 );
   and U15881 ( p3_u3251,n15813,p3_d_reg_14_ );
   and U15882 ( p3_u3250,n15813,p3_d_reg_15_ );
   nor U15883 ( p3_u3249,n15814,n16584 );
   nor U15884 ( p3_u3248,n15814,n16585 );
   nor U15885 ( p3_u3247,n15814,n16586 );
   nor U15886 ( p3_u3246,n15814,n16587 );
   and U15887 ( p3_u3245,n15813,p3_d_reg_20_ );
   and U15888 ( p3_u3244,n15813,p3_d_reg_21_ );
   and U15889 ( p3_u3243,n15813,p3_d_reg_22_ );
   and U15890 ( p3_u3242,n15813,p3_d_reg_23_ );
   and U15891 ( p3_u3241,n15813,p3_d_reg_24_ );
   and U15892 ( p3_u3240,n15813,p3_d_reg_25_ );
   and U15893 ( p3_u3239,n15813,p3_d_reg_26_ );
   nor U15894 ( p3_u3238,n15814,n16588 );
   and U15895 ( p3_u3237,n15813,p3_d_reg_28_ );
   nor U15896 ( p3_u3236,n15814,n16589 );
   and U15897 ( p3_u3235,n15813,p3_d_reg_30_ );
   and U15898 ( p3_u3234,n15813,p3_d_reg_31_ );
   nand U15899 ( p3_u3233,n16591,n16592,n16593,n16594 );
   nor U15900 ( n16594,n16595,n16596,n16597 );
   nor U15901 ( n16597,n15796,n16598 );
   nor U15902 ( n16596,n15797,n16599 );
   not U15903 ( n15797,n15557 );
   nor U15904 ( n16595,n16600,n16601 );
   nand U15905 ( n16593,n16602,n15561 );
   nand U15906 ( n16592,p3_reg2_reg_0_,n16603 );
   nand U15907 ( n16591,n16604,n15565 );
   nand U15908 ( n15565,n16605,n16606 );
   nand U15909 ( n16606,n15557,n16607 );
   nand U15910 ( n16605,n16293,n16608 );
   and U15911 ( n16293,n16609,n16610 );
   nand U15912 ( n16609,n16170,n16611 );
   nand U15913 ( p3_u3232,n16612,n16613,n16614,n16615 );
   nor U15914 ( n16615,n16616,n16617,n16618 );
   nor U15915 ( n16618,n15552,n16603 );
   and U15916 ( n15552,n16619,n16620,n16621,n16622 );
   nor U15917 ( n16622,n16623,n16624,n16625,n16626 );
   nor U15918 ( n16626,n16627,n16628 );
   nor U15919 ( n16625,n16627,n15828 );
   nor U15920 ( n16624,n16629,n16630 );
   nor U15921 ( n16623,n16627,n16631 );
   nor U15922 ( n16621,n16632,n16633 );
   nor U15923 ( n16633,n16629,n16634 );
   not U15924 ( n16629,n15547 );
   nor U15925 ( n16632,n16627,n15831 );
   xor U15926 ( n16627,n16635,n16283 );
   nand U15927 ( n16620,n16636,n15285 );
   nand U15928 ( n16619,n16637,n15547 );
   nor U15929 ( n16617,n16604,n16638 );
   nor U15930 ( n16616,n16639,n16640 );
   nand U15931 ( n16614,n16641,p3_reg3_reg_1_ );
   nand U15932 ( n16613,n16642,n15547 );
   xor U15933 ( n15547,n16643,n16283 );
   nand U15934 ( n16283,n16644,n16645 );
   nand U15935 ( n16612,n16646,n15279 );
   nand U15936 ( p3_u3231,n16647,n16648,n16649,n16650 );
   nor U15937 ( n16650,n16651,n16652,n16653 );
   nor U15938 ( n16653,n15783,n16598 );
   nor U15939 ( n16652,n15537,n16599 );
   and U15940 ( n16651,p3_reg3_reg_2_,n16641 );
   nand U15941 ( n16649,n16602,n15538 );
   nand U15942 ( n16648,p3_reg2_reg_2_,n16603 );
   nand U15943 ( n16647,n16604,n15541 );
   nand U15944 ( n15541,n16654,n16655,n16656,n16657 );
   nand U15945 ( n16657,n16658,n16659,n16660 );
   nand U15946 ( n16658,n16661,n16662,n16663 );
   or U15947 ( n16656,n15537,n16664 );
   nand U15948 ( n15537,n16665,n16659 );
   nand U15949 ( n16659,n16666,n16667 );
   nand U15950 ( n16665,n16668,n16662 );
   not U15951 ( n16668,n16669 );
   nand U15952 ( n16655,n16670,n16671,n16608 );
   nand U15953 ( n16671,n16666,n16672 );
   not U15954 ( n16666,n16274 );
   xor U15955 ( n16274,n16673,n15279 );
   nand U15956 ( n16670,n16661,n16662,n16674 );
   not U15957 ( n16674,n16672 );
   nand U15958 ( n16672,n16675,n16644 );
   nand U15959 ( n16654,n16636,n15282 );
   nand U15960 ( p3_u3230,n16676,n16677,n16678,n16679 );
   nor U15961 ( n16679,n16680,n16681,n16682 );
   nor U15962 ( n16682,n15532,n16603 );
   and U15963 ( n15532,n16683,n16684,n16685,n16686 );
   nor U15964 ( n16686,n16687,n16688,n16689,n16690 );
   nor U15965 ( n16690,n16691,n16692 );
   nor U15966 ( n16689,n15828,n16693 );
   nor U15967 ( n16688,n16631,n16693 );
   and U15968 ( n16687,n15527,n16637 );
   nor U15969 ( n16685,n16694,n16695 );
   nor U15970 ( n16695,n16696,n16634 );
   nor U15971 ( n16696,n16697,n16698 );
   not U15972 ( n16698,n16699 );
   nor U15973 ( n16697,n16700,n16275 );
   nor U15974 ( n16694,n16628,n16693 );
   or U15975 ( n16684,n16693,n15831 );
   xor U15976 ( n16693,n16701,n16702 );
   nor U15977 ( n16701,n16703,n16704 );
   nand U15978 ( n16683,n16705,n15527 );
   nor U15979 ( n16681,n16604,n16706 );
   nor U15980 ( n16680,n16707,n16640 );
   nand U15981 ( n16678,n16641,n16708 );
   nand U15982 ( n16677,n16642,n15527 );
   nand U15983 ( n15527,n16709,n16699 );
   nand U15984 ( n16699,n16275,n16700 );
   nand U15985 ( n16709,n16710,n16661,n16702 );
   not U15986 ( n16702,n16275 );
   xor U15987 ( n16275,n16707,n15276 );
   nand U15988 ( n16710,n16667,n16662 );
   nand U15989 ( n16676,n16646,n15273 );
   nand U15990 ( p3_u3229,n16711,n16712,n16713,n16714 );
   nor U15991 ( n16714,n16715,n16716,n16717 );
   nor U15992 ( n16717,n16718,n16598 );
   and U15993 ( n16716,n15769,n16642 );
   and U15994 ( n16715,n16719,n16641 );
   nand U15995 ( n16713,n16602,n15522 );
   nand U15996 ( n16712,p3_reg2_reg_4_,n16603 );
   nand U15997 ( n16711,n16604,n15770 );
   nand U15998 ( n15770,n16720,n16721,n16722 );
   nand U15999 ( n16722,n16636,n15276 );
   nand U16000 ( n16721,n16723,n16608 );
   xor U16001 ( n16723,n16724,n16284 );
   nand U16002 ( n16720,n15769,n16607 );
   nand U16003 ( n15769,n16725,n16726 );
   nand U16004 ( n16726,n16284,n16727 );
   nand U16005 ( n16284,n16728,n16729 );
   nand U16006 ( n16725,n16730,n16731 );
   nand U16007 ( n16731,n16732,n16733 );
   nand U16008 ( p3_u3228,n16734,n16735,n16736,n16737 );
   nor U16009 ( n16737,n16738,n16739,n16740 );
   nor U16010 ( n16740,n16741,n16598 );
   and U16011 ( n16739,n15761,n16642 );
   and U16012 ( n16738,n16742,n16641 );
   nand U16013 ( n16736,n16602,n15516 );
   nand U16014 ( n16735,p3_reg2_reg_5_,n16603 );
   nand U16015 ( n16734,n16604,n15762 );
   nand U16016 ( n15762,n16743,n16744,n16745 );
   nand U16017 ( n16745,n16636,n15273 );
   nand U16018 ( n16744,n16746,n16747,n16608 );
   nand U16019 ( n16747,n16748,n16285 );
   nand U16020 ( n16748,n16749,n16729 );
   nand U16021 ( n16746,n16749,n16729,n16750 );
   not U16022 ( n16750,n16285 );
   nand U16023 ( n16749,n16724,n16728 );
   not U16024 ( n16724,n16751 );
   nand U16025 ( n16743,n15761,n16607 );
   nand U16026 ( n15761,n16752,n16753 );
   nand U16027 ( n16753,n15916,n16285 );
   nand U16028 ( n16285,n16754,n16755 );
   not U16029 ( n15916,n16756 );
   nand U16030 ( n16752,n16757,n16756 );
   nand U16031 ( n16757,n16758,n16759 );
   nand U16032 ( p3_u3227,n16760,n16761,n16762,n16763 );
   nor U16033 ( n16763,n16764,n16765,n16766 );
   nor U16034 ( n16766,n15507,n16598 );
   nor U16035 ( n16765,n15508,n16599 );
   and U16036 ( n15508,n16767,n16768 );
   and U16037 ( n16764,n16769,n16641 );
   nand U16038 ( n16762,n16602,n15509 );
   nand U16039 ( n16761,p3_reg2_reg_6_,n16603 );
   nand U16040 ( n16760,n16604,n15510 );
   nand U16041 ( n15510,n16770,n16771,n16772,n16773 );
   nor U16042 ( n16773,n16774,n16775,n16776,n16777 );
   and U16043 ( n16777,n16778,n16705 );
   nor U16044 ( n16776,n16779,n15828 );
   nor U16045 ( n16775,n16718,n16692 );
   nor U16046 ( n16774,n16779,n15831 );
   nand U16047 ( n16772,n16637,n16778 );
   or U16048 ( n16771,n16779,n16780 );
   xor U16049 ( n16779,n16781,n16782 );
   nand U16050 ( n16770,n16660,n16778 );
   nand U16051 ( n16778,n16767,n16768 );
   nand U16052 ( n16768,n16783,n16781 );
   not U16053 ( n16783,n16758 );
   and U16054 ( n16767,n16784,n16785 );
   nand U16055 ( n16785,n16756,n16759,n16781 );
   not U16056 ( n16781,n16286 );
   nand U16057 ( n16286,n16786,n16787 );
   nand U16058 ( n16784,n16788,n15912,n15917 );
   nand U16059 ( n16788,n16756,n16759 );
   nand U16060 ( n16756,n16733,n16789 );
   nand U16061 ( n16789,n16730,n16732 );
   nand U16062 ( p3_u3226,n16790,n16791,n16792,n16793 );
   nor U16063 ( n16793,n16794,n16795,n16796 );
   nor U16064 ( n16796,n15908,n16598 );
   nor U16065 ( n16795,n16797,n16599 );
   and U16066 ( n16794,n16798,n16641 );
   nand U16067 ( n16792,n16602,n15496 );
   nand U16068 ( n16791,p3_reg2_reg_7_,n16603 );
   nand U16069 ( n16790,n16604,n15748 );
   nand U16070 ( n15748,n16799,n16800,n16801,n16802 );
   nor U16071 ( n16802,n16803,n16804,n16805,n16806 );
   nor U16072 ( n16806,n16631,n16807 );
   nor U16073 ( n16805,n15828,n16807 );
   nor U16074 ( n16804,n16634,n16797 );
   nor U16075 ( n16803,n16630,n16797 );
   nor U16076 ( n16801,n16808,n16809 );
   nor U16077 ( n16809,n16741,n16692 );
   nor U16078 ( n16808,n15831,n16807 );
   nand U16079 ( n16800,n15495,n16637 );
   not U16080 ( n15495,n16797 );
   nand U16081 ( n16797,n16810,n16811 );
   nand U16082 ( n16811,n16812,n15910 );
   not U16083 ( n16812,n16813 );
   nand U16084 ( n16810,n16814,n16815 );
   or U16085 ( n16799,n16807,n16628 );
   nand U16086 ( n16807,n16816,n16817 );
   nand U16087 ( n16817,n16818,n16287 );
   nand U16088 ( n16818,n16819,n16787 );
   nand U16089 ( n16816,n16819,n16787,n16814 );
   not U16090 ( n16814,n16287 );
   nand U16091 ( n16287,n16820,n16821 );
   nand U16092 ( n16819,n16786,n16782 );
   nand U16093 ( p3_u3225,n16822,n16823,n16824,n16825 );
   nor U16094 ( n16825,n16826,n16827,n16828 );
   nor U16095 ( n16828,n15487,n16598 );
   nor U16096 ( n16827,n15488,n16599 );
   not U16097 ( n15488,n16829 );
   nor U16098 ( n16826,n16830,n16601 );
   nand U16099 ( n16824,n16602,n15489 );
   nand U16100 ( n16823,p3_reg2_reg_8_,n16603 );
   nand U16101 ( n16822,n16604,n15490 );
   nand U16102 ( n15490,n16831,n16832,n16833,n16834 );
   nand U16103 ( n16834,n16835,n16288 );
   nand U16104 ( n16835,n16836,n16837 );
   nand U16105 ( n16837,n16838,n16839 );
   nand U16106 ( n16836,n16840,n16608 );
   nand U16107 ( n16833,n16841,n16842 );
   nand U16108 ( n16842,n16843,n16844 );
   nand U16109 ( n16844,n16839,n16845 );
   nand U16110 ( n16843,n16608,n16846 );
   nand U16111 ( n16832,n16637,n16829 );
   nand U16112 ( n16829,n16847,n16848 );
   nand U16113 ( n16848,n16838,n16288 );
   not U16114 ( n16288,n16841 );
   nand U16115 ( n16847,n16849,n15906,n16841 );
   nor U16116 ( n16841,n16850,n16851 );
   nor U16117 ( n16851,n15261,n15489 );
   nand U16118 ( n16849,n16815,n15910 );
   not U16119 ( n16815,n16852 );
   nand U16120 ( n16831,n16636,n15264 );
   nand U16121 ( p3_u3224,n16853,n16854,n16855,n16856 );
   nor U16122 ( n16856,n16857,n16858,n16859 );
   nor U16123 ( n16859,n16860,n16598 );
   and U16124 ( n16858,n15734,n16642 );
   and U16125 ( n16857,n16861,n16641 );
   nand U16126 ( n16855,n16602,n15480 );
   nand U16127 ( n16854,p3_reg2_reg_9_,n16603 );
   nand U16128 ( n16853,n16604,n15735 );
   nand U16129 ( n15735,n16862,n16863,n16864 );
   nand U16130 ( n16864,n16636,n15261 );
   nand U16131 ( n16863,n16865,n16866 );
   nand U16132 ( n16866,n15831,n15828,n16780 );
   xor U16133 ( n16865,n16289,n16867 );
   nand U16134 ( n16862,n15734,n16607 );
   nand U16135 ( n15734,n16868,n16869 );
   nand U16136 ( n16869,n16870,n16871 );
   nand U16137 ( n16870,n16872,n15900 );
   nand U16138 ( n16868,n16873,n16289 );
   nand U16139 ( n16289,n16874,n16875 );
   not U16140 ( n16873,n16871 );
   nand U16141 ( p3_u3223,n16876,n16877,n16878,n16879 );
   nor U16142 ( n16879,n16880,n16881,n16882 );
   nor U16143 ( n16882,n16883,n16598 );
   and U16144 ( n16881,n15726,n16642 );
   and U16145 ( n16880,n16884,n16641 );
   nand U16146 ( n16878,n16602,n15474 );
   nand U16147 ( n16877,p3_reg2_reg_10_,n16603 );
   nand U16148 ( n16876,n16604,n15727 );
   nand U16149 ( n15727,n16885,n16886,n16887 );
   nand U16150 ( n16887,n16636,n15258 );
   nand U16151 ( n16886,n16888,n16889,n16608 );
   not U16152 ( n16608,n16890 );
   nand U16153 ( n16889,n16891,n16874,n16290 );
   nand U16154 ( n16891,n16892,n16875 );
   not U16155 ( n16892,n16867 );
   nand U16156 ( n16888,n16893,n16875,n16894 );
   not U16157 ( n16894,n16290 );
   nand U16158 ( n16893,n16867,n16874 );
   nor U16159 ( n16867,n16895,n16850 );
   nand U16160 ( n16885,n15726,n16896 );
   nand U16161 ( n16896,n16664,n16634 );
   nor U16162 ( n16664,n16705,n16637 );
   nand U16163 ( n15726,n16897,n16898 );
   nand U16164 ( n16898,n16899,n16290 );
   nand U16165 ( n16290,n16900,n16901 );
   nand U16166 ( n16897,n16902,n16903 );
   nand U16167 ( n16902,n15899,n16904 );
   nand U16168 ( p3_u3222,n16905,n16906,n16907,n16908 );
   nor U16169 ( n16908,n16909,n16910,n16911 );
   nor U16170 ( n16911,n15468,n16603 );
   and U16171 ( n15468,n16912,n16913,n16914,n16915 );
   nor U16172 ( n16915,n16916,n16917,n16918,n16919 );
   nor U16173 ( n16919,n16628,n16920 );
   nor U16174 ( n16918,n16631,n16920 );
   xor U16175 ( n16920,n16921,n16297 );
   nor U16176 ( n16917,n16922,n16923 );
   nor U16177 ( n16916,n15831,n16924 );
   xor U16178 ( n16924,n16297,n16925 );
   nor U16179 ( n16914,n16926,n16927 );
   nor U16180 ( n16927,n16860,n16692 );
   nor U16181 ( n16926,n16922,n16634 );
   not U16182 ( n16922,n15463 );
   nand U16183 ( n16913,n16928,n16929 );
   xor U16184 ( n16928,n16297,n16930 );
   nand U16185 ( n16912,n16705,n15463 );
   nor U16186 ( n16910,n16604,n16931 );
   nor U16187 ( n16909,n16932,n16640 );
   nand U16188 ( n16907,n16641,n16933 );
   nand U16189 ( n16906,n16642,n15463 );
   nand U16190 ( n15463,n16934,n16935 );
   nand U16191 ( n16935,n16936,n15923,n16937 );
   nand U16192 ( n16936,n15899,n16903 );
   not U16193 ( n16903,n16899 );
   nand U16194 ( n16934,n16938,n15899,n16297 );
   nor U16195 ( n16297,n16939,n16940 );
   nand U16196 ( n16938,n16899,n16904 );
   nor U16197 ( n16899,n16941,n16942 );
   nand U16198 ( n16905,n16646,n15249 );
   nand U16199 ( p3_u3221,n16943,n16944,n16945,n16946 );
   nor U16200 ( n16946,n16947,n16948,n16949 );
   nor U16201 ( n16949,n15458,n16603 );
   and U16202 ( n15458,n16950,n16951,n16952,n16953 );
   nor U16203 ( n16953,n16954,n16955,n16956,n16957 );
   nor U16204 ( n16957,n16628,n16958 );
   nor U16205 ( n16956,n15828,n16959 );
   nor U16206 ( n16955,n16960,n16630 );
   nor U16207 ( n16954,n16631,n16958 );
   xor U16208 ( n16958,n16309,n16961 );
   nor U16209 ( n16952,n16962,n16963 );
   nor U16210 ( n16963,n16960,n16634 );
   nor U16211 ( n16962,n15831,n16959 );
   xor U16212 ( n16959,n16309,n16964 );
   nand U16213 ( n16951,n16636,n15252 );
   nand U16214 ( n16950,n16637,n15453 );
   nor U16215 ( n16948,n16604,n16965 );
   nor U16216 ( n16947,n16966,n16640 );
   nand U16217 ( n16945,n16641,n16967 );
   nand U16218 ( n16944,n16642,n15453 );
   not U16219 ( n15453,n16960 );
   xor U16220 ( n16960,n16309,n16968 );
   nand U16221 ( n16309,n16969,n16970 );
   nand U16222 ( n16943,n16646,n15246 );
   nand U16223 ( p3_u3220,n16971,n16972,n16973,n16974 );
   nor U16224 ( n16974,n16975,n16976,n16977 );
   nor U16225 ( n16977,n15448,n16603 );
   and U16226 ( n15448,n16978,n16979 );
   nor U16227 ( n16979,n16980,n16981,n16982,n16983 );
   nor U16228 ( n16983,n16630,n16984 );
   nor U16229 ( n16982,n16985,n16692 );
   nor U16230 ( n16981,n16923,n16984 );
   nor U16231 ( n16980,n16628,n16986,n16987 );
   nor U16232 ( n16978,n16988,n16989,n16990,n16991 );
   nor U16233 ( n16991,n16634,n16984 );
   nor U16234 ( n16990,n16631,n16986,n16987 );
   and U16235 ( n16987,n16992,n16993 );
   nand U16236 ( n16993,n16994,n16970 );
   and U16237 ( n16986,n16308,n16970,n16995 );
   nand U16238 ( n16995,n16969,n16961 );
   not U16239 ( n16961,n16994 );
   nor U16240 ( n16994,n16996,n16940 );
   nor U16241 ( n16989,n15828,n16997 );
   nor U16242 ( n16988,n15831,n16997 );
   nand U16243 ( n16997,n16998,n16999 );
   nand U16244 ( n16999,n16992,n17000 );
   nand U16245 ( n17000,n17001,n16970 );
   and U16246 ( n16992,n17002,n17003 );
   nand U16247 ( n16998,n16308,n16970,n17004 );
   nand U16248 ( n17004,n16964,n16969 );
   not U16249 ( n16964,n17001 );
   nor U16250 ( n17001,n17005,n16940 );
   nor U16251 ( n16976,n16604,n17006 );
   nor U16252 ( n16975,n17007,n16640 );
   nand U16253 ( n16973,n16641,n17008 );
   nand U16254 ( n16972,n16642,n15443 );
   not U16255 ( n15443,n16984 );
   xor U16256 ( n16984,n17009,n16308 );
   nand U16257 ( n16308,n17003,n17010 );
   nand U16258 ( n16971,n16646,n15243 );
   nand U16259 ( p3_u3219,n17011,n17012,n17013,n17014 );
   nor U16260 ( n17014,n17015,n17016,n17017 );
   nor U16261 ( n17017,n15435,n16598 );
   nor U16262 ( n17016,n15436,n16599 );
   not U16263 ( n15436,n17018 );
   nor U16264 ( n17015,n17019,n16601 );
   nand U16265 ( n17013,n16602,n15437 );
   nand U16266 ( n17012,p3_reg2_reg_14_,n16603 );
   nand U16267 ( n17011,n16604,n15438 );
   nand U16268 ( n15438,n17020,n17021,n17022,n17023 );
   nand U16269 ( n17023,n17024,n16307 );
   nand U16270 ( n17024,n17025,n17026 );
   nand U16271 ( n17026,n17027,n17028 );
   nand U16272 ( n17025,n17029,n17030 );
   nand U16273 ( n17022,n17031,n17032 );
   nand U16274 ( n17032,n17033,n17034 );
   nand U16275 ( n17034,n17035,n17027 );
   nand U16276 ( n17033,n17036,n17029 );
   not U16277 ( n17031,n16307 );
   nand U16278 ( n17021,n17018,n16607 );
   nand U16279 ( n17018,n17037,n17038 );
   nand U16280 ( n17038,n16307,n17039 );
   nand U16281 ( n16307,n17040,n17041 );
   nand U16282 ( n17037,n17042,n17043 );
   nand U16283 ( n17043,n15894,n15890 );
   not U16284 ( n17042,n17039 );
   nand U16285 ( n17020,n16636,n15246 );
   nand U16286 ( p3_u3218,n17044,n17045,n17046,n17047 );
   nor U16287 ( n17047,n17048,n17049,n17050 );
   nor U16288 ( n17050,n17051,n16598 );
   and U16289 ( n17049,n15694,n16642 );
   and U16290 ( n17048,n17052,n16641 );
   nand U16291 ( n17046,n16602,n15428 );
   nand U16292 ( n17045,p3_reg2_reg_15_,n16603 );
   nand U16293 ( n17044,n16604,n15695 );
   nand U16294 ( n15695,n17053,n17054,n17055,n17056 );
   nand U16295 ( n17056,n17057,n17029 );
   xor U16296 ( n17057,n16306,n17058 );
   nand U16297 ( n17055,n17059,n17027 );
   xor U16298 ( n17059,n16306,n17060 );
   nand U16299 ( n17054,n15694,n16607 );
   nand U16300 ( n15694,n17061,n17062 );
   nand U16301 ( n17062,n17063,n16306 );
   nand U16302 ( n16306,n17064,n17065 );
   nand U16303 ( n17061,n17066,n17067 );
   nand U16304 ( n17066,n15887,n15886 );
   nand U16305 ( n17053,n16636,n15243 );
   nand U16306 ( p3_u3217,n17068,n17069,n17070,n17071 );
   nor U16307 ( n17071,n17072,n17073,n17074 );
   nor U16308 ( n17074,n15422,n16603 );
   and U16309 ( n15422,n17075,n17076 );
   nor U16310 ( n17076,n17077,n17078,n17079,n17080 );
   nor U16311 ( n17080,n17081,n16630 );
   nor U16312 ( n17079,n17082,n15828 );
   nor U16313 ( n17078,n15435,n16692 );
   nor U16314 ( n17077,n17081,n16634 );
   nor U16315 ( n17075,n17083,n17084,n17085,n17086 );
   nor U16316 ( n17086,n17087,n16628 );
   nor U16317 ( n17085,n17081,n16923 );
   not U16318 ( n17081,n15417 );
   nor U16319 ( n17084,n17087,n16631 );
   xor U16320 ( n17087,n16305,n17088 );
   nor U16321 ( n17083,n17082,n15831 );
   xor U16322 ( n17082,n16305,n17089 );
   nor U16323 ( n17073,n16604,n17090 );
   nor U16324 ( n17072,n17091,n16640 );
   nand U16325 ( n17070,n16641,n17092 );
   nand U16326 ( n17069,n16642,n15417 );
   nand U16327 ( n15417,n17093,n17094 );
   nand U16328 ( n17094,n17095,n15883,n17096 );
   nand U16329 ( n17095,n15887,n17067 );
   not U16330 ( n17067,n17063 );
   nand U16331 ( n17093,n17097,n15887,n16305 );
   and U16332 ( n16305,n17098,n17099 );
   nand U16333 ( n17097,n17063,n15886 );
   nor U16334 ( n17063,n17100,n17101 );
   nand U16335 ( n17068,n16646,n15234 );
   nand U16336 ( p3_u3216,n17102,n17103,n17104,n17105 );
   nor U16337 ( n17105,n17106,n17107,n17108 );
   nor U16338 ( n17108,n15409,n16598 );
   nor U16339 ( n17107,n15410,n16599 );
   not U16340 ( n15410,n17109 );
   nor U16341 ( n17106,n17110,n16601 );
   not U16342 ( n16601,n16641 );
   nand U16343 ( n17104,n16602,n15411 );
   nand U16344 ( n17103,p3_reg2_reg_17_,n16603 );
   nand U16345 ( n17102,n16604,n15412 );
   nand U16346 ( n15412,n17111,n17112,n17113,n17114 );
   nand U16347 ( n17114,n17029,n17115,n17116 );
   nand U16348 ( n17116,n17117,n17118 );
   nand U16349 ( n17118,n17088,n17099 );
   nand U16350 ( n17115,n17119,n17099,n16276 );
   nand U16351 ( n17119,n17120,n17098 );
   nand U16352 ( n17113,n17121,n17027,n17122 );
   nand U16353 ( n17122,n17117,n17123 );
   nand U16354 ( n17123,n17089,n17099 );
   and U16355 ( n17117,n17124,n17125 );
   nand U16356 ( n17125,n15411,n15234 );
   nand U16357 ( n17121,n17126,n17099,n16276 );
   nand U16358 ( n17126,n17127,n17098 );
   nand U16359 ( n17112,n17109,n16607 );
   xor U16360 ( n17109,n16276,n17128 );
   xor U16361 ( n16276,n15411,n17129 );
   nand U16362 ( n17111,n16636,n15237 );
   nand U16363 ( p3_u3215,n17130,n17131,n17132,n17133 );
   nor U16364 ( n17133,n17134,n17135,n17136 );
   nor U16365 ( n17136,n15397,n16598 );
   nor U16366 ( n17135,n15400,n16599 );
   and U16367 ( n17134,n17137,n16641 );
   nand U16368 ( n17132,n16602,n15401 );
   nand U16369 ( n17131,p3_reg2_reg_18_,n16603 );
   nand U16370 ( n17130,n16604,n15402 );
   nand U16371 ( n15402,n17138,n17139,n17140,n17141 );
   nor U16372 ( n17141,n17142,n17143,n17144,n17145 );
   nor U16373 ( n17145,n17129,n16692 );
   nor U16374 ( n17144,n15831,n17146 );
   xor U16375 ( n17146,n17147,n17148 );
   nor U16376 ( n17143,n16630,n15400 );
   not U16377 ( n15400,n17149 );
   nor U16378 ( n17142,n16628,n17150 );
   xor U16379 ( n17150,n17151,n17148 );
   nand U16380 ( n17140,n17152,n16929 );
   not U16381 ( n16929,n15828 );
   xor U16382 ( n17152,n17147,n16304 );
   nand U16383 ( n17139,n17149,n17153 );
   nand U16384 ( n17153,n16634,n16923 );
   xor U16385 ( n17149,n16304,n17154 );
   nand U16386 ( n17138,n17155,n17156 );
   xor U16387 ( n17155,n17151,n16304 );
   not U16388 ( n16304,n17148 );
   nand U16389 ( n17148,n17157,n17158 );
   nand U16390 ( p3_u3214,n17159,n17160,n17161,n17162 );
   nor U16391 ( n17162,n17163,n17164,n17165 );
   nor U16392 ( n17165,n15390,n16603 );
   and U16393 ( n15390,n17166,n17167,n17168,n17169 );
   nor U16394 ( n17169,n17170,n17171,n17172,n17173 );
   nor U16395 ( n17173,n16628,n17174 );
   xor U16396 ( n17174,n17175,n16295 );
   nor U16397 ( n17172,n15828,n17176 );
   nor U16398 ( n17171,n15409,n16692 );
   nor U16399 ( n17170,n16923,n17177 );
   nor U16400 ( n17168,n17178,n17179 );
   nor U16401 ( n17179,n15831,n17176 );
   xor U16402 ( n17176,n17180,n16295 );
   nor U16403 ( n17178,n16630,n17177 );
   not U16404 ( n17177,n15386 );
   nand U16405 ( n17167,n17181,n17156 );
   xor U16406 ( n17181,n17175,n17182 );
   nand U16407 ( n17166,n15386,n16660 );
   and U16408 ( n17164,n16603,p3_reg2_reg_19_ );
   nor U16409 ( n17163,n15874,n16640 );
   nand U16410 ( n17161,n16641,n17183 );
   nand U16411 ( n17160,n16642,n15386 );
   xor U16412 ( n15386,n17184,n16295 );
   not U16413 ( n16295,n17182 );
   nand U16414 ( n17182,n17185,n17186 );
   nand U16415 ( n17159,n16646,n15225 );
   nand U16416 ( p3_u3213,n17187,n17188,n17189,n17190 );
   nor U16417 ( n17190,n17191,n17192,n17193 );
   nor U16418 ( n17193,n15379,n16603 );
   and U16419 ( n15379,n17194,n17195,n17196,n17197 );
   nor U16420 ( n17197,n17198,n17199,n17200,n17201 );
   nor U16421 ( n17201,n16631,n17202,n17203 );
   nor U16422 ( n17200,n15397,n16692 );
   and U16423 ( n17199,n16637,n15381 );
   nor U16424 ( n17198,n15831,n17204,n17205 );
   nor U16425 ( n17196,n17206,n17207 );
   nor U16426 ( n17207,n15828,n17204,n17205 );
   and U16427 ( n17205,n17208,n17209 );
   nand U16428 ( n17209,n17180,n17186 );
   and U16429 ( n17204,n17210,n17186,n17211 );
   nand U16430 ( n17211,n17185,n17212 );
   nor U16431 ( n17206,n16628,n17202,n17203 );
   and U16432 ( n17203,n17208,n17213 );
   nand U16433 ( n17213,n17175,n17186 );
   and U16434 ( n17208,n17214,n17215 );
   and U16435 ( n17202,n17210,n17186,n17216 );
   nand U16436 ( n17216,n17185,n17217 );
   nand U16437 ( n17195,n15381,n16660 );
   nand U16438 ( n17194,n15381,n16705 );
   and U16439 ( n17192,n16603,p3_reg2_reg_20_ );
   nor U16440 ( n17191,n15380,n16640 );
   nand U16441 ( n17189,n16641,n17218 );
   nand U16442 ( n17188,n16642,n15381 );
   xor U16443 ( n15381,n16303,n17219 );
   not U16444 ( n16303,n17210 );
   nand U16445 ( n17210,n17215,n17220 );
   nand U16446 ( n17187,n16646,n15222 );
   nand U16447 ( p3_u3212,n17221,n17222,n17223,n17224 );
   nor U16448 ( n17224,n17225,n17226,n17227 );
   nor U16449 ( n17227,n17228,n16598 );
   and U16450 ( n17226,n15655,n16642 );
   and U16451 ( n17225,n17229,n16641 );
   nand U16452 ( n17223,n16602,n15372 );
   nand U16453 ( n17222,p3_reg2_reg_21_,n16603 );
   nand U16454 ( n17221,n16604,n15656 );
   nand U16455 ( n15656,n17230,n17231,n17232,n17233 );
   nand U16456 ( n17233,n17234,n17235,n17029 );
   nand U16457 ( n17235,n17236,n17237,n17238 );
   nand U16458 ( n17236,n17214,n17217 );
   nand U16459 ( n17234,n17239,n17240 );
   nand U16460 ( n17240,n17175,n17238 );
   not U16461 ( n17175,n17217 );
   nand U16462 ( n17217,n17241,n17157 );
   nand U16463 ( n17241,n17158,n17151 );
   nand U16464 ( n17232,n17242,n17243,n17027 );
   nand U16465 ( n17243,n17244,n17237,n17238 );
   nand U16466 ( n17244,n17214,n17212 );
   nand U16467 ( n17242,n17239,n17245 );
   nand U16468 ( n17245,n17180,n17238 );
   not U16469 ( n17180,n17212 );
   nand U16470 ( n17212,n17246,n17157 );
   nand U16471 ( n17246,n17158,n17147 );
   and U16472 ( n17239,n16302,n17247 );
   nand U16473 ( n17247,n17238,n17248 );
   not U16474 ( n16302,n17237 );
   nand U16475 ( n17231,n15655,n16607 );
   nand U16476 ( n15655,n17249,n17250 );
   nand U16477 ( n17250,n17237,n17251 );
   nand U16478 ( n17237,n17252,n17253 );
   nand U16479 ( n17249,n17254,n17255 );
   nand U16480 ( n17255,n15928,n15877 );
   nand U16481 ( n17230,n16636,n15225 );
   nand U16482 ( p3_u3211,n17256,n17257,n17258,n17259 );
   nor U16483 ( n17259,n17260,n17261,n17262 );
   nor U16484 ( n17262,n17263,n16598 );
   and U16485 ( n17261,n15647,n16642 );
   and U16486 ( n17260,n17264,n16641 );
   nand U16487 ( n17258,n16602,n15366 );
   nand U16488 ( n17257,p3_reg2_reg_22_,n16603 );
   nand U16489 ( n17256,n16604,n15648 );
   nand U16490 ( n15648,n17265,n17266,n17267,n17268 );
   nand U16491 ( n17268,n17269,n17029 );
   xor U16492 ( n17269,n17270,n16298 );
   nand U16493 ( n17267,n17271,n17027 );
   xor U16494 ( n17271,n17272,n16298 );
   nand U16495 ( n17266,n15647,n16607 );
   nand U16496 ( n15647,n17273,n17274 );
   nand U16497 ( n17274,n17275,n16298 );
   nand U16498 ( n16298,n17276,n17277 );
   not U16499 ( n17275,n17278 );
   nand U16500 ( n17273,n17279,n17278 );
   nand U16501 ( n17279,n15878,n17280 );
   nand U16502 ( n17265,n16636,n15222 );
   nand U16503 ( p3_u3210,n17281,n17282,n17283,n17284 );
   nor U16504 ( n17284,n17285,n17286,n17287 );
   nor U16505 ( n17287,n15360,n16603 );
   and U16506 ( n15360,n17288,n17289 );
   nor U16507 ( n17289,n17290,n17291,n17292,n17293 );
   nor U16508 ( n17293,n17294,n16630 );
   nor U16509 ( n17292,n17295,n15828 );
   nor U16510 ( n17291,n17228,n16692 );
   nor U16511 ( n17290,n17294,n16634 );
   nor U16512 ( n17288,n17296,n17297,n17298,n17299 );
   nor U16513 ( n17299,n17300,n16628 );
   nor U16514 ( n17298,n17294,n16923 );
   not U16515 ( n17294,n15356 );
   nor U16516 ( n17297,n17300,n16631 );
   xor U16517 ( n17300,n17301,n17302 );
   nor U16518 ( n17296,n17295,n15831 );
   xor U16519 ( n17295,n17301,n17303 );
   and U16520 ( n17286,n16603,p3_reg2_reg_23_ );
   nor U16521 ( n17285,n17304,n16640 );
   nand U16522 ( n17283,n16641,n17305 );
   nand U16523 ( n17282,n16642,n15356 );
   nand U16524 ( n15356,n17306,n17307 );
   nand U16525 ( n17307,n17308,n15863,n15864 );
   nand U16526 ( n17306,n17301,n17309 );
   nand U16527 ( n17309,n17308,n17280 );
   not U16528 ( n17301,n16299 );
   nand U16529 ( n16299,n17310,n17311 );
   nand U16530 ( n17281,n16646,n15213 );
   nand U16531 ( p3_u3209,n17312,n17313,n17314,n17315 );
   nor U16532 ( n17315,n17316,n17317,n17318 );
   nor U16533 ( n17318,n15349,n16603 );
   and U16534 ( n15349,n17319,n17320 );
   nor U16535 ( n17320,n17321,n17322,n17323,n17324 );
   nor U16536 ( n17324,n17325,n16628 );
   nor U16537 ( n17323,n17326,n15831 );
   nor U16538 ( n17322,n16630,n17327 );
   nor U16539 ( n17321,n17326,n15828 );
   xor U16540 ( n17326,n17328,n17329 );
   nor U16541 ( n17319,n17330,n17331,n17332,n17333 );
   nor U16542 ( n17333,n17263,n16692 );
   nor U16543 ( n17332,n17325,n16631 );
   xor U16544 ( n17325,n17328,n17334 );
   nor U16545 ( n17331,n16923,n17327 );
   nor U16546 ( n17330,n16634,n17327 );
   not U16547 ( n17327,n15351 );
   and U16548 ( n17317,n16603,p3_reg2_reg_24_ );
   nor U16549 ( n17316,n15350,n16640 );
   nand U16550 ( n17314,n16641,n17335 );
   nand U16551 ( n17313,n16642,n15351 );
   xor U16552 ( n15351,n17328,n17336 );
   not U16553 ( n17328,n16300 );
   nand U16554 ( n16300,n17337,n17338 );
   nand U16555 ( n17312,n16646,n15210 );
   nand U16556 ( p3_u3208,n17339,n17340,n17341,n17342 );
   nor U16557 ( n17342,n17343,n17344,n17345 );
   nor U16558 ( n17345,n15339,n16603 );
   and U16559 ( n15339,n17346,n17347,n17348,n17349 );
   nor U16560 ( n17349,n17350,n17351,n17352,n17353 );
   nor U16561 ( n17353,n17354,n16628 );
   nor U16562 ( n17352,n17355,n15828 );
   nor U16563 ( n17351,n16630,n17356 );
   nor U16564 ( n17350,n17354,n16631 );
   xor U16565 ( n17354,n17357,n17358 );
   nor U16566 ( n17348,n17359,n17360 );
   nor U16567 ( n17360,n16634,n17356 );
   not U16568 ( n17356,n15342 );
   nor U16569 ( n17359,n17355,n15831 );
   xor U16570 ( n17355,n17357,n17361 );
   nand U16571 ( n17347,n16636,n15213 );
   nand U16572 ( n17346,n15342,n16637 );
   and U16573 ( n17344,n16603,p3_reg2_reg_25_ );
   nor U16574 ( n17343,n15340,n16640 );
   nand U16575 ( n17341,n16641,n17362 );
   nand U16576 ( n17340,n16642,n15342 );
   xor U16577 ( n15342,n17357,n17363 );
   not U16578 ( n17357,n16301 );
   nand U16579 ( n16301,n17364,n17365 );
   nand U16580 ( n17339,n16646,n15207 );
   nand U16581 ( p3_u3207,n17366,n17367,n17368,n17369 );
   nor U16582 ( n17369,n17370,n17371,n17372 );
   nor U16583 ( n17372,n15617,n16598 );
   nor U16584 ( n17371,n15619,n16599 );
   and U16585 ( n17370,n17373,n16641 );
   nand U16586 ( n17368,n16602,n15329 );
   nand U16587 ( n17367,p3_reg2_reg_26_,n16603 );
   nand U16588 ( n17366,n16604,n15332 );
   nand U16589 ( n15332,n17374,n17375,n17376,n17377 );
   nor U16590 ( n17377,n17378,n17379,n17380,n17381 );
   nor U16591 ( n17381,n16631,n17382,n17383 );
   nor U16592 ( n17380,n16630,n15619 );
   nor U16593 ( n17379,n16923,n15619 );
   nor U16594 ( n17378,n15831,n17384,n17385 );
   nor U16595 ( n17376,n17386,n17387 );
   nor U16596 ( n17387,n15828,n17384,n17385 );
   nor U16597 ( n17385,n17388,n17389 );
   and U16598 ( n17389,n17361,n17365 );
   and U16599 ( n17384,n17390,n17365,n16280 );
   or U16600 ( n17390,n17361,n17391 );
   nand U16601 ( n17361,n17338,n17392 );
   nand U16602 ( n17392,n17337,n17329 );
   nor U16603 ( n17386,n16628,n17382,n17383 );
   nor U16604 ( n17383,n17393,n17388 );
   nand U16605 ( n17388,n17394,n17364 );
   nor U16606 ( n17393,n17395,n17396 );
   not U16607 ( n17396,n17358 );
   nor U16608 ( n17382,n17394,n17395,n17397 );
   nor U16609 ( n17397,n17391,n17358 );
   nand U16610 ( n17358,n17338,n17398 );
   nand U16611 ( n17398,n17334,n17337 );
   not U16612 ( n17395,n17365 );
   nand U16613 ( n17375,n16636,n15210 );
   not U16614 ( n16636,n16692 );
   nand U16615 ( n17374,n15328,n16660 );
   not U16616 ( n16660,n16634 );
   not U16617 ( n15328,n15619 );
   nand U16618 ( n15619,n17399,n17400 );
   nand U16619 ( n17400,n17394,n17401 );
   not U16620 ( n17394,n16280 );
   xor U16621 ( n16280,n17402,n15207 );
   nand U16622 ( n17399,n15855,n15851,n17403 );
   nand U16623 ( p3_u3206,n17404,n17405,n17406,n17407 );
   nor U16624 ( n17407,n17408,n17409,n17410 );
   nor U16625 ( n17410,n15323,n16603 );
   and U16626 ( n15323,n17411,n17412 );
   nor U16627 ( n17412,n17413,n17414,n17415,n17416 );
   nor U16628 ( n17416,n15831,n17417 );
   nor U16629 ( n17415,n17418,n16630 );
   nor U16630 ( n17414,n17418,n16923 );
   nor U16631 ( n17413,n16628,n17419 );
   xor U16632 ( n17419,n16294,n17420 );
   nor U16633 ( n17420,n17421,n17422 );
   nor U16634 ( n17411,n17423,n17424,n17425,n17426 );
   nor U16635 ( n17426,n17427,n16692 );
   nor U16636 ( n17425,n15828,n17417 );
   nand U16637 ( n17417,n17428,n17429,n17430 );
   not U16638 ( n17430,n17431 );
   nand U16639 ( n17429,n17432,n17329 );
   nand U16640 ( n17428,n16294,n17433,n17434 );
   nor U16641 ( n17424,n17418,n16634 );
   not U16642 ( n17418,n15319 );
   nor U16643 ( n17423,n17435,n17436,n16631,n17431 );
   nand U16644 ( n17431,n17437,n17438 );
   nand U16645 ( n17438,n17432,n17439 );
   nand U16646 ( n17437,n16294,n17422 );
   and U16647 ( n17436,n17421,n16294 );
   and U16648 ( n17435,n17334,n17432 );
   nor U16649 ( n17432,n17422,n16294 );
   and U16650 ( n17409,n16603,p3_reg2_reg_27_ );
   nor U16651 ( n17408,n17440,n16640 );
   nand U16652 ( n17406,n16641,n17441 );
   nand U16653 ( n17405,n16642,n15319 );
   nand U16654 ( n15319,n17442,n17443 );
   or U16655 ( n17443,n17444,n16294 );
   nand U16656 ( n17442,n17445,n15855,n16294 );
   and U16657 ( n16294,n17446,n17447 );
   nand U16658 ( n17445,n15851,n17401 );
   nand U16659 ( n17404,n16646,n15201 );
   nand U16660 ( p3_u3205,n17448,n17449,n17450,n17451 );
   nor U16661 ( n17451,n17452,n17453,n17454 );
   nor U16662 ( n17454,n15314,n16603 );
   and U16663 ( n15314,n17455,n17456 );
   nor U16664 ( n17456,n17457,n17458,n17459,n17460 );
   nor U16665 ( n17460,n16628,n17461 );
   nor U16666 ( n17459,n17462,n15831 );
   nor U16667 ( n17458,n17463,n16630 );
   nor U16668 ( n17457,n17462,n15828 );
   xor U16669 ( n17462,n17464,n16296 );
   nor U16670 ( n17455,n17465,n17466,n17467,n17468 );
   nor U16671 ( n17468,n15617,n16692 );
   nor U16672 ( n17467,n16631,n17461 );
   xor U16673 ( n17461,n17469,n16296 );
   nor U16674 ( n17466,n17463,n16923 );
   nor U16675 ( n17465,n17463,n16634 );
   and U16676 ( n17453,n16603,p3_reg2_reg_28_ );
   nor U16677 ( n17452,n17470,n16640 );
   nand U16678 ( n17450,n16641,n17471 );
   nand U16679 ( n17449,n16642,n15309 );
   not U16680 ( n15309,n17463 );
   xor U16681 ( n17463,n16296,n17472 );
   nand U16682 ( n17448,n16646,n15198 );
   not U16683 ( n16646,n16598 );
   nand U16684 ( p3_u3204,n17473,n17474,n17475,n17476 );
   nor U16685 ( n17476,n17477,n17478 );
   nor U16686 ( n17478,n15930,n16640 );
   not U16687 ( n15930,n15304 );
   and U16688 ( n17477,n15303,n16642 );
   nand U16689 ( n16599,n17479,n17480,n16604 );
   nand U16690 ( n17474,p3_reg2_reg_29_,n16603 );
   nand U16691 ( n17473,n16604,n15301 );
   nand U16692 ( n15301,n17481,n17482,n17483,n17484 );
   nor U16693 ( n17484,n17485,n17486,n17487 );
   nor U16694 ( n17487,n17488,n17489,n17490 );
   nor U16695 ( n17490,n17491,n17492 );
   nor U16696 ( n17492,n16780,n17493 );
   nor U16697 ( n17491,n17469,n17494 );
   not U16698 ( n17469,n17495 );
   nor U16699 ( n17486,n17496,n16281 );
   nor U16700 ( n17496,n17497,n17498 );
   nor U16701 ( n17498,n16780,n17499 );
   not U16702 ( n16780,n17029 );
   nor U16703 ( n17497,n17495,n17500,n17494 );
   nor U16704 ( n17494,n17156,n17501 );
   not U16705 ( n17501,n16628 );
   not U16706 ( n17156,n16631 );
   nand U16707 ( n17495,n17502,n17503 );
   nand U16708 ( n17503,n17421,n17446 );
   nor U16709 ( n17421,n17334,n17439 );
   nand U16710 ( n17334,n17311,n17504 );
   nand U16711 ( n17504,n17302,n17310 );
   nand U16712 ( n17302,n17277,n17505 );
   nand U16713 ( n17505,n17270,n17276 );
   and U16714 ( n17270,n17506,n17507 );
   nand U16715 ( n17507,n17508,n17151 );
   nand U16716 ( n17151,n17509,n17510 );
   nand U16717 ( n17510,n17120,n17124 );
   not U16718 ( n17120,n17088 );
   nand U16719 ( n17088,n17065,n17511 );
   nand U16720 ( n17511,n17058,n17064 );
   nand U16721 ( n17058,n17041,n17512 );
   nand U16722 ( n17512,n17036,n17040 );
   not U16723 ( n17036,n17030 );
   nand U16724 ( n17030,n17513,n17514 );
   nand U16725 ( n17513,n16996,n17002 );
   nor U16726 ( n16996,n16939,n16921 );
   and U16727 ( n16921,n17515,n17516 );
   nand U16728 ( n17516,n16900,n17517 );
   nand U16729 ( n17517,n17518,n16901,n16874 );
   nor U16730 ( n17485,n17519,n16692 );
   nand U16731 ( n17483,n15303,n16607 );
   nand U16732 ( n16607,n17521,n16923 );
   not U16733 ( n16923,n16637 );
   nor U16734 ( n16637,n16172,n17522 );
   not U16735 ( n17521,n16839 );
   nand U16736 ( n16839,n16630,n16634 );
   nand U16737 ( n15303,n17523,n17524 );
   nand U16738 ( n17524,n17488,n17525 );
   nand U16739 ( n17525,n15845,n17526 );
   nand U16740 ( n17526,n17472,n15848 );
   not U16741 ( n17488,n16281 );
   nand U16742 ( n17523,n16281,n17527 );
   nand U16743 ( n17527,n15848,n17528 );
   nand U16744 ( n17528,n17529,n15845 );
   not U16745 ( n17529,n17472 );
   nand U16746 ( n17472,n15852,n17530 );
   nand U16747 ( n17530,n17444,n15847 );
   nand U16748 ( n15847,n15617,n15320 );
   nand U16749 ( n17444,n15851,n17531 );
   nand U16750 ( n17531,n17403,n15855 );
   nand U16751 ( n15855,n17427,n15329 );
   not U16752 ( n17403,n17401 );
   nand U16753 ( n17401,n15856,n17532 );
   nand U16754 ( n17532,n17363,n15858 );
   nand U16755 ( n15858,n15340,n15210 );
   nand U16756 ( n17363,n15859,n17533 );
   nand U16757 ( n17533,n15862,n17336 );
   nand U16758 ( n17336,n17534,n15863 );
   nand U16759 ( n15863,n17263,n15357 );
   nand U16760 ( n17534,n15864,n17308 );
   nand U16761 ( n17308,n15878,n17278 );
   nand U16762 ( n17278,n17535,n15928 );
   nand U16763 ( n15928,n17536,n15222 );
   nand U16764 ( n17535,n17254,n15877 );
   nand U16765 ( n15877,n17537,n15372 );
   not U16766 ( n17254,n17251 );
   nand U16767 ( n17251,n17538,n17539 );
   nand U16768 ( n17539,n17540,n15661 );
   or U16769 ( n17540,n17219,n17541 );
   nand U16770 ( n17538,n17541,n17219 );
   nand U16771 ( n17219,n17542,n17543 );
   nand U16772 ( n17543,n15924,n17184 );
   nand U16773 ( n17184,n17544,n17545 );
   nand U16774 ( n17545,n17546,n15401 );
   or U16775 ( n17546,n17154,n15409 );
   nand U16776 ( n17544,n15409,n17154 );
   nand U16777 ( n17154,n17547,n17548 );
   nand U16778 ( n17548,n17549,n15411 );
   nand U16779 ( n17549,n15234,n17128 );
   or U16780 ( n17547,n17128,n15234 );
   nand U16781 ( n17128,n17550,n17551 );
   nand U16782 ( n17551,n15883,n17552 );
   nand U16783 ( n17552,n17096,n17553 );
   nand U16784 ( n17553,n17101,n15887 );
   not U16785 ( n17101,n15890 );
   nand U16786 ( n15890,n17554,n15243 );
   and U16787 ( n17096,n15886,n15881 );
   nand U16788 ( n15881,n17091,n15237 );
   nand U16789 ( n15886,n17555,n15240 );
   nand U16790 ( n17550,n15883,n15887,n17100 );
   nor U16791 ( n17100,n17039,n17556 );
   nand U16792 ( n17039,n15891,n17557 );
   nand U16793 ( n17557,n17009,n15897 );
   nand U16794 ( n15897,n17007,n15246 );
   nand U16795 ( n17009,n15920,n17558 );
   nand U16796 ( n17558,n16968,n15898 );
   nand U16797 ( n15898,n16966,n15249 );
   and U16798 ( n16968,n17559,n17560 );
   nand U16799 ( n17560,n15899,n15923,n16941 );
   and U16800 ( n16941,n16871,n15900 );
   nand U16801 ( n15900,n15487,n15480 );
   nand U16802 ( n16871,n17561,n17562 );
   nand U16803 ( n17562,n17563,n15261 );
   nand U16804 ( n17563,n16838,n15489 );
   not U16805 ( n16838,n16845 );
   nand U16806 ( n17561,n15904,n16845 );
   nand U16807 ( n16845,n15910,n16813 );
   nand U16808 ( n16813,n15906,n16852 );
   nand U16809 ( n16852,n17564,n17565 );
   nand U16810 ( n17565,n17566,n15912 );
   nand U16811 ( n17566,n15917,n17567 );
   or U16812 ( n17567,n16733,n15914 );
   not U16813 ( n15914,n16759 );
   nand U16814 ( n16733,n17568,n15273 );
   and U16815 ( n15917,n16758,n15915 );
   nand U16816 ( n15915,n17569,n15267 );
   nand U16817 ( n16758,n17570,n15270 );
   nand U16818 ( n17564,n16730,n16732,n16759,n15912 );
   nand U16819 ( n15912,n16741,n15509 );
   nand U16820 ( n16759,n16718,n15516 );
   nand U16821 ( n16732,n17571,n15522 );
   not U16822 ( n16730,n16727 );
   nand U16823 ( n16727,n17572,n17573 );
   nand U16824 ( n17573,n15783,n15528 );
   nand U16825 ( n17572,n16700,n17574 );
   nand U16826 ( n17574,n16707,n15276 );
   and U16827 ( n16700,n16662,n16669 );
   nand U16828 ( n16669,n16663,n16661 );
   nand U16829 ( n16661,n16691,n15538 );
   not U16830 ( n16663,n16667 );
   nand U16831 ( n16667,n17575,n17576 );
   nand U16832 ( n17576,n17577,n15548 );
   nand U16833 ( n17577,n15282,n16643 );
   or U16834 ( n17575,n15282,n16643 );
   nand U16835 ( n16662,n16673,n15279 );
   not U16836 ( n16673,n15538 );
   nand U16837 ( n15906,n15507,n15496 );
   nand U16838 ( n15910,n17578,n15264 );
   nand U16839 ( n17559,n15918,n15923 );
   nand U16840 ( n15923,n16883,n15464 );
   nand U16841 ( n15918,n16937,n17579 );
   nand U16842 ( n17579,n16942,n15899 );
   nand U16843 ( n15899,n16860,n15474 );
   not U16844 ( n16942,n16872 );
   nand U16845 ( n16872,n17580,n15258 );
   and U16846 ( n16937,n16904,n17581 );
   nand U16847 ( n17581,n16932,n15252 );
   nand U16848 ( n15920,n16985,n15454 );
   nand U16849 ( n15891,n17582,n15444 );
   nand U16850 ( n15887,n15435,n15428 );
   nand U16851 ( n15883,n17051,n15418 );
   nand U16852 ( n15924,n15874,n15228 );
   nand U16853 ( n17542,n15397,n15387 );
   nand U16854 ( n15878,n17228,n15366 );
   and U16855 ( n15864,n17280,n17583 );
   nand U16856 ( n17583,n17304,n15216 );
   nand U16857 ( n17280,n17584,n15219 );
   nand U16858 ( n15862,n15350,n15213 );
   nand U16859 ( n15851,n17402,n15207 );
   nand U16860 ( n15852,n17440,n15204 );
   nand U16861 ( n17482,n17585,n15195,n15559 );
   nand U16862 ( n15195,n17586,n17587,n17588,n17589 );
   nand U16863 ( n17588,p3_reg2_reg_30_,n17590 );
   nand U16864 ( n17587,p3_reg1_reg_30_,n17591 );
   nand U16865 ( n17586,p3_reg0_reg_30_,n17592 );
   nand U16866 ( n17481,n17593,n17027 );
   xor U16867 ( n17593,n16281,n17594 );
   nand U16868 ( n17594,n17499,n17595 );
   nand U16869 ( n17595,n17464,n17493 );
   and U16870 ( n17464,n17502,n17596 );
   nand U16871 ( n17596,n17434,n17446,n17433 );
   not U16872 ( n17433,n17439 );
   nand U16873 ( n17439,n17597,n17338 );
   not U16874 ( n17434,n17329 );
   nand U16875 ( n17329,n17311,n17598 );
   nand U16876 ( n17598,n17310,n17303 );
   nand U16877 ( n17303,n17277,n17599 );
   nand U16878 ( n17599,n17272,n17276 );
   nand U16879 ( n17276,n15366,n15219 );
   and U16880 ( n17272,n17506,n17600 );
   nand U16881 ( n17600,n17508,n17147 );
   nand U16882 ( n17147,n17509,n17601 );
   nand U16883 ( n17601,n17124,n17127 );
   not U16884 ( n17127,n17089 );
   nand U16885 ( n17089,n17065,n17602 );
   nand U16886 ( n17602,n17064,n17060 );
   nand U16887 ( n17060,n17041,n17603 );
   nand U16888 ( n17603,n17035,n17040 );
   nand U16889 ( n17040,n15437,n15243 );
   not U16890 ( n17035,n17028 );
   nand U16891 ( n17028,n17604,n17514 );
   nand U16892 ( n17514,n17605,n17010 );
   nand U16893 ( n17605,n16970,n17003,n17606 );
   nand U16894 ( n17606,n17002,n16940 );
   nor U16895 ( n16940,n16932,n16883 );
   nand U16896 ( n17003,n15444,n15246 );
   nand U16897 ( n16970,n15454,n15249 );
   nand U16898 ( n17604,n17005,n17002 );
   and U16899 ( n17002,n17010,n16969 );
   nand U16900 ( n16969,n16985,n16966 );
   nand U16901 ( n17010,n17582,n17007 );
   nor U16902 ( n17005,n16939,n16925 );
   not U16903 ( n16925,n16930 );
   nand U16904 ( n16930,n16901,n17515,n17607 );
   nand U16905 ( n17607,n17608,n16900 );
   nand U16906 ( n17608,n17518,n16874 );
   nand U16907 ( n16874,n15480,n15258 );
   nand U16908 ( n17518,n16850,n16875 );
   nor U16909 ( n16850,n15904,n15908 );
   nand U16910 ( n17515,n16900,n16875,n16895 );
   and U16911 ( n16895,n16840,n17609 );
   nand U16912 ( n17609,n15908,n15904 );
   not U16913 ( n15904,n15489 );
   not U16914 ( n16840,n16846 );
   nand U16915 ( n16846,n17610,n16820 );
   nand U16916 ( n16820,n17578,n15507 );
   nand U16917 ( n17610,n17611,n16786,n16821 );
   nand U16918 ( n16821,n15496,n15264 );
   nand U16919 ( n16786,n15267,n15509 );
   nand U16920 ( n17611,n17612,n16787 );
   nand U16921 ( n16787,n17569,n16741 );
   not U16922 ( n17612,n16782 );
   nand U16923 ( n16782,n17613,n16754 );
   nand U16924 ( n16754,n16718,n17570 );
   not U16925 ( n17570,n15516 );
   nand U16926 ( n17613,n17614,n16728,n16755 );
   nand U16927 ( n16755,n15516,n15270 );
   nand U16928 ( n16728,n15522,n15273 );
   nand U16929 ( n17614,n16751,n16729 );
   nand U16930 ( n16729,n17571,n17568 );
   nand U16931 ( n16751,n17615,n17616 );
   nand U16932 ( n17616,n17617,n17618 );
   nand U16933 ( n17618,n16707,n15783 );
   or U16934 ( n17617,n16704,n16703 );
   nor U16935 ( n16703,n16675,n17619 );
   nor U16936 ( n17619,n15538,n15279 );
   nand U16937 ( n16675,n16635,n16645 );
   nand U16938 ( n16645,n16639,n15796 );
   not U16939 ( n16635,n16610 );
   nand U16940 ( n16704,n17620,n17621 );
   nand U16941 ( n17621,n17622,n15538 );
   nand U16942 ( n17622,n16691,n16644 );
   or U16943 ( n17620,n16644,n16691 );
   nand U16944 ( n16644,n15548,n15282 );
   nand U16945 ( n17615,n15528,n15276 );
   nand U16946 ( n16875,n17580,n15487 );
   nand U16947 ( n16900,n17623,n16860 );
   nor U16948 ( n16939,n15464,n15252 );
   nand U16949 ( n17064,n15428,n15240 );
   nand U16950 ( n17065,n15435,n17555 );
   not U16951 ( n15435,n15240 );
   and U16952 ( n17124,n17624,n17098 );
   nand U16953 ( n17098,n17051,n17091 );
   nand U16954 ( n17624,n15873,n17129 );
   nand U16955 ( n17509,n17625,n17626 );
   nand U16956 ( n17626,n15873,n17627 );
   or U16957 ( n17627,n17099,n17129 );
   nand U16958 ( n17625,n17129,n17099 );
   nand U16959 ( n17099,n15418,n15237 );
   and U16960 ( n17508,n17158,n17253,n17214 );
   not U16961 ( n17214,n17248 );
   nand U16962 ( n17158,n15926,n15409 );
   not U16963 ( n15926,n15401 );
   and U16964 ( n17506,n17628,n17252 );
   nand U16965 ( n17252,n15372,n15222 );
   nand U16966 ( n17628,n17253,n17629 );
   nand U16967 ( n17629,n17238,n17630 );
   or U16968 ( n17630,n17157,n17248 );
   nand U16969 ( n17248,n17185,n17220 );
   nand U16970 ( n17185,n15397,n15874 );
   nand U16971 ( n17157,n15401,n15231 );
   and U16972 ( n17238,n17215,n17631 );
   nand U16973 ( n17631,n17632,n17220 );
   nand U16974 ( n17220,n15380,n17541 );
   not U16975 ( n15380,n15661 );
   not U16976 ( n17632,n17186 );
   nand U16977 ( n17186,n15387,n15228 );
   nand U16978 ( n17215,n15661,n15225 );
   nand U16979 ( n17253,n17537,n17536 );
   nand U16980 ( n17277,n17228,n17584 );
   not U16981 ( n17228,n15219 );
   nand U16982 ( n17310,n15357,n15216 );
   nand U16983 ( n17311,n17304,n17263 );
   and U16984 ( n17502,n17447,n17633 );
   nand U16985 ( n17633,n17422,n17446 );
   nand U16986 ( n17446,n17440,n15617 );
   nand U16987 ( n17422,n17634,n17635 );
   nand U16988 ( n17635,n17597,n17636 );
   nand U16989 ( n17636,n17365,n17337 );
   nand U16990 ( n17337,n15632,n15213 );
   nand U16991 ( n17365,n15625,n15210 );
   and U16992 ( n17597,n17364,n17637 );
   nand U16993 ( n17637,n17402,n17427 );
   nand U16994 ( n17634,n15329,n15207 );
   nand U16995 ( n17447,n15320,n15204 );
   xor U16996 ( n16281,n15844,n15304 );
   nand U16997 ( n15304,n17638,n17639 );
   nand U16998 ( n17639,n16562,n17640 );
   xor U16999 ( n16562,n17641,n17642 );
   xor U17000 ( n17641,p2_datao_reg_29_,p1_datao_reg_29_ );
   nand U17001 ( n17638,si_29_,n17643 );
   not U17002 ( n15844,n15198 );
   nand U17003 ( p3_u3203,n17644,n17645,n17646 );
   nand U17004 ( n17645,n16602,n15296 );
   nand U17005 ( n15296,n17647,n17648 );
   nand U17006 ( n17648,n17640,n16571 );
   xor U17007 ( n16571,n17649,n17650 );
   xor U17008 ( n17649,p2_datao_reg_30_,p1_datao_reg_30_ );
   nand U17009 ( n17647,si_30_,n17643 );
   nand U17010 ( n17644,p3_reg2_reg_30_,n16603 );
   nand U17011 ( p3_u3202,n17651,n17652,n17646 );
   and U17012 ( n17646,n17475,n17653 );
   nand U17013 ( n17653,n16604,n15294 );
   and U17014 ( n15294,n17585,n15192,n15559 );
   nand U17015 ( n15192,n17654,n17655,n17656,n17589 );
   nand U17016 ( n17656,p3_reg2_reg_31_,n17590 );
   nand U17017 ( n17655,p3_reg1_reg_31_,n17591 );
   nand U17018 ( n17654,p3_reg0_reg_31_,n17592 );
   nand U17019 ( n17585,n17657,n17658 );
   nand U17020 ( n17658,n17659,n17660 );
   nand U17021 ( n17475,n16641,n17661 );
   nand U17022 ( n17652,n16602,n15291 );
   nand U17023 ( n15291,n17663,n17664 );
   nand U17024 ( n17664,n16579,n17657 );
   nand U17025 ( n16579,n17665,n17666 );
   nand U17026 ( n17666,n16576,n17667,n17668 );
   xor U17027 ( n17668,p2_datao_reg_31_,n17669 );
   nand U17028 ( n17667,n17670,n17671 );
   nand U17029 ( n17665,n17672,n16576,n17670,n17671 );
   nand U17030 ( n17671,n17650,n17673 );
   or U17031 ( n17673,n17674,p2_datao_reg_30_ );
   and U17032 ( n17650,n17675,n17676 );
   nand U17033 ( n17676,n17677,n17678 );
   nand U17034 ( n17677,n17679,n17642 );
   or U17035 ( n17675,n17679,n17642 );
   nand U17036 ( n17642,n17680,n17681 );
   nand U17037 ( n17681,p2_datao_reg_28_,n17682 );
   or U17038 ( n17682,n17683,n17684 );
   nand U17039 ( n17680,n17684,n17683 );
   nand U17040 ( n17670,p2_datao_reg_30_,n17674 );
   xor U17041 ( n17672,p2_datao_reg_31_,p1_datao_reg_31_ );
   nand U17042 ( n17663,si_31_,n17643 );
   nand U17043 ( n17651,p3_reg2_reg_31_,n16603 );
   nand U17044 ( n17686,n17662,n17687 );
   nand U17045 ( n17687,n17688,n17689,n15566 );
   nand U17046 ( n17689,n17690,n15582 );
   nand U17047 ( n17690,n15583,n17691 );
   nand U17048 ( n17691,n17692,n15580,n15943 );
   nand U17049 ( n17692,n17480,n15809 );
   nand U17050 ( n17688,n15570,n17693 );
   nand U17051 ( n17693,n15584,n15572 );
   nand U17052 ( n15584,n17694,n17695 );
   nand U17053 ( n17694,n17479,n16260 );
   nand U17054 ( p3_u3201,n17696,n17697,n17698,n17699 );
   nor U17055 ( n17699,n17700,n17701,n17702 );
   nor U17056 ( n17702,n17703,n17704 );
   nor U17057 ( n17701,n15577,n17705 );
   nand U17058 ( n17698,n17706,n17707,n17708 );
   nand U17059 ( n17707,n17709,n17710,n17711 );
   not U17060 ( n17711,n17712 );
   nand U17061 ( n17709,p3_reg2_reg_18_,n17713 );
   nand U17062 ( n17706,n17714,n17713,n17712 );
   or U17063 ( n17713,n17715,n17716 );
   nand U17064 ( n17714,n17710,n17717 );
   nand U17065 ( n17710,n17716,n17715 );
   nand U17066 ( n17697,n17718,n17719 );
   xor U17067 ( n17718,n17720,n17721 );
   nand U17068 ( n17721,n17722,n17723 );
   nand U17069 ( n17723,n17724,n17725 );
   or U17070 ( n17725,n17726,n17727 );
   nand U17071 ( n17722,n17727,n17726 );
   nand U17072 ( n17720,n17728,n17729 );
   nand U17073 ( n17729,n17730,n15937 );
   nand U17074 ( n17728,n17712,n17731 );
   xor U17075 ( n17712,p3_reg2_reg_19_,n17480 );
   nand U17076 ( n17696,n17732,n17733,n17734 );
   nand U17077 ( n17733,n17735,n17736,n17737 );
   not U17078 ( n17737,n17730 );
   nand U17079 ( n17735,p3_reg1_reg_18_,n17738 );
   nand U17080 ( n17732,n17739,n17738,n17730 );
   xor U17081 ( n17730,p3_reg1_reg_19_,n17480 );
   or U17082 ( n17738,n17740,n17716 );
   nand U17083 ( n17739,n17736,n17741 );
   nand U17084 ( n17736,n17716,n17740 );
   nand U17085 ( p3_u3200,n17742,n17743,n17744,n17745 );
   nand U17086 ( n17745,n17724,n17746 );
   nand U17087 ( n17746,n17705,n17747,n17748,n17749 );
   nand U17088 ( n17749,n17750,n17719 );
   nand U17089 ( n17748,n17734,n17751 );
   xor U17090 ( n17751,n17740,n17741 );
   nand U17091 ( n17747,n17708,n17752 );
   xor U17092 ( n17752,n17715,n17717 );
   nand U17093 ( n17744,n17753,n17716 );
   nand U17094 ( n17753,n17754,n17755,n17756 );
   nand U17095 ( n17756,n17757,n17708 );
   xor U17096 ( n17757,p3_reg2_reg_18_,n17715 );
   nand U17097 ( n17715,n17758,n17759 );
   nand U17098 ( n17759,p3_reg2_reg_17_,n17760 );
   or U17099 ( n17760,n17761,n17762 );
   nand U17100 ( n17758,n17761,n17762 );
   or U17101 ( n17755,n17763,n17750 );
   xor U17102 ( n17750,n17727,n17726 );
   nand U17103 ( n17726,n17764,n17765 );
   nand U17104 ( n17765,n17766,n17767 );
   or U17105 ( n17767,n17768,n17769 );
   nand U17106 ( n17764,n17769,n17768 );
   nand U17107 ( n17727,n17770,n17771 );
   nand U17108 ( n17771,n17731,n17717 );
   not U17109 ( n17717,p3_reg2_reg_18_ );
   nand U17110 ( n17770,n15937,n17741 );
   not U17111 ( n17741,p3_reg1_reg_18_ );
   nand U17112 ( n17754,n17772,n17734 );
   xor U17113 ( n17772,p3_reg1_reg_18_,n17740 );
   nand U17114 ( n17740,n17773,n17774 );
   nand U17115 ( n17774,p3_reg1_reg_17_,n17775 );
   or U17116 ( n17775,n17776,n17762 );
   nand U17117 ( n17773,n17776,n17762 );
   nand U17118 ( n17743,n17777,p3_addr_reg_18_ );
   nand U17119 ( n17742,p3_reg3_reg_18_,p3_u3151 );
   nand U17120 ( p3_u3199,n17778,n17779,n17780,n17781 );
   nand U17121 ( n17781,n17766,n17782 );
   nand U17122 ( n17782,n17705,n17783,n17784,n17785 );
   nand U17123 ( n17785,n17786,n17719 );
   nand U17124 ( n17784,n17734,n17787 );
   xor U17125 ( n17787,n17776,n17788 );
   nand U17126 ( n17783,n17708,n17789 );
   xor U17127 ( n17789,n17761,n17790 );
   nand U17128 ( n17780,n17791,n17762 );
   nand U17129 ( n17791,n17792,n17793,n17794 );
   nand U17130 ( n17794,n17795,n17708 );
   xor U17131 ( n17795,p3_reg2_reg_17_,n17761 );
   nand U17132 ( n17761,n17796,n17797 );
   nand U17133 ( n17797,p3_reg2_reg_16_,n17798 );
   or U17134 ( n17798,n17799,n17800 );
   nand U17135 ( n17796,n17800,n17799 );
   or U17136 ( n17793,n17763,n17786 );
   xor U17137 ( n17786,n17769,n17768 );
   nand U17138 ( n17768,n17801,n17802 );
   nand U17139 ( n17801,n17803,n17804 );
   nand U17140 ( n17769,n17805,n17806 );
   nand U17141 ( n17806,n17731,n17790 );
   not U17142 ( n17790,p3_reg2_reg_17_ );
   nand U17143 ( n17805,n15937,n17788 );
   not U17144 ( n17788,p3_reg1_reg_17_ );
   nand U17145 ( n17792,n17807,n17734 );
   xor U17146 ( n17807,p3_reg1_reg_17_,n17776 );
   nand U17147 ( n17776,n17808,n17809 );
   nand U17148 ( n17809,p3_reg1_reg_16_,n17810 );
   or U17149 ( n17810,n17811,n17800 );
   nand U17150 ( n17808,n17800,n17811 );
   nand U17151 ( n17779,n17777,p3_addr_reg_17_ );
   nand U17152 ( n17778,p3_reg3_reg_17_,p3_u3151 );
   nand U17153 ( p3_u3198,n17812,n17813,n17814 );
   nor U17154 ( n17814,n17815,n17816,n17817 );
   nor U17155 ( n17817,n17818,n17800 );
   nor U17156 ( n17818,n17819,n17820,n17821 );
   nor U17157 ( n17821,n17822,n17823 );
   xor U17158 ( n17822,p3_reg2_reg_16_,n17799 );
   nor U17159 ( n17820,n17824,n17825 );
   xor U17160 ( n17824,p3_reg1_reg_16_,n17811 );
   nor U17161 ( n17816,n17826,n17827 );
   nor U17162 ( n17826,n17828,n17829 );
   nor U17163 ( n17829,n17823,n17830 );
   xor U17164 ( n17830,n17799,n17090 );
   nand U17165 ( n17799,n17831,n17832 );
   nand U17166 ( n17832,p3_reg2_reg_15_,n17833 );
   or U17167 ( n17833,n17834,n17835 );
   nand U17168 ( n17831,n17834,n17835 );
   nor U17169 ( n17828,n17825,n17836 );
   xor U17170 ( n17836,n17811,n15421 );
   nand U17171 ( n17811,n17837,n17838 );
   nand U17172 ( n17838,p3_reg1_reg_15_,n17839 );
   or U17173 ( n17839,n17840,n17835 );
   nand U17174 ( n17837,n17840,n17835 );
   nand U17175 ( n17813,n17719,n17841 );
   nand U17176 ( n17841,n17842,n17843 );
   nand U17177 ( n17843,n17804,n17802,n17803 );
   and U17178 ( n17803,n17844,n17845 );
   or U17179 ( n17845,n17846,n17827 );
   nand U17180 ( n17802,n17827,n17846 );
   nand U17181 ( n17804,n17847,n17848 );
   nand U17182 ( n17842,n17849,n17847,n17850 );
   xor U17183 ( n17850,n17800,n17846 );
   nand U17184 ( n17846,n17851,n17852 );
   nand U17185 ( n17852,n17731,n17090 );
   not U17186 ( n17090,p3_reg2_reg_16_ );
   nand U17187 ( n17851,n15937,n15421 );
   not U17188 ( n15421,p3_reg1_reg_16_ );
   nand U17189 ( n17849,n17853,n17844 );
   nand U17190 ( n17844,n17854,n17835 );
   nand U17191 ( n17812,n17777,p3_addr_reg_16_ );
   nand U17192 ( p3_u3197,n17855,n17856,n17857,n17858 );
   nor U17193 ( n17858,n17859,n17860 );
   and U17194 ( n17860,p3_addr_reg_15_,n17777 );
   nor U17195 ( n17859,n17847,n17853,n17763 );
   nand U17196 ( n17847,n17861,n17862 );
   nand U17197 ( n17857,p3_reg3_reg_15_,p3_u3151 );
   nand U17198 ( n17856,n17863,n17835 );
   nand U17199 ( n17863,n17864,n17865,n17866 );
   nand U17200 ( n17866,n17867,n17708 );
   xor U17201 ( n17867,p3_reg2_reg_15_,n17834 );
   nand U17202 ( n17865,n17868,n17719 );
   xor U17203 ( n17868,n17853,n17854 );
   nand U17204 ( n17864,n17869,n17734 );
   xor U17205 ( n17869,p3_reg1_reg_15_,n17840 );
   nand U17206 ( n17855,n17861,n17870 );
   nand U17207 ( n17870,n17705,n17871,n17872,n17873 );
   nand U17208 ( n17873,n17854,n17719,n17853 );
   not U17209 ( n17853,n17848 );
   nand U17210 ( n17848,n17874,n17875 );
   nand U17211 ( n17875,n17876,n17877 );
   nand U17212 ( n17877,n17878,n17879 );
   nand U17213 ( n17874,n17880,n17881 );
   not U17214 ( n17854,n17862 );
   nand U17215 ( n17862,n17882,n17883 );
   nand U17216 ( n17883,n17731,n17884 );
   nand U17217 ( n17882,n15937,n17885 );
   nand U17218 ( n17872,n17734,n17886 );
   xor U17219 ( n17886,n17840,n17885 );
   not U17220 ( n17885,p3_reg1_reg_15_ );
   nand U17221 ( n17840,n17887,n17888 );
   nand U17222 ( n17888,p3_reg1_reg_14_,n17889 );
   or U17223 ( n17889,n17890,n17881 );
   nand U17224 ( n17887,n17881,n17890 );
   nand U17225 ( n17871,n17708,n17891 );
   xor U17226 ( n17891,n17834,n17884 );
   not U17227 ( n17884,p3_reg2_reg_15_ );
   nand U17228 ( n17834,n17892,n17893 );
   nand U17229 ( n17893,p3_reg2_reg_14_,n17894 );
   or U17230 ( n17894,n17895,n17881 );
   nand U17231 ( n17892,n17881,n17895 );
   nand U17232 ( p3_u3196,n17896,n17897,n17898,n17899 );
   nand U17233 ( n17899,n17881,n17900 );
   nand U17234 ( n17900,n17901,n17902,n17903 );
   nand U17235 ( n17903,n17904,n17708 );
   xor U17236 ( n17904,p3_reg2_reg_14_,n17895 );
   nand U17237 ( n17902,n17719,n17905 );
   xor U17238 ( n17905,n17879,n17876 );
   nand U17239 ( n17901,n17906,n17734 );
   xor U17240 ( n17906,p3_reg1_reg_14_,n17890 );
   nand U17241 ( n17898,n17878,n17907 );
   nand U17242 ( n17907,n17705,n17908,n17909,n17910 );
   nand U17243 ( n17910,n17911,n17719 );
   xor U17244 ( n17911,n17880,n17876 );
   and U17245 ( n17876,n17912,n17913 );
   nand U17246 ( n17913,n17914,n17915 );
   or U17247 ( n17915,n17916,n17917 );
   nand U17248 ( n17912,n17917,n17916 );
   not U17249 ( n17880,n17879 );
   nand U17250 ( n17879,n17918,n17919 );
   nand U17251 ( n17919,n17731,n17920 );
   nand U17252 ( n17918,n15937,n17921 );
   nand U17253 ( n17909,n17734,n17922 );
   xor U17254 ( n17922,n17890,n17921 );
   not U17255 ( n17921,p3_reg1_reg_14_ );
   nand U17256 ( n17890,n17923,n17924 );
   nand U17257 ( n17924,p3_reg1_reg_13_,n17925 );
   or U17258 ( n17925,n17926,n17927 );
   nand U17259 ( n17923,n17926,n17927 );
   nand U17260 ( n17908,n17708,n17928 );
   xor U17261 ( n17928,n17895,n17920 );
   not U17262 ( n17920,p3_reg2_reg_14_ );
   nand U17263 ( n17895,n17929,n17930 );
   nand U17264 ( n17930,p3_reg2_reg_13_,n17931 );
   or U17265 ( n17931,n17932,n17927 );
   nand U17266 ( n17929,n17932,n17927 );
   nand U17267 ( n17897,n17777,p3_addr_reg_14_ );
   nand U17268 ( n17896,p3_reg3_reg_14_,p3_u3151 );
   nand U17269 ( p3_u3195,n17933,n17934,n17935,n17936 );
   nand U17270 ( n17936,n17914,n17937 );
   nand U17271 ( n17937,n17705,n17938,n17939,n17940 );
   nand U17272 ( n17940,n17941,n17719 );
   nand U17273 ( n17939,n17734,n17942 );
   xor U17274 ( n17942,n17926,n15447 );
   nand U17275 ( n17938,n17708,n17943 );
   xor U17276 ( n17943,n17932,n17006 );
   nand U17277 ( n17935,n17944,n17927 );
   nand U17278 ( n17944,n17945,n17946,n17947 );
   nand U17279 ( n17947,n17948,n17708 );
   xor U17280 ( n17948,p3_reg2_reg_13_,n17932 );
   nand U17281 ( n17932,n17949,n17950 );
   nand U17282 ( n17950,p3_reg2_reg_12_,n17951 );
   or U17283 ( n17951,n17952,n17953 );
   nand U17284 ( n17949,n17953,n17952 );
   or U17285 ( n17946,n17763,n17941 );
   xor U17286 ( n17941,n17917,n17916 );
   nand U17287 ( n17916,n17954,n17955 );
   nand U17288 ( n17955,n17956,n17957 );
   nand U17289 ( n17957,n17958,n17959 );
   or U17290 ( n17954,n17959,n17958 );
   nand U17291 ( n17917,n17960,n17961 );
   nand U17292 ( n17961,n17731,n17006 );
   not U17293 ( n17006,p3_reg2_reg_13_ );
   nand U17294 ( n17960,n15937,n15447 );
   not U17295 ( n15447,p3_reg1_reg_13_ );
   nand U17296 ( n17945,n17962,n17734 );
   xor U17297 ( n17962,p3_reg1_reg_13_,n17926 );
   nand U17298 ( n17926,n17963,n17964 );
   nand U17299 ( n17964,p3_reg1_reg_12_,n17965 );
   or U17300 ( n17965,n17966,n17953 );
   nand U17301 ( n17963,n17953,n17966 );
   nand U17302 ( n17934,n17777,p3_addr_reg_13_ );
   nand U17303 ( n17933,p3_reg3_reg_13_,p3_u3151 );
   nand U17304 ( p3_u3194,n17967,n17968,n17969,n17970 );
   nand U17305 ( n17970,n17953,n17971 );
   nand U17306 ( n17971,n17972,n17973,n17974 );
   nand U17307 ( n17974,n17975,n17708 );
   xor U17308 ( n17975,p3_reg2_reg_12_,n17952 );
   nand U17309 ( n17973,n17976,n17719 );
   xor U17310 ( n17976,n17959,n17977 );
   nand U17311 ( n17972,n17978,n17734 );
   xor U17312 ( n17978,p3_reg1_reg_12_,n17966 );
   nand U17313 ( n17969,n17956,n17979 );
   nand U17314 ( n17979,n17705,n17980,n17981,n17982 );
   nand U17315 ( n17982,n17719,n17983 );
   xor U17316 ( n17983,n17959,n17958 );
   not U17317 ( n17958,n17977 );
   nand U17318 ( n17977,n17984,n17985 );
   nand U17319 ( n17985,n17731,n16965 );
   nand U17320 ( n17984,n15937,n15457 );
   nand U17321 ( n17959,n17986,n17987 );
   nand U17322 ( n17987,n17988,n17989,n17990 );
   not U17323 ( n17990,n17991 );
   nand U17324 ( n17986,n17992,n17989 );
   nand U17325 ( n17992,n17993,n17994 );
   nand U17326 ( n17994,n17988,n17995,n17996 );
   nand U17327 ( n17981,n17734,n17997 );
   xor U17328 ( n17997,n17966,n15457 );
   not U17329 ( n15457,p3_reg1_reg_12_ );
   nand U17330 ( n17966,n17998,n17999 );
   nand U17331 ( n17999,p3_reg1_reg_11_,n18000 );
   or U17332 ( n18000,n18001,n18002 );
   nand U17333 ( n17998,n18001,n18002 );
   nand U17334 ( n17980,n17708,n18003 );
   xor U17335 ( n18003,n17952,n16965 );
   not U17336 ( n16965,p3_reg2_reg_12_ );
   nand U17337 ( n17952,n18004,n18005 );
   nand U17338 ( n18005,p3_reg2_reg_11_,n18006 );
   or U17339 ( n18006,n18007,n18002 );
   nand U17340 ( n18004,n18007,n18002 );
   nand U17341 ( n17968,n17777,p3_addr_reg_12_ );
   nand U17342 ( n17967,p3_reg3_reg_12_,p3_u3151 );
   nand U17343 ( p3_u3193,n18008,n18009,n18010 );
   nor U17344 ( n18010,n18011,n18012,n18013 );
   nor U17345 ( n18013,n18014,n18015 );
   nor U17346 ( n18015,n18016,n18017 );
   nor U17347 ( n18017,n17823,n18018 );
   xor U17348 ( n18018,n18007,n16931 );
   nor U17349 ( n18016,n17825,n18019 );
   xor U17350 ( n18019,n18001,n15467 );
   nor U17351 ( n18012,n18020,n18002 );
   nor U17352 ( n18020,n17819,n18021,n18022 );
   nor U17353 ( n18022,n18023,n17823 );
   xor U17354 ( n18023,p3_reg2_reg_11_,n18007 );
   nand U17355 ( n18007,n18024,n18025 );
   nand U17356 ( n18025,p3_reg2_reg_10_,n18026 );
   or U17357 ( n18026,n18027,n18028 );
   nand U17358 ( n18024,n18028,n18027 );
   nor U17359 ( n18021,n18029,n17825 );
   xor U17360 ( n18029,p3_reg1_reg_11_,n18001 );
   nand U17361 ( n18001,n18030,n18031 );
   nand U17362 ( n18031,p3_reg1_reg_10_,n18032 );
   or U17363 ( n18032,n18033,n18028 );
   nand U17364 ( n18030,n18028,n18033 );
   nand U17365 ( n18009,n17719,n18034 );
   nand U17366 ( n18034,n18035,n18036 );
   nand U17367 ( n18036,n18037,n17989,n17993 );
   and U17368 ( n17993,n18038,n18039 );
   or U17369 ( n18039,n18040,n18014 );
   nand U17370 ( n17989,n18014,n18040 );
   nand U17371 ( n18037,n17988,n18041 );
   nand U17372 ( n18035,n18042,n17988,n18043 );
   xor U17373 ( n18043,n18002,n18040 );
   nand U17374 ( n18040,n18044,n18045 );
   nand U17375 ( n18045,n17731,n16931 );
   not U17376 ( n16931,p3_reg2_reg_11_ );
   nand U17377 ( n18044,n15937,n15467 );
   not U17378 ( n15467,p3_reg1_reg_11_ );
   nand U17379 ( n18042,n18046,n18038 );
   nand U17380 ( n18038,n18047,n18028 );
   nand U17381 ( n18008,n17777,p3_addr_reg_11_ );
   nand U17382 ( p3_u3192,n18048,n18049,n18050,n18051 );
   nor U17383 ( n18051,n18052,n18053 );
   and U17384 ( n18053,p3_addr_reg_10_,n17777 );
   nor U17385 ( n18052,n17988,n18046,n17763 );
   nand U17386 ( n17988,n18054,n18055 );
   nand U17387 ( n18050,p3_reg3_reg_10_,p3_u3151 );
   nand U17388 ( n18049,n18028,n18056 );
   nand U17389 ( n18056,n18057,n18058,n18059 );
   nand U17390 ( n18059,n18060,n17708 );
   xor U17391 ( n18060,p3_reg2_reg_10_,n18027 );
   nand U17392 ( n18058,n18061,n17719 );
   xor U17393 ( n18061,n18055,n18041 );
   nand U17394 ( n18057,n18062,n17734 );
   xor U17395 ( n18062,p3_reg1_reg_10_,n18033 );
   nand U17396 ( n18048,n18054,n18063 );
   nand U17397 ( n18063,n17705,n18064,n18065,n18066 );
   nand U17398 ( n18066,n18047,n17719,n18046 );
   not U17399 ( n18046,n18041 );
   nand U17400 ( n18041,n18067,n17991 );
   nand U17401 ( n17991,n18068,n18069 );
   nand U17402 ( n18068,n18070,n18071 );
   nand U17403 ( n18067,n17996,n17995 );
   not U17404 ( n18047,n18055 );
   nand U17405 ( n18055,n18072,n18073 );
   nand U17406 ( n18073,n17731,n18074 );
   nand U17407 ( n18072,n15937,n18075 );
   nand U17408 ( n18065,n17734,n18076 );
   xor U17409 ( n18076,n18033,n18075 );
   not U17410 ( n18075,p3_reg1_reg_10_ );
   nand U17411 ( n18033,n18077,n18078 );
   nand U17412 ( n18078,p3_reg1_reg_9_,n18079 );
   or U17413 ( n18079,n18080,n17995 );
   nand U17414 ( n18077,n18080,n17995 );
   nand U17415 ( n18064,n17708,n18081 );
   xor U17416 ( n18081,n18027,n18074 );
   not U17417 ( n18074,p3_reg2_reg_10_ );
   nand U17418 ( n18027,n18082,n18083 );
   nand U17419 ( n18083,p3_reg2_reg_9_,n18084 );
   or U17420 ( n18084,n18085,n17995 );
   nand U17421 ( n18082,n18085,n17995 );
   nand U17422 ( p3_u3191,n18086,n18087,n18088,n18089 );
   nand U17423 ( n18089,n18070,n18090 );
   nand U17424 ( n18090,n17705,n18091,n18092,n18093 );
   nand U17425 ( n18093,n17719,n18094 );
   xor U17426 ( n18094,n17996,n18069 );
   not U17427 ( n17996,n18071 );
   nand U17428 ( n18092,n17734,n18095 );
   xor U17429 ( n18095,n18080,n18096 );
   nand U17430 ( n18091,n17708,n18097 );
   xor U17431 ( n18097,n18085,n18098 );
   nand U17432 ( n18088,n18099,n17995 );
   nand U17433 ( n18099,n18100,n18101,n18102 );
   nand U17434 ( n18102,n18103,n17708 );
   xor U17435 ( n18103,p3_reg2_reg_9_,n18085 );
   nand U17436 ( n18085,n18104,n18105 );
   nand U17437 ( n18105,p3_reg2_reg_8_,n18106 );
   or U17438 ( n18106,n18107,n18108 );
   nand U17439 ( n18104,n18108,n18107 );
   nand U17440 ( n18101,n18109,n17719 );
   xor U17441 ( n18109,n18071,n18069 );
   nand U17442 ( n18069,n18110,n18111 );
   nand U17443 ( n18111,n18108,n18112 );
   nand U17444 ( n18112,n18113,n18114 );
   nand U17445 ( n18110,n18115,n18116 );
   nand U17446 ( n18071,n18117,n18118 );
   nand U17447 ( n18118,n17731,n18098 );
   not U17448 ( n18098,p3_reg2_reg_9_ );
   nand U17449 ( n18117,n15937,n18096 );
   not U17450 ( n18096,p3_reg1_reg_9_ );
   nand U17451 ( n18100,n18119,n17734 );
   xor U17452 ( n18119,p3_reg1_reg_9_,n18080 );
   nand U17453 ( n18080,n18120,n18121 );
   nand U17454 ( n18121,p3_reg1_reg_8_,n18122 );
   or U17455 ( n18122,n18123,n18108 );
   nand U17456 ( n18120,n18108,n18123 );
   nand U17457 ( n18087,n17777,p3_addr_reg_9_ );
   nand U17458 ( n18086,p3_reg3_reg_9_,p3_u3151 );
   nand U17459 ( p3_u3190,n18124,n18125,n18126,n18127 );
   nor U17460 ( n18127,n18128,n18129 );
   and U17461 ( n18129,p3_addr_reg_8_,n17777 );
   nor U17462 ( n18128,n17763,n18113,n18130 );
   xor U17463 ( n18130,n18115,n18108 );
   nand U17464 ( n18126,p3_reg3_reg_8_,p3_u3151 );
   nand U17465 ( n18125,n18108,n18131 );
   nand U17466 ( n18131,n18132,n18133,n18134 );
   nand U17467 ( n18134,n18135,n17708 );
   xor U17468 ( n18135,p3_reg2_reg_8_,n18107 );
   nand U17469 ( n18133,n18113,n18114,n17719 );
   nand U17470 ( n18132,n18136,n17734 );
   xor U17471 ( n18136,p3_reg1_reg_8_,n18123 );
   nand U17472 ( n18124,n18137,n18138 );
   nand U17473 ( n18138,n17705,n18139,n18140,n18141 );
   nand U17474 ( n18141,n18115,n18113,n17719 );
   not U17475 ( n18113,n18116 );
   nand U17476 ( n18116,n18142,n18143 );
   nand U17477 ( n18143,n18144,n18145 );
   nand U17478 ( n18145,n18146,n18147 );
   not U17479 ( n18144,n18148 );
   not U17480 ( n18115,n18114 );
   nand U17481 ( n18114,n18149,n18150 );
   nand U17482 ( n18150,n17731,n18151 );
   nand U17483 ( n18149,n15937,n18152 );
   nand U17484 ( n18140,n17734,n18153 );
   xor U17485 ( n18153,n18123,n18152 );
   not U17486 ( n18152,p3_reg1_reg_8_ );
   nand U17487 ( n18123,n18154,n18155 );
   nand U17488 ( n18155,p3_reg1_reg_7_,n18156 );
   or U17489 ( n18156,n18157,n18158 );
   nand U17490 ( n18154,n18157,n18158 );
   nand U17491 ( n18139,n17708,n18159 );
   xor U17492 ( n18159,n18107,n18151 );
   not U17493 ( n18151,p3_reg2_reg_8_ );
   nand U17494 ( n18107,n18160,n18161 );
   nand U17495 ( n18161,p3_reg2_reg_7_,n18162 );
   or U17496 ( n18162,n18163,n18158 );
   nand U17497 ( n18160,n18163,n18158 );
   nand U17498 ( p3_u3189,n18164,n18165,n18166,n18167 );
   nor U17499 ( n18167,n18168,n18169 );
   and U17500 ( n18169,p3_addr_reg_7_,n17777 );
   nor U17501 ( n18168,n18142,n18148,n17763 );
   or U17502 ( n18142,n18147,n18146 );
   nand U17503 ( n18166,p3_reg3_reg_7_,p3_u3151 );
   nand U17504 ( n18165,n18146,n18170 );
   nand U17505 ( n18170,n17705,n18171,n18172,n18173 );
   nand U17506 ( n18173,n18174,n17719 );
   xor U17507 ( n18174,n18147,n18148 );
   nand U17508 ( n18172,n17734,n18175 );
   xor U17509 ( n18175,n18157,n15499 );
   nand U17510 ( n18171,n17708,n18176 );
   xor U17511 ( n18176,n18163,n18177 );
   nand U17512 ( n18164,n18178,n18158 );
   nand U17513 ( n18178,n18179,n18180,n18181 );
   nand U17514 ( n18181,n18182,n17708 );
   xor U17515 ( n18182,p3_reg2_reg_7_,n18163 );
   nand U17516 ( n18163,n18183,n18184 );
   nand U17517 ( n18184,p3_reg2_reg_6_,n18185 );
   or U17518 ( n18185,n18186,n18187 );
   nand U17519 ( n18183,n18187,n18186 );
   nand U17520 ( n18180,n18147,n18148,n17719 );
   nand U17521 ( n18148,n18188,n18189 );
   nand U17522 ( n18188,n18190,n18191 );
   nand U17523 ( n18147,n18192,n18193 );
   nand U17524 ( n18193,n17731,n18177 );
   not U17525 ( n18177,p3_reg2_reg_7_ );
   nand U17526 ( n18192,n15937,n15499 );
   not U17527 ( n15499,p3_reg1_reg_7_ );
   nand U17528 ( n18179,n18194,n17734 );
   xor U17529 ( n18194,p3_reg1_reg_7_,n18157 );
   nand U17530 ( n18157,n18195,n18196 );
   nand U17531 ( n18196,p3_reg1_reg_6_,n18197 );
   or U17532 ( n18197,n18198,n18187 );
   nand U17533 ( n18195,n18187,n18198 );
   nand U17534 ( p3_u3188,n18199,n18200,n18201 );
   nor U17535 ( n18201,n18202,n18203,n18204 );
   nor U17536 ( n18204,n18205,n18187 );
   nor U17537 ( n18205,n17819,n18206,n18207 );
   nor U17538 ( n18207,n18208,n17823 );
   xor U17539 ( n18208,p3_reg2_reg_6_,n18186 );
   nor U17540 ( n18206,n18209,n17825 );
   xor U17541 ( n18209,p3_reg1_reg_6_,n18198 );
   nor U17542 ( n18203,n18210,n18211 );
   nor U17543 ( n18210,n18212,n18213 );
   nor U17544 ( n18213,n17823,n18214 );
   xor U17545 ( n18214,n18186,n18215 );
   nand U17546 ( n18186,n18216,n18217 );
   nand U17547 ( n18217,p3_reg2_reg_5_,n18218 );
   or U17548 ( n18218,n18219,n18220 );
   nand U17549 ( n18216,n18219,n18220 );
   nor U17550 ( n18212,n17825,n18221 );
   xor U17551 ( n18221,n18198,n18222 );
   nand U17552 ( n18198,n18223,n18224 );
   nand U17553 ( n18224,p3_reg1_reg_5_,n18225 );
   or U17554 ( n18225,n18226,n18220 );
   nand U17555 ( n18223,n18226,n18220 );
   nand U17556 ( n18200,n17719,n18227 );
   nand U17557 ( n18227,n18228,n18229 );
   nand U17558 ( n18229,n18191,n18189,n18190 );
   and U17559 ( n18190,n18230,n18231 );
   or U17560 ( n18231,n18232,n18211 );
   nand U17561 ( n18189,n18211,n18232 );
   nand U17562 ( n18191,n18233,n18234 );
   nand U17563 ( n18228,n18235,n18233,n18236 );
   xor U17564 ( n18236,n18187,n18232 );
   nand U17565 ( n18232,n18237,n18238 );
   nand U17566 ( n18238,n17731,n18215 );
   not U17567 ( n18215,p3_reg2_reg_6_ );
   nand U17568 ( n18237,n15937,n18222 );
   not U17569 ( n18222,p3_reg1_reg_6_ );
   nand U17570 ( n18235,n18239,n18230 );
   nand U17571 ( n18230,n18240,n18220 );
   nand U17572 ( n18199,n17777,p3_addr_reg_6_ );
   nand U17573 ( p3_u3187,n18241,n18242,n18243,n18244 );
   nor U17574 ( n18244,n18245,n18246 );
   and U17575 ( n18246,p3_addr_reg_5_,n17777 );
   nor U17576 ( n18245,n18233,n18239,n17763 );
   nand U17577 ( n18233,n18247,n18248 );
   nand U17578 ( n18243,p3_reg3_reg_5_,p3_u3151 );
   nand U17579 ( n18242,n18249,n18220 );
   nand U17580 ( n18249,n18250,n18251,n18252 );
   nand U17581 ( n18252,n18253,n17708 );
   xor U17582 ( n18253,p3_reg2_reg_5_,n18219 );
   nand U17583 ( n18251,n18254,n17719 );
   xor U17584 ( n18254,n18248,n18234 );
   nand U17585 ( n18250,n18255,n17734 );
   xor U17586 ( n18255,p3_reg1_reg_5_,n18226 );
   nand U17587 ( n18241,n18247,n18256 );
   nand U17588 ( n18256,n17705,n18257,n18258,n18259 );
   nand U17589 ( n18259,n18240,n17719,n18239 );
   not U17590 ( n18239,n18234 );
   nand U17591 ( n18234,n18260,n18261 );
   nand U17592 ( n18261,n18262,n18263 );
   nand U17593 ( n18262,n18264,n18265 );
   nand U17594 ( n18260,n18266,n18267 );
   not U17595 ( n18240,n18248 );
   nand U17596 ( n18248,n18268,n18269 );
   nand U17597 ( n18269,n17731,n18270 );
   nand U17598 ( n18268,n15937,n18271 );
   nand U17599 ( n18258,n17734,n18272 );
   xor U17600 ( n18272,n18226,n18271 );
   not U17601 ( n18271,p3_reg1_reg_5_ );
   nand U17602 ( n18226,n18273,n18274 );
   nand U17603 ( n18274,p3_reg1_reg_4_,n18275 );
   or U17604 ( n18275,n18276,n18267 );
   nand U17605 ( n18273,n18267,n18276 );
   nand U17606 ( n18257,n17708,n18277 );
   xor U17607 ( n18277,n18219,n18270 );
   not U17608 ( n18270,p3_reg2_reg_5_ );
   nand U17609 ( n18219,n18278,n18279 );
   nand U17610 ( n18279,p3_reg2_reg_4_,n18280 );
   or U17611 ( n18280,n18281,n18267 );
   nand U17612 ( n18278,n18267,n18281 );
   nand U17613 ( p3_u3186,n18282,n18283,n18284,n18285 );
   nand U17614 ( n18285,n18267,n18286 );
   nand U17615 ( n18286,n18287,n18288,n18289 );
   nand U17616 ( n18289,n18290,n17708 );
   xor U17617 ( n18290,p3_reg2_reg_4_,n18281 );
   nand U17618 ( n18288,n18291,n17719 );
   xor U17619 ( n18291,n18265,n18263 );
   nand U17620 ( n18287,n18292,n17734 );
   xor U17621 ( n18292,p3_reg1_reg_4_,n18276 );
   nand U17622 ( n18284,n18264,n18293 );
   nand U17623 ( n18293,n17705,n18294,n18295,n18296 );
   nand U17624 ( n18296,n17719,n18297 );
   xor U17625 ( n18297,n18266,n18263 );
   nand U17626 ( n18263,n18298,n18299 );
   nand U17627 ( n18299,n18300,n18301 );
   nand U17628 ( n18300,n18302,n18303 );
   nand U17629 ( n18298,n18304,n18305 );
   not U17630 ( n18266,n18265 );
   nand U17631 ( n18265,n18306,n18307 );
   nand U17632 ( n18307,n17731,n18308 );
   nand U17633 ( n18306,n15937,n18309 );
   nand U17634 ( n18295,n17734,n18310 );
   xor U17635 ( n18310,n18276,n18309 );
   not U17636 ( n18309,p3_reg1_reg_4_ );
   nand U17637 ( n18276,n18311,n18312 );
   nand U17638 ( n18312,p3_reg1_reg_3_,n18313 );
   or U17639 ( n18313,n18314,n18301 );
   nand U17640 ( n18311,n18314,n18301 );
   nand U17641 ( n18294,n17708,n18315 );
   xor U17642 ( n18315,n18281,n18308 );
   not U17643 ( n18308,p3_reg2_reg_4_ );
   nand U17644 ( n18281,n18316,n18317 );
   nand U17645 ( n18317,p3_reg2_reg_3_,n18318 );
   or U17646 ( n18318,n18319,n18301 );
   nand U17647 ( n18316,n18319,n18301 );
   nand U17648 ( n18283,n17777,p3_addr_reg_4_ );
   nand U17649 ( n18282,p3_reg3_reg_4_,p3_u3151 );
   nand U17650 ( p3_u3185,n18320,n18321,n18322 );
   nor U17651 ( n18322,n18323,n18324,n18325 );
   nor U17652 ( n18325,n18326,n18327 );
   nor U17653 ( n18327,n18328,n18329,n18330 );
   nor U17654 ( n18330,n17825,n18331 );
   xor U17655 ( n18331,n18314,n15531 );
   nor U17656 ( n18329,n17763,n18304,n18305 );
   nor U17657 ( n18328,n17823,n18332 );
   xor U17658 ( n18332,n18319,n16706 );
   nor U17659 ( n18324,n18333,n18301 );
   nor U17660 ( n18333,n18334,n18335,n18336,n17819 );
   nor U17661 ( n18336,n18337,n17823 );
   xor U17662 ( n18337,p3_reg2_reg_3_,n18319 );
   nand U17663 ( n18319,n18338,n18339 );
   nand U17664 ( n18339,p3_reg2_reg_2_,n18340 );
   or U17665 ( n18340,n18341,n18342 );
   nand U17666 ( n18338,n18342,n18341 );
   nor U17667 ( n18335,n18343,n17825 );
   xor U17668 ( n18343,p3_reg1_reg_3_,n18314 );
   nand U17669 ( n18314,n18344,n18345 );
   nand U17670 ( n18345,p3_reg1_reg_2_,n18346 );
   or U17671 ( n18346,n18347,n18342 );
   nand U17672 ( n18344,n18342,n18347 );
   nor U17673 ( n18334,n17763,n18305,n18303 );
   nand U17674 ( n18321,n17719,n18305,n18348 );
   xor U17675 ( n18348,n18326,n18304 );
   not U17676 ( n18304,n18303 );
   nand U17677 ( n18303,n18349,n18350 );
   nand U17678 ( n18350,n17731,n16706 );
   not U17679 ( n16706,p3_reg2_reg_3_ );
   nand U17680 ( n18349,n15937,n15531 );
   not U17681 ( n15531,p3_reg1_reg_3_ );
   not U17682 ( n18305,n18302 );
   nor U17683 ( n18302,n18351,n18352 );
   and U17684 ( n18352,n18353,n18354 );
   nand U17685 ( n18354,n18355,n18356 );
   nand U17686 ( n18320,n17777,p3_addr_reg_3_ );
   nand U17687 ( p3_u3184,n18357,n18358,n18359,n18360 );
   nand U17688 ( n18360,n17719,n18353,n18351 );
   nor U17689 ( n18351,n18356,n18355 );
   nand U17690 ( n18359,n17777,p3_addr_reg_2_ );
   nand U17691 ( n18358,p3_reg3_reg_2_,p3_u3151 );
   nor U17692 ( n18357,n18361,n18362 );
   nor U17693 ( n18362,n18363,n18342 );
   nor U17694 ( n18363,n18364,n18365,n18366,n17819 );
   nor U17695 ( n18366,n18367,n17823 );
   xor U17696 ( n18367,p3_reg2_reg_2_,n18341 );
   nor U17697 ( n18365,n18368,n17825 );
   xor U17698 ( n18368,p3_reg1_reg_2_,n18347 );
   nor U17699 ( n18364,n17763,n18369 );
   xor U17700 ( n18369,n18356,n18353 );
   nor U17701 ( n18361,n18370,n18355 );
   nor U17702 ( n18370,n18371,n18372,n18373 );
   nor U17703 ( n18373,n17825,n18374 );
   xor U17704 ( n18374,n18347,n15542 );
   nand U17705 ( n18347,n18375,n18376 );
   nand U17706 ( n18376,p3_reg1_reg_1_,n18377 );
   nand U17707 ( n18377,n18378,n18379 );
   nand U17708 ( n18375,n18380,n18381 );
   nor U17709 ( n18372,n17763,n18353,n18382 );
   not U17710 ( n18382,n18356 );
   nand U17711 ( n18356,n18383,n18384 );
   nand U17712 ( n18384,n17731,n18385 );
   nand U17713 ( n18383,n15937,n15542 );
   not U17714 ( n15542,p3_reg1_reg_2_ );
   and U17715 ( n18353,n18386,n18387 );
   nand U17716 ( n18387,n18378,n18388 );
   nand U17717 ( n18388,n18389,n18390 );
   or U17718 ( n18386,n18390,n18389 );
   nor U17719 ( n18371,n17823,n18391 );
   xor U17720 ( n18391,n18341,n18385 );
   not U17721 ( n18385,p3_reg2_reg_2_ );
   nand U17722 ( n18341,n18392,n18393 );
   nand U17723 ( n18393,p3_reg2_reg_1_,n18394 );
   nand U17724 ( n18394,n18378,n18395 );
   nand U17725 ( n18392,n18396,n18381 );
   nand U17726 ( p3_u3183,n18397,n18398,n18399,n18400 );
   nand U17727 ( n18400,n18378,n18401 );
   nand U17728 ( n18401,n17705,n18402,n18403 );
   nor U17729 ( n18403,n18404,n18405,n18406,n18407 );
   nor U17730 ( n18407,n15551,n18408 );
   nor U17731 ( n18406,p3_reg1_reg_1_,n18380,n17825 );
   nor U17732 ( n18405,n16638,n18409 );
   nor U17733 ( n18404,p3_reg2_reg_1_,n18396,n17823 );
   nand U17734 ( n18402,n17719,n18410 );
   nand U17735 ( n18399,n18411,n18381 );
   nand U17736 ( n18411,n18412,n18413,n18414 );
   nor U17737 ( n18414,n18415,n18416,n18417 );
   nor U17738 ( n18417,n15551,n18380,n17825 );
   nor U17739 ( n18416,p3_reg1_reg_1_,n18408 );
   nor U17740 ( n18415,n17763,n18410 );
   xor U17741 ( n18410,n18389,n18390 );
   and U17742 ( n18389,n18418,n18419 );
   nand U17743 ( n18419,n17731,n16638 );
   not U17744 ( n16638,p3_reg2_reg_1_ );
   nand U17745 ( n18418,n15937,n15551 );
   not U17746 ( n15551,p3_reg1_reg_1_ );
   or U17747 ( n18413,n18409,p3_reg2_reg_1_ );
   nand U17748 ( n18412,n17708,n18395,p3_reg2_reg_1_ );
   nand U17749 ( n18398,n17777,p3_addr_reg_1_ );
   not U17750 ( n17777,n17704 );
   nand U17751 ( n18397,p3_reg3_reg_1_,p3_u3151 );
   nand U17752 ( p3_u3182,n18408,n18409,n18420,n18421 );
   nor U17753 ( n18421,n18422,n18423,n18424 );
   nor U17754 ( n18424,n15076,n17704 );
   not U17755 ( n15076,p3_addr_reg_0_ );
   nor U17756 ( n18423,n18425,n16326 );
   nor U17757 ( n18425,n17819,n18426,n18427 );
   nor U17758 ( n18427,p3_reg2_reg_0_,n17823 );
   nor U17759 ( n18426,p3_reg1_reg_0_,n17825 );
   not U17760 ( n17819,n17705 );
   nand U17761 ( n17705,n18428,n18429 );
   nand U17762 ( n18429,n15939,n15191 );
   or U17763 ( n18428,n18430,n15939 );
   not U17764 ( n15939,n18431 );
   nor U17765 ( n18422,p3_state_reg,n16600 );
   not U17766 ( n16600,p3_reg3_reg_0_ );
   nand U17767 ( n18420,n17719,n18432 );
   nand U17768 ( n18432,n18433,n18434,n18390 );
   nand U17769 ( n18390,n18435,n18436,p3_ir_reg_0_ );
   nand U17770 ( n18436,p3_reg1_reg_0_,n15937 );
   nand U17771 ( n18435,n17731,p3_reg2_reg_0_ );
   nand U17772 ( n18434,n18380,n15937 );
   nand U17773 ( n18433,n18396,n17731 );
   nand U17774 ( n18409,n17708,n18396 );
   not U17775 ( n18396,n18395 );
   nand U17776 ( n18395,p3_reg2_reg_0_,n16326 );
   nand U17777 ( n18408,n17734,n18380 );
   not U17778 ( n18380,n18379 );
   nand U17779 ( n18379,p3_reg1_reg_0_,n16326 );
   nand U17780 ( n18430,n18438,n18439 );
   nand U17781 ( n18439,n17704,p3_state_reg,n15944 );
   nand U17782 ( n18438,n18440,n17704,n15567 );
   nand U17783 ( n17704,n18441,n18442,n18443 );
   nand U17784 ( n18442,n17657,n16262 );
   nand U17785 ( n18441,n18437,n15824 );
   nand U17786 ( n18440,n16890,n17662,n18444 );
   nor U17787 ( n18444,n17685,n17479,n16260 );
   nor U17788 ( n16890,n17027,n17029 );
   nand U17789 ( n17029,n16628,n16631 );
   nand U17790 ( n17027,n15828,n15831 );
   nand U17791 ( p3_u3181,n18445,n18446,n18447,n18448 );
   nor U17792 ( n18448,n18449,n18450,n18451 );
   nor U17793 ( n18451,n17051,n18452 );
   nor U17794 ( n18450,n17555,n18453 );
   and U17795 ( n18449,p3_u3151,p3_reg3_reg_15_ );
   nand U17796 ( n18447,n18454,n15243 );
   nand U17797 ( n18446,n18455,n18456 );
   xor U17798 ( n18455,n18457,n18458 );
   xor U17799 ( n18458,n18459,n15240 );
   not U17800 ( n18457,n18460 );
   nand U17801 ( n18445,n17052,n18461 );
   nand U17802 ( p3_u3180,n18462,n18463,n18464,n18465 );
   nor U17803 ( n18465,n18466,n18467,n18468 );
   nor U17804 ( n18468,n18469,n18470 );
   nor U17805 ( n18467,n17402,n18453 );
   not U17806 ( n17402,n15329 );
   and U17807 ( n18466,p3_u3151,p3_reg3_reg_26_ );
   nand U17808 ( n18464,n18471,n15204 );
   nand U17809 ( n18463,n18472,n18473,n18456 );
   nand U17810 ( n18473,n18474,n18475 );
   nand U17811 ( n18474,n18476,n18477 );
   nand U17812 ( n18472,n18476,n18477,n18478 );
   not U17813 ( n18478,n18475 );
   nand U17814 ( n18475,n18479,n18480 );
   or U17815 ( n18477,n18481,n18482 );
   nand U17816 ( n18462,n17373,n18483 );
   nand U17817 ( p3_u3179,n18484,n18485,n18486,n18487 );
   nor U17818 ( n18487,n18202,n18488,n18489 );
   nor U17819 ( n18489,n16718,n18470 );
   nor U17820 ( n18488,n15507,n18452 );
   nor U17821 ( n18202,p3_state_reg,n18490 );
   not U17822 ( n18490,p3_reg3_reg_6_ );
   nand U17823 ( n18486,n16769,n18461 );
   nand U17824 ( n18485,n18491,n18492,n18456 );
   nand U17825 ( n18492,n18493,n18494 );
   xor U17826 ( n18493,n18495,n15267 );
   nand U17827 ( n18491,n18496,n18497,n18498 );
   nand U17828 ( n18484,n18499,n15509 );
   nand U17829 ( p3_u3178,n18500,n18501,n18502,n18503 );
   nor U17830 ( n18503,n18504,n18505,n18506 );
   nor U17831 ( n18506,n15397,n18452 );
   nor U17832 ( n18505,n17129,n18470 );
   nor U17833 ( n18504,p3_state_reg,n18507 );
   nand U17834 ( n18502,n18499,n15401 );
   nand U17835 ( n18501,n18508,n18456 );
   xor U17836 ( n18508,n18509,n18510 );
   xor U17837 ( n18510,n18511,n15409 );
   not U17838 ( n15409,n15231 );
   nand U17839 ( n18500,n17137,n18461 );
   nand U17840 ( p3_u3177,n18512,n18513,n18514,n18515 );
   nor U17841 ( n18515,n18516,n18517 );
   nor U17842 ( n18517,n15796,n18470 );
   nor U17843 ( n18516,n15783,n18452 );
   nand U17844 ( n18514,n18499,n15538 );
   nand U17845 ( n18513,n18456,n18518 );
   nand U17846 ( n18518,n18519,n18520,n18521 );
   nand U17847 ( n18521,n18522,n18523 );
   or U17848 ( n18520,n18523,n16691,n18524 );
   nand U17849 ( n18519,n18525,n18524 );
   xor U17850 ( n18525,n16691,n18523 );
   nand U17851 ( n18512,p3_reg3_reg_2_,n18526 );
   nand U17852 ( p3_u3176,n18527,n18528,n18529,n18530 );
   nor U17853 ( n18530,n18011,n18531,n18532 );
   nor U17854 ( n18532,n16985,n18452 );
   nor U17855 ( n18531,n16932,n18453 );
   nor U17856 ( n18011,p3_state_reg,n18533 );
   nand U17857 ( n18529,n16933,n18461 );
   nand U17858 ( n18528,n18534,n18535,n18456 );
   nand U17859 ( n18535,n18536,n18537 );
   nand U17860 ( n18536,n18538,n18539 );
   nand U17861 ( n18534,n18540,n18541 );
   xor U17862 ( n18540,n16883,n18542 );
   nand U17863 ( n18527,n18454,n15255 );
   nand U17864 ( p3_u3175,n18543,n18544,n18545,n18546 );
   nor U17865 ( n18546,n18547,n18548,n18549 );
   nor U17866 ( n18549,n17537,n18470 );
   nor U17867 ( n18548,n17584,n18453 );
   not U17868 ( n17584,n15366 );
   nor U17869 ( n18547,p3_state_reg,n18550 );
   nand U17870 ( n18545,n18471,n15216 );
   nand U17871 ( n18544,n18551,n18456 );
   xor U17872 ( n18551,n18552,n18553 );
   xor U17873 ( n18553,n18554,n15219 );
   nand U17874 ( n18543,n17264,n18483 );
   nand U17875 ( p3_u3174,n18555,n18556,n18557,n18558 );
   nor U17876 ( n18558,n18559,n18560,n18561 );
   nor U17877 ( n18561,n18562,n18452 );
   nor U17878 ( n18560,n16985,n18470 );
   and U17879 ( n18559,p3_u3151,p3_reg3_reg_13_ );
   nand U17880 ( n18557,n18499,n15444 );
   nand U17881 ( n18556,n18563,n18564,n18456 );
   nand U17882 ( n18564,n18565,n18566,n18567 );
   nand U17883 ( n18567,n18568,n18569 );
   nand U17884 ( n18565,n18570,n18571 );
   nand U17885 ( n18563,n18572,n18568,n18573 );
   nand U17886 ( n18572,n18574,n18566 );
   nand U17887 ( n18555,n17008,n18461 );
   nand U17888 ( p3_u3173,n18575,n18576,n18577,n18578 );
   nor U17889 ( n18578,n18579,n18580,n18581 );
   nor U17890 ( n18581,n17537,n18452 );
   nor U17891 ( n18580,n15397,n18470 );
   nor U17892 ( n18579,p3_state_reg,n18582 );
   nand U17893 ( n18577,n18499,n15661 );
   nand U17894 ( n18576,n18456,n18583 );
   xor U17895 ( n18583,n18584,n18585 );
   xor U17896 ( n18584,n15225,n18586 );
   nand U17897 ( n18575,n17218,n18483 );
   nand U17898 ( p3_u3172,n18587,n18588,n18589,n18590 );
   nand U17899 ( n18590,p3_reg3_reg_0_,n18526 );
   nand U17900 ( n18589,n18456,n15557 );
   nand U17901 ( n15557,n16643,n18591 );
   nand U17902 ( n18591,n16170,n15285 );
   nand U17903 ( n16643,n16611,n15561 );
   nand U17904 ( n18588,n18499,n15561 );
   nand U17905 ( n18587,n18471,n15282 );
   nand U17906 ( p3_u3171,n18592,n18593,n18594,n18595 );
   nor U17907 ( n18595,n18596,n18597,n18598 );
   nor U17908 ( n18598,n15908,n18470 );
   nor U17909 ( n18597,n16860,n18452 );
   and U17910 ( n18596,p3_u3151,p3_reg3_reg_9_ );
   nand U17911 ( n18594,n18499,n15480 );
   nand U17912 ( n18593,n18456,n18599 );
   xor U17913 ( n18599,n18600,n18601 );
   xor U17914 ( n18600,n15258,n18602 );
   nand U17915 ( n18592,n16861,n18461 );
   nand U17916 ( p3_u3170,n18603,n18604,n18605,n18606 );
   nor U17917 ( n18606,n18607,n18608,n18609 );
   nor U17918 ( n18609,n15783,n18470 );
   nor U17919 ( n18608,n16718,n18452 );
   and U17920 ( n18607,p3_u3151,p3_reg3_reg_4_ );
   nand U17921 ( n18605,n16719,n18461 );
   nand U17922 ( n18604,n18610,n18456 );
   xor U17923 ( n18610,n18611,n18612 );
   xor U17924 ( n18611,n18613,n15273 );
   nand U17925 ( n18603,n18499,n15522 );
   nand U17926 ( p3_u3169,n18614,n18615,n18616,n18617 );
   nor U17927 ( n18617,n18618,n18619,n18620 );
   nor U17928 ( n18620,n18469,n18452 );
   nor U17929 ( n18619,n15350,n18453 );
   nor U17930 ( n18618,p3_state_reg,n18621 );
   nand U17931 ( n18616,n18454,n15216 );
   nand U17932 ( n18615,n18456,n18622 );
   xor U17933 ( n18622,n18623,n18624 );
   nand U17934 ( n18623,n18625,n18626 );
   nand U17935 ( n18614,n17335,n18483 );
   nand U17936 ( p3_u3168,n18627,n18628,n18629,n18630 );
   nor U17937 ( n18630,n18631,n18632,n18633 );
   nor U17938 ( n18632,n18634,n17110 );
   and U17939 ( n18631,p3_u3151,p3_reg3_reg_17_ );
   nand U17940 ( n18629,n18454,n15237 );
   nand U17941 ( n18628,n18635,n18636,n18456 );
   nand U17942 ( n18636,n18637,n18638 );
   nand U17943 ( n18638,n18639,n18640 );
   nand U17944 ( n18635,n18639,n18640,n18641 );
   nand U17945 ( n18627,n18471,n15231 );
   nand U17946 ( p3_u3167,n18642,n18643,n18644,n18645 );
   nor U17947 ( n18645,n18646,n18647,n18648 );
   nor U17948 ( n18648,n17571,n18470 );
   nor U17949 ( n18647,n16741,n18452 );
   and U17950 ( n18646,p3_u3151,p3_reg3_reg_5_ );
   nand U17951 ( n18644,n16742,n18461 );
   nand U17952 ( n18643,n18456,n18649 );
   nand U17953 ( n18649,n18650,n18651,n18652 );
   nand U17954 ( n18652,n18653,n18654 );
   nand U17955 ( n18651,n18655,n18656,n16718 );
   not U17956 ( n16718,n15270 );
   nand U17957 ( n18650,n18657,n15270 );
   xor U17958 ( n18657,n18656,n18655 );
   nand U17959 ( n18642,n18499,n15516 );
   nand U17960 ( p3_u3166,n18658,n18659,n18660,n18661 );
   nor U17961 ( n18661,n17815,n18662,n18663 );
   nor U17962 ( n18663,n17129,n18452 );
   nor U17963 ( n18662,n17091,n18453 );
   not U17964 ( n17091,n15418 );
   nor U17965 ( n17815,p3_state_reg,n18664 );
   nand U17966 ( n18660,n17092,n18461 );
   nand U17967 ( n18659,n18665,n18456 );
   xor U17968 ( n18665,n18666,n18667 );
   xor U17969 ( n18666,n18668,n17051 );
   nand U17970 ( n18658,n18454,n15240 );
   nand U17971 ( p3_u3165,n18669,n18670,n18671,n18672 );
   nor U17972 ( n18672,n18673,n18674,n18675 );
   nor U17973 ( n18675,n17427,n18452 );
   and U17974 ( n18673,p3_u3151,p3_reg3_reg_25_ );
   nand U17975 ( n18671,n18454,n15213 );
   nand U17976 ( n18670,n18676,n18456 );
   xor U17977 ( n18676,n18677,n18481 );
   nand U17978 ( n18481,n18678,n18626 );
   nand U17979 ( n18678,n18679,n18625 );
   nor U17980 ( n18677,n18482,n18680 );
   not U17981 ( n18482,n18681 );
   nand U17982 ( n18669,n17362,n18483 );
   nand U17983 ( p3_u3164,n18682,n18683,n18684,n18685 );
   nor U17984 ( n18685,n18686,n18687,n18688 );
   nor U17985 ( n18688,n16966,n18453 );
   and U17986 ( n18687,n18461,n16967 );
   nor U17987 ( n18686,p3_state_reg,n18689 );
   nand U17988 ( n18684,n18454,n15252 );
   nand U17989 ( n18683,n18690,n18691,n18456 );
   nand U17990 ( n18691,n18571,n18566,n18570 );
   nand U17991 ( n18690,n18692,n18574 );
   not U17992 ( n18574,n18570 );
   nand U17993 ( n18570,n18538,n18693 );
   nand U17994 ( n18693,n18541,n18539 );
   not U17995 ( n18541,n18537 );
   nand U17996 ( n18537,n18694,n18695 );
   xor U17997 ( n18692,n18696,n15249 );
   nand U17998 ( n18682,n18471,n15246 );
   nand U17999 ( p3_u3163,n18697,n18698,n18699,n18700 );
   nor U18000 ( n18700,n18701,n18702,n18703 );
   nor U18001 ( n18702,n17541,n18470 );
   not U18002 ( n17541,n15225 );
   and U18003 ( n18701,p3_u3151,p3_reg3_reg_21_ );
   nand U18004 ( n18699,n18471,n15219 );
   nand U18005 ( n18698,n18704,n18705,n18456 );
   nand U18006 ( n18705,n18706,n18707 );
   nand U18007 ( n18707,n18708,n18709 );
   nand U18008 ( n18704,n18708,n18709,n18710 );
   nand U18009 ( n18697,n17229,n18483 );
   nand U18010 ( p3_u3162,n18711,n18712,n18713,n18714 );
   nor U18011 ( n18714,n18715,n18716 );
   nor U18012 ( n18716,n16611,n18470 );
   not U18013 ( n16611,n15285 );
   nor U18014 ( n18715,n16691,n18452 );
   nand U18015 ( n18713,n18499,n15548 );
   nand U18016 ( n18712,n18717,n18456 );
   xor U18017 ( n18717,n18718,n18719 );
   and U18018 ( n18718,n18720,n18721 );
   nand U18019 ( n18711,p3_reg3_reg_1_,n18526 );
   nand U18020 ( n18526,n18634,p3_state_reg );
   nand U18021 ( p3_u3161,n18722,n18723,n18724,n18725 );
   nor U18022 ( n18725,n18726,n18727,n18728 );
   nor U18023 ( n18728,n15507,n18470 );
   nor U18024 ( n18727,n18634,n16830 );
   nor U18025 ( n18726,p3_state_reg,n18729 );
   nand U18026 ( n18724,n18499,n15489 );
   nand U18027 ( n18723,n18456,n18730 );
   xor U18028 ( n18730,n18731,n18732 );
   xor U18029 ( n18731,n15261,n18733 );
   nand U18030 ( n18722,n18471,n15258 );
   nand U18031 ( p3_u3160,n18734,n18735,n18736,n18737 );
   nor U18032 ( n18737,n18738,n18739,n18740 );
   nor U18033 ( n18740,n15617,n18470 );
   and U18034 ( n18739,n18483,n17471 );
   and U18035 ( n18738,p3_u3151,p3_reg3_reg_28_ );
   nand U18036 ( n18736,n18499,n15311 );
   nand U18037 ( n18735,n18741,n18742,n18456 );
   nand U18038 ( n18742,n18743,n18744 );
   nand U18039 ( n18744,n18745,n18746 );
   nand U18040 ( n18746,n18747,n18748 );
   not U18041 ( n18747,n18749 );
   nand U18042 ( n18741,n18750,n18751 );
   nand U18043 ( n18751,n18748,n18752 );
   nand U18044 ( n18752,n18749,n18745 );
   not U18045 ( n18750,n18743 );
   nand U18046 ( n18743,n18753,n18754 );
   or U18047 ( n18754,n18755,n16296 );
   nor U18048 ( n16296,n17489,n17500 );
   not U18049 ( n17500,n17493 );
   nand U18050 ( n17493,n15311,n15201 );
   not U18051 ( n17489,n17499 );
   nand U18052 ( n17499,n17519,n17470 );
   nand U18053 ( n18753,n18756,n18755 );
   nand U18054 ( n18756,n15848,n15845 );
   nand U18055 ( n15845,n17470,n15201 );
   not U18056 ( n17470,n15311 );
   nand U18057 ( n15848,n17519,n15311 );
   nand U18058 ( n15311,n18757,n18758 );
   nand U18059 ( n18758,n16555,n17640 );
   xor U18060 ( n16555,n18759,n17684 );
   nand U18061 ( n17684,n18760,n18761 );
   nand U18062 ( n18761,p2_datao_reg_27_,n18762 );
   or U18063 ( n18762,n18763,n18764 );
   nand U18064 ( n18760,n18764,n18763 );
   xor U18065 ( n18759,p2_datao_reg_28_,p1_datao_reg_28_ );
   nand U18066 ( n18757,si_28_,n17643 );
   not U18067 ( n17519,n15201 );
   nand U18068 ( n18734,n18471,n15198 );
   nand U18069 ( n15198,n18765,n18766,n18767,n17589 );
   nand U18070 ( n17589,n18768,n17661 );
   nand U18071 ( n18767,p3_reg2_reg_29_,n17590 );
   nand U18072 ( n18766,p3_reg1_reg_29_,n17591 );
   nand U18073 ( n18765,p3_reg0_reg_29_,n17592 );
   nand U18074 ( p3_u3159,n18769,n18770,n18771,n18772 );
   nor U18075 ( n18772,n17700,n18773,n18774 );
   nor U18076 ( n18774,n15874,n18453 );
   and U18077 ( n18773,n18461,n17183 );
   nor U18078 ( n17700,p3_state_reg,n18775 );
   nand U18079 ( n18771,n18471,n15225 );
   nand U18080 ( n18770,n18776,n18456 );
   xor U18081 ( n18776,n18777,n18778 );
   xor U18082 ( n18777,n15397,n18779 );
   nand U18083 ( n18769,n18454,n15231 );
   nand U18084 ( p3_u3158,n18780,n18781,n18782,n18783 );
   nor U18085 ( n18783,n18784,n18323,n18785 );
   nor U18086 ( n18785,p3_reg3_reg_3_,n18634 );
   nor U18087 ( n18323,p3_state_reg,n16708 );
   nor U18088 ( n18784,n16691,n18470 );
   not U18089 ( n16691,n15279 );
   nand U18090 ( n18782,n18471,n15273 );
   nand U18091 ( n18781,n18786,n18787,n18456 );
   nand U18092 ( n18787,n18788,n18789 );
   nand U18093 ( n18789,n18790,n18791 );
   nand U18094 ( n18786,n18792,n18793,n18790,n18791 );
   nand U18095 ( n18792,n18794,n18795 );
   not U18096 ( n18794,n18523 );
   nand U18097 ( n18780,n18499,n15528 );
   nand U18098 ( p3_u3157,n18796,n18797,n18798,n18799 );
   nor U18099 ( n18799,n18800,n18801,n18802 );
   nor U18100 ( n18802,n16883,n18452 );
   nor U18101 ( n18801,n17623,n18453 );
   nor U18102 ( n18800,p3_state_reg,n18803 );
   nand U18103 ( n18798,n16884,n18461 );
   nand U18104 ( n18797,n18456,n18804 );
   nand U18105 ( n18804,n18805,n18806 );
   nand U18106 ( n18806,n18807,n18808 );
   nand U18107 ( n18808,n18809,n18694 );
   nand U18108 ( n18805,n18810,n18694 );
   not U18109 ( n18810,n18695 );
   nand U18110 ( n18695,n18809,n18811 );
   nand U18111 ( n18796,n18454,n15258 );
   nand U18112 ( p3_u3156,n18812,n18813,n18814,n18815 );
   nor U18113 ( n18815,n18816,n18817,n18818 );
   nor U18114 ( n18818,n18819,n18452 );
   nor U18115 ( n18817,n17304,n18453 );
   and U18116 ( n18816,p3_u3151,p3_reg3_reg_23_ );
   nand U18117 ( n18814,n18454,n15219 );
   nand U18118 ( n18813,n18456,n18820 );
   xor U18119 ( n18820,n18821,n18822 );
   xor U18120 ( n18821,n17263,n18823 );
   not U18121 ( n17263,n15216 );
   nand U18122 ( n18812,n17305,n18483 );
   nand U18123 ( p3_u3155,n18824,n18825,n18826,n18827 );
   nor U18124 ( n18827,n18828,n18829,n18830 );
   nor U18125 ( n18829,n18634,n17019 );
   not U18126 ( n18634,n18461 );
   nor U18127 ( n18828,p3_state_reg,n18831 );
   nand U18128 ( n18826,n18454,n15246 );
   not U18129 ( n18454,n18470 );
   nand U18130 ( n18825,n18832,n18456 );
   xor U18131 ( n18832,n18833,n18834 );
   nor U18132 ( n18833,n18835,n18836 );
   nand U18133 ( n18824,n18471,n15240 );
   nand U18134 ( p3_u3154,n18837,n18838,n18839,n18840 );
   nor U18135 ( n18840,n18841,n18842,n18843 );
   nor U18136 ( n18843,n17427,n18470 );
   not U18137 ( n17427,n15207 );
   nor U18138 ( n18841,p3_state_reg,n18844 );
   nand U18139 ( n18839,n18471,n15201 );
   nand U18140 ( n15201,n18845,n18846,n18847,n18848 );
   nand U18141 ( n18848,n18768,n17471 );
   or U18142 ( n17471,n17661,n18849 );
   and U18143 ( n18849,p3_reg3_reg_28_,n18850 );
   nand U18144 ( n18850,n18851,n18844 );
   not U18145 ( n18844,p3_reg3_reg_27_ );
   nor U18146 ( n17661,p3_reg3_reg_27_,p3_reg3_reg_28_,n18852 );
   nand U18147 ( n18847,p3_reg2_reg_28_,n17590 );
   nand U18148 ( n18846,p3_reg1_reg_28_,n17591 );
   nand U18149 ( n18845,p3_reg0_reg_28_,n17592 );
   not U18150 ( n18471,n18452 );
   nand U18151 ( n18838,n18853,n18456 );
   xor U18152 ( n18853,n18854,n18749 );
   nand U18153 ( n18749,n18855,n18479,n18856 );
   nand U18154 ( n18856,n18476,n18679,n18625,n18480 );
   and U18155 ( n18625,n18857,n18858 );
   or U18156 ( n18858,n15859,n18859 );
   nand U18157 ( n15859,n18819,n15632 );
   or U18158 ( n18857,n17338,n18755 );
   nand U18159 ( n17338,n18819,n15350 );
   not U18160 ( n18819,n15213 );
   not U18161 ( n18679,n18624 );
   nand U18162 ( n18624,n18860,n18861 );
   nand U18163 ( n18861,n18822,n18862 );
   nand U18164 ( n18862,n18823,n15216 );
   xor U18165 ( n18822,n17304,n18755 );
   not U18166 ( n17304,n15357 );
   nand U18167 ( n15357,n18863,n18864 );
   nand U18168 ( n18864,n16511,n17640 );
   xor U18169 ( n16511,n18865,n18866 );
   xor U18170 ( n18865,p2_datao_reg_23_,p1_datao_reg_23_ );
   nand U18171 ( n18863,si_23_,n17643 );
   or U18172 ( n18860,n18823,n15216 );
   nand U18173 ( n15216,n18867,n18868,n18869,n18870 );
   nand U18174 ( n18870,n18768,n17305 );
   nand U18175 ( n17305,n18871,n18872 );
   nand U18176 ( n18872,p3_reg3_reg_23_,n18873 );
   nand U18177 ( n18873,n18874,n18550 );
   nand U18178 ( n18869,p3_reg2_reg_23_,n17590 );
   nand U18179 ( n18868,p3_reg1_reg_23_,n17591 );
   nand U18180 ( n18867,p3_reg0_reg_23_,n17592 );
   nand U18181 ( n18823,n18875,n18876 );
   nand U18182 ( n18876,n18554,n18877 );
   or U18183 ( n18877,n18552,n15219 );
   and U18184 ( n18554,n18878,n18709 );
   nand U18185 ( n18709,n18879,n17537 );
   not U18186 ( n17537,n15222 );
   xor U18187 ( n18879,n17536,n18755 );
   nand U18188 ( n18878,n18706,n18708 );
   nand U18189 ( n18708,n18880,n15222 );
   nand U18190 ( n15222,n18881,n18882,n18883,n18884 );
   nand U18191 ( n18884,n18768,n17229 );
   nand U18192 ( n17229,n18885,n18886 );
   nand U18193 ( n18886,p3_reg3_reg_21_,n18887 );
   or U18194 ( n18887,n18888,p3_reg3_reg_20_ );
   nand U18195 ( n18883,p3_reg2_reg_21_,n17590 );
   nand U18196 ( n18882,p3_reg1_reg_21_,n17591 );
   nand U18197 ( n18881,p3_reg0_reg_21_,n17592 );
   xor U18198 ( n18880,n18859,n17536 );
   not U18199 ( n17536,n15372 );
   nand U18200 ( n15372,n18889,n18890 );
   nand U18201 ( n18890,n16494,n17640 );
   xor U18202 ( n16494,n18891,n18892 );
   xor U18203 ( n18891,p2_datao_reg_21_,p1_datao_reg_21_ );
   nand U18204 ( n18889,si_21_,n17643 );
   not U18205 ( n18706,n18710 );
   nand U18206 ( n18710,n18893,n18894 );
   nand U18207 ( n18894,n18585,n18895 );
   or U18208 ( n18895,n18586,n15225 );
   xor U18209 ( n18585,n15661,n18755 );
   nand U18210 ( n15661,n18896,n18897 );
   nand U18211 ( n18897,n16485,n17640 );
   xor U18212 ( n16485,n18898,n18899 );
   xor U18213 ( n18898,p2_datao_reg_20_,p1_datao_reg_20_ );
   nand U18214 ( n18896,si_20_,n17643 );
   nand U18215 ( n18893,n15225,n18586 );
   nand U18216 ( n18586,n18900,n18901 );
   nand U18217 ( n18901,n18779,n18902 );
   nand U18218 ( n18902,n18778,n15397 );
   and U18219 ( n18779,n18903,n18904 );
   nand U18220 ( n18904,n18905,n18511 );
   nand U18221 ( n18511,n18906,n18640 );
   nand U18222 ( n18640,n18907,n17129 );
   not U18223 ( n17129,n15234 );
   xor U18224 ( n18907,n15873,n18755 );
   nand U18225 ( n18906,n18637,n18639 );
   nand U18226 ( n18639,n18908,n15234 );
   nand U18227 ( n15234,n18909,n18910,n18911,n18912 );
   nand U18228 ( n18912,n18768,n18913 );
   not U18229 ( n18913,n17110 );
   nor U18230 ( n17110,n18914,n18915 );
   and U18231 ( n18915,p3_reg3_reg_17_,n18916 );
   nand U18232 ( n18916,n18917,n18664 );
   not U18233 ( n18664,p3_reg3_reg_16_ );
   nand U18234 ( n18911,p3_reg2_reg_17_,n17590 );
   nand U18235 ( n18910,p3_reg1_reg_17_,n17591 );
   nand U18236 ( n18909,p3_reg0_reg_17_,n17592 );
   xor U18237 ( n18908,n18859,n15873 );
   not U18238 ( n15873,n15411 );
   nand U18239 ( n15411,n18918,n18919,n18920 );
   nand U18240 ( n18920,si_17_,n17643 );
   nand U18241 ( n18919,n17766,n18921 );
   not U18242 ( n17766,n17762 );
   nand U18243 ( n17762,n18922,n18923,n16469 );
   nand U18244 ( n18923,n16460,n16578 );
   nand U18245 ( n18922,p3_ir_reg_17_,n16459,p3_ir_reg_31_ );
   nand U18246 ( n18918,n16461,n17640 );
   xor U18247 ( n16461,n18924,n18925 );
   xor U18248 ( n18924,p2_datao_reg_17_,p1_datao_reg_17_ );
   not U18249 ( n18637,n18641 );
   nand U18250 ( n18641,n18926,n18927 );
   nand U18251 ( n18927,n18667,n18928 );
   nand U18252 ( n18928,n17051,n18668 );
   xor U18253 ( n18667,n15418,n18755 );
   nand U18254 ( n15418,n18929,n18930,n18931 );
   nand U18255 ( n18931,si_16_,n17643 );
   nand U18256 ( n18930,n17827,n18921 );
   not U18257 ( n17827,n17800 );
   nand U18258 ( n17800,n18932,n18933 );
   or U18259 ( n18933,p3_ir_reg_16_,p3_ir_reg_31_ );
   nand U18260 ( n18932,p3_ir_reg_31_,n16450 );
   nand U18261 ( n16450,n16459,n18934 );
   nand U18262 ( n18934,p3_ir_reg_16_,n18935 );
   not U18263 ( n16459,n16458 );
   nand U18264 ( n18929,n16451,n17640 );
   xor U18265 ( n16451,n18936,n18937 );
   xor U18266 ( n18936,p2_datao_reg_16_,p1_datao_reg_16_ );
   or U18267 ( n18926,n18668,n17051 );
   not U18268 ( n17051,n15237 );
   nand U18269 ( n15237,n18938,n18939,n18940,n18941 );
   nand U18270 ( n18941,n18768,n17092 );
   xor U18271 ( n17092,p3_reg3_reg_16_,n18917 );
   nand U18272 ( n18940,p3_reg2_reg_16_,n17590 );
   nand U18273 ( n18939,p3_reg1_reg_16_,n17591 );
   nand U18274 ( n18938,p3_reg0_reg_16_,n17592 );
   nand U18275 ( n18668,n18942,n18943 );
   nand U18276 ( n18943,n18460,n18944 );
   nand U18277 ( n18944,n18459,n15240 );
   xor U18278 ( n18460,n17555,n18755 );
   not U18279 ( n17555,n15428 );
   nand U18280 ( n15428,n18945,n18946,n18947 );
   nand U18281 ( n18947,si_15_,n17643 );
   nand U18282 ( n18946,n17861,n18921 );
   not U18283 ( n17861,n17835 );
   nand U18284 ( n17835,n18948,n18949,n18935 );
   nand U18285 ( n18949,n16443,n16578 );
   nand U18286 ( n18948,p3_ir_reg_15_,n16442,p3_ir_reg_31_ );
   nand U18287 ( n18945,n16444,n17640 );
   xor U18288 ( n16444,n18950,n18951 );
   xor U18289 ( n18950,p2_datao_reg_15_,p1_datao_reg_15_ );
   or U18290 ( n18942,n15240,n18459 );
   nor U18291 ( n18459,n18836,n18952 );
   nor U18292 ( n18952,n18834,n18835 );
   and U18293 ( n18835,n18953,n15243 );
   xor U18294 ( n18953,n18859,n17554 );
   nand U18295 ( n18834,n18954,n18568,n18955 );
   nand U18296 ( n18955,n18956,n18569 );
   not U18297 ( n18956,n18566 );
   nand U18298 ( n18566,n18957,n15249 );
   not U18299 ( n18957,n18696 );
   nand U18300 ( n18568,n18958,n15246 );
   xor U18301 ( n18958,n18859,n17007 );
   nand U18302 ( n18954,n18573,n18959 );
   nand U18303 ( n18959,n18538,n18960 );
   nand U18304 ( n18960,n18961,n18539 );
   nand U18305 ( n18539,n18542,n16883 );
   not U18306 ( n16883,n15252 );
   nand U18307 ( n18961,n18809,n18962 );
   nand U18308 ( n18962,n18807,n18694 );
   nand U18309 ( n18694,n18963,n16860 );
   not U18310 ( n16860,n15255 );
   xor U18311 ( n18963,n17623,n18755 );
   not U18312 ( n18807,n18811 );
   nand U18313 ( n18811,n18964,n18965 );
   nand U18314 ( n18965,n18602,n18966 );
   or U18315 ( n18966,n18601,n15487 );
   and U18316 ( n18602,n18967,n18968 );
   nand U18317 ( n18968,n18969,n15261 );
   or U18318 ( n18969,n18733,n18732 );
   nand U18319 ( n18967,n18732,n18733 );
   nand U18320 ( n18733,n18970,n18971 );
   nand U18321 ( n18971,n18972,n18973,n18654 );
   not U18322 ( n18654,n18656 );
   and U18323 ( n18970,n18974,n18975,n18976 );
   nand U18324 ( n18975,n18655,n15270,n18972 );
   nand U18325 ( n18974,n18977,n18978 );
   not U18326 ( n18977,n18497 );
   xor U18327 ( n18732,n15489,n18755 );
   nand U18328 ( n15489,n18979,n18980,n18981 );
   nand U18329 ( n18981,si_8_,n17643 );
   nand U18330 ( n18980,n16384,n17657 );
   and U18331 ( n16384,n18982,n16576 );
   xor U18332 ( n18982,n18983,n18984 );
   xor U18333 ( n18983,p2_datao_reg_8_,p1_datao_reg_8_ );
   nand U18334 ( n18979,n18137,n18921 );
   not U18335 ( n18137,n18108 );
   nand U18336 ( n18108,n18985,n18986 );
   or U18337 ( n18986,p3_ir_reg_31_,p3_ir_reg_8_ );
   nand U18338 ( n18985,p3_ir_reg_31_,n18987 );
   nand U18339 ( n18987,n16383,n16382 );
   nand U18340 ( n16382,p3_ir_reg_8_,n18988 );
   nand U18341 ( n18964,n18601,n15487 );
   not U18342 ( n15487,n15258 );
   nand U18343 ( n15258,n18989,n18990,n18991,n18992 );
   nand U18344 ( n18992,n18768,n16861 );
   nand U18345 ( n16861,n18993,n18994 );
   nand U18346 ( n18994,p3_reg3_reg_9_,n18995 );
   nand U18347 ( n18995,n18996,n18729 );
   not U18348 ( n18729,p3_reg3_reg_8_ );
   nand U18349 ( n18991,p3_reg2_reg_9_,n17590 );
   nand U18350 ( n18990,p3_reg1_reg_9_,n17591 );
   nand U18351 ( n18989,p3_reg0_reg_9_,n17592 );
   xor U18352 ( n18601,n17580,n18755 );
   not U18353 ( n17580,n15480 );
   nand U18354 ( n15480,n18997,n18998,n18999 );
   nand U18355 ( n18999,si_9_,n17643 );
   nand U18356 ( n18998,n18070,n18921 );
   not U18357 ( n18070,n17995 );
   nand U18358 ( n17995,n19000,n19001,n19002 );
   nand U18359 ( n19001,n16578,n16392 );
   nand U18360 ( n19000,p3_ir_reg_31_,n16383,p3_ir_reg_9_ );
   not U18361 ( n16383,n16391 );
   nand U18362 ( n18997,n17640,n16393 );
   nand U18363 ( n16393,n19003,n19004,n19005 );
   nand U18364 ( n19005,n19006,n19007 );
   or U18365 ( n19004,n19007,p1_datao_reg_9_,p2_datao_reg_9_ );
   nand U18366 ( n19003,n19008,p2_datao_reg_9_ );
   xor U18367 ( n19008,p1_datao_reg_9_,n19007 );
   and U18368 ( n18809,n19009,n19010 );
   or U18369 ( n19010,n16904,n18859 );
   nand U18370 ( n16904,n17623,n15255 );
   not U18371 ( n17623,n15474 );
   or U18372 ( n19009,n16901,n18755 );
   nand U18373 ( n16901,n15474,n15255 );
   nand U18374 ( n15255,n19011,n19012,n19013,n19014 );
   nand U18375 ( n19014,n18768,n16884 );
   xor U18376 ( n16884,n18803,n18993 );
   not U18377 ( n18993,n19015 );
   nand U18378 ( n19013,p3_reg2_reg_10_,n17590 );
   nand U18379 ( n19012,p3_reg1_reg_10_,n17591 );
   nand U18380 ( n19011,p3_reg0_reg_10_,n17592 );
   nand U18381 ( n15474,n19016,n19017,n19018 );
   nand U18382 ( n19018,si_10_,n17643 );
   nand U18383 ( n19017,n18054,n18921 );
   not U18384 ( n18054,n18028 );
   nand U18385 ( n18028,n19019,n19020 );
   or U18386 ( n19020,p3_ir_reg_10_,p3_ir_reg_31_ );
   nand U18387 ( n19019,p3_ir_reg_31_,n16399 );
   nand U18388 ( n16399,n16408,n19021 );
   nand U18389 ( n19021,p3_ir_reg_10_,n19002 );
   nand U18390 ( n19016,n17640,n16400 );
   xor U18391 ( n16400,n19022,n19023 );
   nand U18392 ( n19023,n19024,n19025 );
   nand U18393 ( n19025,n19026,n19007 );
   xor U18394 ( n19022,p2_datao_reg_10_,n19027 );
   nand U18395 ( n18538,n19028,n15252 );
   nand U18396 ( n15252,n19029,n19030,n19031,n19032 );
   nand U18397 ( n19032,n18768,n16933 );
   nand U18398 ( n16933,n19033,n19034 );
   nand U18399 ( n19034,p3_reg3_reg_11_,n19035 );
   nand U18400 ( n19035,n19015,n18803 );
   nand U18401 ( n19031,p3_reg2_reg_11_,n17590 );
   nand U18402 ( n19030,p3_reg1_reg_11_,n17591 );
   nand U18403 ( n19029,p3_reg0_reg_11_,n17592 );
   not U18404 ( n19028,n18542 );
   xor U18405 ( n18542,n16932,n18755 );
   not U18406 ( n16932,n15464 );
   nand U18407 ( n15464,n19036,n19037,n19038 );
   nand U18408 ( n19038,si_11_,n17643 );
   nand U18409 ( n19037,n16410,n17657 );
   and U18410 ( n16410,n16576,n19039 );
   nand U18411 ( n19039,n19040,n19041,n19042 );
   nand U18412 ( n19042,n19043,n19044 );
   or U18413 ( n19041,n19044,n19045,n19046 );
   nand U18414 ( n19040,n19047,n19046 );
   xor U18415 ( n19047,n19044,n19045 );
   nand U18416 ( n19044,n19048,n19049 );
   nand U18417 ( n19036,n18014,n18921 );
   not U18418 ( n18014,n18002 );
   nand U18419 ( n18002,n19050,n19051,n19052 );
   nand U18420 ( n19051,n16409,n16578 );
   nand U18421 ( n19050,p3_ir_reg_11_,n16408,p3_ir_reg_31_ );
   not U18422 ( n16408,n16407 );
   and U18423 ( n18573,n18571,n18569 );
   nand U18424 ( n18569,n19053,n17582 );
   not U18425 ( n17582,n15246 );
   nand U18426 ( n15246,n19054,n19055,n19056,n19057 );
   nand U18427 ( n19057,n18768,n17008 );
   nand U18428 ( n17008,n19058,n19059 );
   nand U18429 ( n19059,p3_reg3_reg_13_,n19060 );
   nand U18430 ( n19060,n19061,n18689 );
   not U18431 ( n19061,n19033 );
   nand U18432 ( n19056,p3_reg2_reg_13_,n17590 );
   nand U18433 ( n19055,p3_reg1_reg_13_,n17591 );
   nand U18434 ( n19054,p3_reg0_reg_13_,n17592 );
   xor U18435 ( n19053,n17007,n18755 );
   not U18436 ( n17007,n15444 );
   nand U18437 ( n15444,n19062,n19063,n19064 );
   nand U18438 ( n19064,si_13_,n17643 );
   nand U18439 ( n19063,n17914,n18921 );
   not U18440 ( n17914,n17927 );
   nand U18441 ( n17927,n19065,n19066,n19067 );
   nand U18442 ( n19066,n16426,n16578 );
   nand U18443 ( n19065,p3_ir_reg_13_,n16425,p3_ir_reg_31_ );
   nand U18444 ( n19062,n17640,n16427 );
   xor U18445 ( n16427,n19068,n19069 );
   xor U18446 ( n19068,p2_datao_reg_13_,n19070 );
   nand U18447 ( n18571,n18696,n16985 );
   not U18448 ( n16985,n15249 );
   nand U18449 ( n15249,n19071,n19072,n19073,n19074 );
   nand U18450 ( n19074,n18768,n16967 );
   xor U18451 ( n16967,n18689,n19033 );
   not U18452 ( n18689,p3_reg3_reg_12_ );
   nand U18453 ( n19073,p3_reg2_reg_12_,n17590 );
   nand U18454 ( n19072,p3_reg1_reg_12_,n17591 );
   nand U18455 ( n19071,p3_reg0_reg_12_,n17592 );
   xor U18456 ( n18696,n16966,n18755 );
   not U18457 ( n16966,n15454 );
   nand U18458 ( n15454,n19075,n19076,n19077 );
   nand U18459 ( n19077,si_12_,n17643 );
   nand U18460 ( n19076,n16417,n17657 );
   and U18461 ( n16417,n19078,n16576 );
   xor U18462 ( n19078,n19079,n19080 );
   xor U18463 ( n19079,p2_datao_reg_12_,p1_datao_reg_12_ );
   nand U18464 ( n19075,n17956,n18921 );
   not U18465 ( n17956,n17953 );
   nand U18466 ( n17953,n19081,n19082 );
   or U18467 ( n19082,p3_ir_reg_12_,p3_ir_reg_31_ );
   nand U18468 ( n19081,p3_ir_reg_31_,n16416 );
   nand U18469 ( n16416,n16425,n19083 );
   nand U18470 ( n19083,p3_ir_reg_12_,n19052 );
   not U18471 ( n16425,n16424 );
   nand U18472 ( n18836,n19084,n19085 );
   nand U18473 ( n19085,n17556,n18755 );
   not U18474 ( n17556,n15894 );
   nand U18475 ( n15894,n18562,n15437 );
   or U18476 ( n19084,n17041,n18755 );
   nand U18477 ( n17041,n18562,n17554 );
   not U18478 ( n17554,n15437 );
   nand U18479 ( n15437,n19086,n19087,n19088 );
   nand U18480 ( n19088,si_14_,n17643 );
   nand U18481 ( n19087,n17878,n18921 );
   not U18482 ( n17878,n17881 );
   nand U18483 ( n17881,n19089,n19090 );
   or U18484 ( n19090,p3_ir_reg_14_,p3_ir_reg_31_ );
   nand U18485 ( n19089,p3_ir_reg_31_,n16433 );
   nand U18486 ( n16433,n16442,n19091 );
   nand U18487 ( n19091,p3_ir_reg_14_,n19067 );
   not U18488 ( n16442,n16441 );
   nand U18489 ( n19086,n16434,n17640 );
   xor U18490 ( n16434,n19092,n19093 );
   xor U18491 ( n19092,p2_datao_reg_14_,p1_datao_reg_14_ );
   not U18492 ( n18562,n15243 );
   nand U18493 ( n15243,n19094,n19095,n19096,n19097 );
   nand U18494 ( n19097,n18768,n19098 );
   not U18495 ( n19098,n17019 );
   xor U18496 ( n17019,p3_reg3_reg_14_,n19058 );
   nand U18497 ( n19096,p3_reg2_reg_14_,n17590 );
   nand U18498 ( n19095,p3_reg1_reg_14_,n17591 );
   nand U18499 ( n19094,p3_reg0_reg_14_,n17592 );
   nand U18500 ( n15240,n19099,n19100,n19101,n19102 );
   nand U18501 ( n19102,n18768,n17052 );
   nand U18502 ( n17052,n19103,n19104 );
   nand U18503 ( n19104,p3_reg3_reg_15_,n19105 );
   nand U18504 ( n19105,n19106,n18831 );
   not U18505 ( n18831,p3_reg3_reg_14_ );
   nand U18506 ( n19101,p3_reg2_reg_15_,n17590 );
   nand U18507 ( n19100,p3_reg1_reg_15_,n17591 );
   nand U18508 ( n19099,p3_reg0_reg_15_,n17592 );
   nand U18509 ( n18905,n18509,n15231 );
   or U18510 ( n18903,n18509,n15231 );
   nand U18511 ( n15231,n19107,n19108,n19109,n19110 );
   nand U18512 ( n19110,n18768,n17137 );
   xor U18513 ( n17137,p3_reg3_reg_18_,n18914 );
   nand U18514 ( n19109,p3_reg2_reg_18_,n17590 );
   nand U18515 ( n19108,p3_reg1_reg_18_,n17591 );
   nand U18516 ( n19107,p3_reg0_reg_18_,n17592 );
   xor U18517 ( n18509,n15401,n18755 );
   nand U18518 ( n15401,n19111,n19112,n19113 );
   nand U18519 ( n19113,si_18_,n17643 );
   nand U18520 ( n19112,n18921,n17724 );
   not U18521 ( n17724,n17716 );
   nand U18522 ( n17716,n19114,n19115,n19116 );
   nand U18523 ( n19115,n16470,n16578 );
   nand U18524 ( n19114,p3_ir_reg_18_,n16469,p3_ir_reg_31_ );
   nand U18525 ( n19111,n16471,n17640 );
   xor U18526 ( n16471,n19117,n19118 );
   xor U18527 ( n19117,p2_datao_reg_18_,p1_datao_reg_18_ );
   or U18528 ( n18900,n18778,n15397 );
   not U18529 ( n15397,n15228 );
   nand U18530 ( n15228,n19119,n19120,n19121,n19122 );
   nand U18531 ( n19122,n18768,n17183 );
   nand U18532 ( n17183,n18888,n19123 );
   nand U18533 ( n19123,p3_reg3_reg_19_,n19124 );
   nand U18534 ( n19124,n18914,n18507 );
   nand U18535 ( n19121,p3_reg2_reg_19_,n17590 );
   nand U18536 ( n19120,p3_reg1_reg_19_,n17591 );
   nand U18537 ( n19119,p3_reg0_reg_19_,n17592 );
   xor U18538 ( n18778,n15874,n18755 );
   not U18539 ( n15874,n15387 );
   nand U18540 ( n15387,n19125,n19126,n19127 );
   nand U18541 ( n19127,n18921,n17480 );
   nand U18542 ( n19126,n16478,n17640 );
   xor U18543 ( n16478,n19128,n19129 );
   xor U18544 ( n19128,p2_datao_reg_19_,p1_datao_reg_19_ );
   nand U18545 ( n19125,si_19_,n17643 );
   nand U18546 ( n15225,n19130,n19131,n19132,n19133 );
   nand U18547 ( n19133,n18768,n17218 );
   xor U18548 ( n17218,n18582,n18888 );
   not U18549 ( n18582,p3_reg3_reg_20_ );
   nand U18550 ( n19132,p3_reg2_reg_20_,n17590 );
   nand U18551 ( n19131,p3_reg1_reg_20_,n17591 );
   nand U18552 ( n19130,p3_reg0_reg_20_,n17592 );
   nand U18553 ( n18875,n18552,n15219 );
   nand U18554 ( n15219,n19134,n19135,n19136,n19137 );
   nand U18555 ( n19137,n18768,n17264 );
   xor U18556 ( n17264,n18550,n18885 );
   not U18557 ( n18550,p3_reg3_reg_22_ );
   nand U18558 ( n19136,p3_reg2_reg_22_,n17590 );
   nand U18559 ( n19135,p3_reg1_reg_22_,n17591 );
   nand U18560 ( n19134,p3_reg0_reg_22_,n17592 );
   xor U18561 ( n18552,n15366,n18755 );
   nand U18562 ( n15366,n19138,n19139 );
   nand U18563 ( n19139,n16501,n17640 );
   xor U18564 ( n16501,n19140,n19141 );
   xor U18565 ( n19140,p2_datao_reg_22_,p1_datao_reg_22_ );
   nand U18566 ( n19138,si_22_,n17643 );
   nand U18567 ( n18479,n19142,n15207 );
   nand U18568 ( n18855,n19143,n18480,n18476 );
   not U18569 ( n18476,n18680 );
   nand U18570 ( n18680,n19144,n19145 );
   or U18571 ( n19145,n15856,n18859 );
   nand U18572 ( n15856,n18469,n15625 );
   nand U18573 ( n19144,n17391,n18859 );
   not U18574 ( n17391,n17364 );
   nand U18575 ( n17364,n18469,n15340 );
   not U18576 ( n18469,n15210 );
   or U18577 ( n18480,n19142,n15207 );
   nand U18578 ( n15207,n19146,n19147,n19148,n19149 );
   nand U18579 ( n19149,n18768,n17373 );
   nand U18580 ( n17373,n18852,n19150 );
   nand U18581 ( n19150,p3_reg3_reg_26_,n19151 );
   not U18582 ( n18852,n18851 );
   nand U18583 ( n19148,p3_reg2_reg_26_,n17590 );
   nand U18584 ( n19147,p3_reg1_reg_26_,n17591 );
   nand U18585 ( n19146,p3_reg0_reg_26_,n17592 );
   xor U18586 ( n19142,n15329,n18755 );
   nand U18587 ( n15329,n19152,n19153 );
   nand U18588 ( n19153,n16535,n17640 );
   xor U18589 ( n16535,n19154,n19155 );
   xor U18590 ( n19154,p2_datao_reg_26_,p1_datao_reg_26_ );
   nand U18591 ( n19152,si_26_,n17643 );
   nand U18592 ( n19143,n18626,n18681 );
   nand U18593 ( n18681,n19156,n15210 );
   nand U18594 ( n15210,n19157,n19158,n19159,n19160 );
   nand U18595 ( n19160,n18768,n17362 );
   nand U18596 ( n17362,n19151,n19161 );
   nand U18597 ( n19161,p3_reg3_reg_25_,n19162 );
   nand U18598 ( n19162,n19163,n18621 );
   not U18599 ( n18621,p3_reg3_reg_24_ );
   nand U18600 ( n19159,p3_reg2_reg_25_,n17590 );
   nand U18601 ( n19158,p3_reg1_reg_25_,n17591 );
   nand U18602 ( n19157,p3_reg0_reg_25_,n17592 );
   xor U18603 ( n19156,n18859,n15340 );
   not U18604 ( n15340,n15625 );
   nand U18605 ( n15625,n19164,n19165 );
   nand U18606 ( n19165,n16528,n17640 );
   xor U18607 ( n16528,n19166,n19167 );
   xor U18608 ( n19166,p2_datao_reg_25_,p1_datao_reg_25_ );
   nand U18609 ( n19164,si_25_,n17643 );
   nand U18610 ( n18626,n19168,n15213 );
   nand U18611 ( n15213,n19169,n19170,n19171,n19172 );
   nand U18612 ( n19172,n18768,n17335 );
   xor U18613 ( n17335,p3_reg3_reg_24_,n19163 );
   nand U18614 ( n19171,p3_reg2_reg_24_,n17590 );
   nand U18615 ( n19170,p3_reg1_reg_24_,n17591 );
   nand U18616 ( n19169,p3_reg0_reg_24_,n17592 );
   xor U18617 ( n19168,n18859,n15350 );
   not U18618 ( n15350,n15632 );
   nand U18619 ( n15632,n19173,n19174 );
   nand U18620 ( n19174,n16518,n17640 );
   xor U18621 ( n16518,n19175,n19176 );
   xor U18622 ( n19175,p2_datao_reg_24_,p1_datao_reg_24_ );
   nand U18623 ( n19173,si_24_,n17643 );
   and U18624 ( n18854,n18745,n18748 );
   nand U18625 ( n18748,n19177,n15204 );
   xor U18626 ( n19177,n18859,n17440 );
   nand U18627 ( n18745,n19178,n15617 );
   not U18628 ( n15617,n15204 );
   nand U18629 ( n15204,n19179,n19180,n19181,n19182 );
   nand U18630 ( n19182,n18768,n17441 );
   nand U18631 ( n19181,p3_reg2_reg_27_,n17590 );
   nand U18632 ( n19180,p3_reg1_reg_27_,n17591 );
   nand U18633 ( n19179,p3_reg0_reg_27_,n17592 );
   xor U18634 ( n19178,n17440,n18755 );
   not U18635 ( n17440,n15320 );
   nand U18636 ( n15320,n19183,n19184 );
   nand U18637 ( n19184,n16545,n17640 );
   xor U18638 ( n16545,n19185,n18764 );
   nand U18639 ( n18764,n19186,n19187 );
   nand U18640 ( n19187,p2_datao_reg_26_,n19188 );
   or U18641 ( n19188,n19189,n19155 );
   nand U18642 ( n19186,n19155,n19189 );
   nand U18643 ( n19155,n19190,n19191 );
   nand U18644 ( n19191,p2_datao_reg_25_,n19192 );
   or U18645 ( n19192,n19193,n19167 );
   nand U18646 ( n19190,n19167,n19193 );
   nand U18647 ( n19167,n19194,n19195 );
   nand U18648 ( n19195,p2_datao_reg_24_,n19196 );
   or U18649 ( n19196,n19197,n19176 );
   nand U18650 ( n19194,n19176,n19197 );
   nand U18651 ( n19176,n19198,n19199 );
   nand U18652 ( n19199,p2_datao_reg_23_,n19200 );
   or U18653 ( n19200,n19201,n18866 );
   nand U18654 ( n19198,n18866,n19201 );
   nand U18655 ( n18866,n19202,n19203 );
   nand U18656 ( n19203,p2_datao_reg_22_,n19204 );
   or U18657 ( n19204,n19205,n19141 );
   nand U18658 ( n19202,n19141,n19205 );
   nand U18659 ( n19141,n19206,n19207 );
   nand U18660 ( n19207,p2_datao_reg_21_,n19208 );
   or U18661 ( n19208,n19209,n18892 );
   nand U18662 ( n19206,n18892,n19209 );
   nand U18663 ( n18892,n19210,n19211 );
   nand U18664 ( n19211,p2_datao_reg_20_,n19212 );
   or U18665 ( n19212,n19213,n18899 );
   nand U18666 ( n19210,n18899,n19213 );
   nand U18667 ( n18899,n19214,n19215 );
   nand U18668 ( n19215,p2_datao_reg_19_,n19216 );
   or U18669 ( n19216,n19217,n19129 );
   nand U18670 ( n19214,n19129,n19217 );
   nand U18671 ( n19129,n19218,n19219 );
   nand U18672 ( n19219,p2_datao_reg_18_,n19220 );
   or U18673 ( n19220,n19221,n19118 );
   nand U18674 ( n19218,n19118,n19221 );
   nand U18675 ( n19118,n19222,n19223 );
   nand U18676 ( n19223,p2_datao_reg_17_,n19224 );
   or U18677 ( n19224,n19225,n18925 );
   nand U18678 ( n19222,n18925,n19225 );
   nand U18679 ( n18925,n19226,n19227 );
   nand U18680 ( n19227,p2_datao_reg_16_,n19228 );
   or U18681 ( n19228,n19229,n18937 );
   nand U18682 ( n19226,n18937,n19229 );
   nand U18683 ( n18937,n19230,n19231 );
   nand U18684 ( n19231,p2_datao_reg_15_,n19232 );
   or U18685 ( n19232,n19233,n18951 );
   nand U18686 ( n19230,n18951,n19233 );
   nand U18687 ( n18951,n19234,n19235 );
   nand U18688 ( n19235,p2_datao_reg_14_,n19236 );
   or U18689 ( n19236,n19237,n19093 );
   nand U18690 ( n19234,n19093,n19237 );
   nand U18691 ( n19093,n19238,n19239 );
   nand U18692 ( n19239,p2_datao_reg_13_,n19240 );
   nand U18693 ( n19240,p1_datao_reg_13_,n19069 );
   or U18694 ( n19238,n19069,p1_datao_reg_13_ );
   nand U18695 ( n19069,n19241,n19242 );
   nand U18696 ( n19242,n19243,n19244 );
   nand U18697 ( n19243,n19245,n19080 );
   not U18698 ( n19080,n19246 );
   nand U18699 ( n19241,p1_datao_reg_12_,n19246 );
   nor U18700 ( n19246,n19247,n19043 );
   nor U18701 ( n19043,n19046,p1_datao_reg_11_ );
   and U18702 ( n19247,n19248,n19049,n19048 );
   and U18703 ( n19048,n19249,n19250 );
   nand U18704 ( n19250,n19251,n19252 );
   nand U18705 ( n19251,n19027,n19024 );
   not U18706 ( n19024,n19006 );
   nand U18707 ( n19249,p1_datao_reg_10_,n19006 );
   nor U18708 ( n19006,n19253,p2_datao_reg_9_ );
   nand U18709 ( n19049,n19254,n19007,n19026 );
   nand U18710 ( n19026,p2_datao_reg_9_,n19253 );
   nand U18711 ( n19007,n19255,n19256 );
   nand U18712 ( n19256,n19257,n19258 );
   nand U18713 ( n19257,n19259,n18984 );
   not U18714 ( n18984,n19260 );
   nand U18715 ( n19255,p1_datao_reg_8_,n19260 );
   nor U18716 ( n19260,n19261,n19262 );
   and U18717 ( n19261,n19263,n19264,n19265 );
   nand U18718 ( n19263,p1_datao_reg_7_,n19266 );
   nand U18719 ( n19254,p2_datao_reg_10_,n19027 );
   nand U18720 ( n19248,p1_datao_reg_11_,n19046 );
   not U18721 ( n19046,p2_datao_reg_11_ );
   xor U18722 ( n19185,p2_datao_reg_27_,p1_datao_reg_27_ );
   nand U18723 ( n19183,si_27_,n17643 );
   nand U18724 ( n18837,n17441,n18483 );
   nand U18725 ( n18483,n19267,n19268,n19269 );
   nand U18726 ( n19269,n19270,p3_state_reg );
   xor U18727 ( n17441,p3_reg3_reg_27_,n18851 );
   nor U18728 ( n18851,n19151,p3_reg3_reg_26_ );
   or U18729 ( n19151,p3_reg3_reg_24_,p3_reg3_reg_25_,n18871 );
   not U18730 ( n18871,n19163 );
   nor U18731 ( n19163,p3_reg3_reg_22_,p3_reg3_reg_23_,n18885 );
   not U18732 ( n18885,n18874 );
   nor U18733 ( n18874,p3_reg3_reg_20_,p3_reg3_reg_21_,n18888 );
   nand U18734 ( n18888,n18507,n18775,n18914 );
   nor U18735 ( n18914,p3_reg3_reg_16_,p3_reg3_reg_17_,n19103 );
   not U18736 ( n19103,n18917 );
   nor U18737 ( n18917,p3_reg3_reg_14_,p3_reg3_reg_15_,n19058 );
   not U18738 ( n19058,n19106 );
   nor U18739 ( n19106,p3_reg3_reg_12_,p3_reg3_reg_13_,n19033 );
   nand U18740 ( n19033,n18803,n18533,n19015 );
   nor U18741 ( n19015,p3_reg3_reg_8_,p3_reg3_reg_9_,n19271 );
   not U18742 ( n18533,p3_reg3_reg_11_ );
   not U18743 ( n18803,p3_reg3_reg_10_ );
   not U18744 ( n18775,p3_reg3_reg_19_ );
   not U18745 ( n18507,p3_reg3_reg_18_ );
   nand U18746 ( p3_u3153,n19272,n19273,n19274,n19275 );
   nor U18747 ( n19275,n19276,n19277,n19278 );
   nor U18748 ( n19278,n16741,n18470 );
   nor U18749 ( n19277,n15908,n18452 );
   not U18750 ( n15560,n17520 );
   nor U18751 ( n17520,n17659,n18921 );
   nor U18752 ( n17659,n18431,n15937 );
   not U18753 ( n15908,n15261 );
   nand U18754 ( n15261,n19279,n19280,n19281,n19282 );
   nand U18755 ( n19282,n18768,n19283 );
   not U18756 ( n19283,n16830 );
   xor U18757 ( n16830,p3_reg3_reg_8_,n19271 );
   nand U18758 ( n19281,p3_reg2_reg_8_,n17590 );
   nand U18759 ( n19280,p3_reg1_reg_8_,n17591 );
   nand U18760 ( n19279,p3_reg0_reg_8_,n17592 );
   and U18761 ( n19276,p3_u3151,p3_reg3_reg_7_ );
   nand U18762 ( n19274,n16798,n18461 );
   nand U18763 ( n18461,n19267,n19268,n19284 );
   nand U18764 ( n19284,n19270,n15567 );
   and U18765 ( n19270,n17685,n19285 );
   nand U18766 ( n19268,n19286,p3_state_reg );
   nand U18767 ( n19286,n19287,n19288,n19289,n19290 );
   and U18768 ( n19290,n15824,n15938,n16258 );
   nand U18769 ( n16258,n15559,n17480 );
   nand U18770 ( n19289,n15559,n16264 );
   not U18771 ( n15559,n16262 );
   nand U18772 ( n19288,n15803,n19291 );
   nand U18773 ( n19287,n19292,n19285 );
   nand U18774 ( n19267,n15810,n19291 );
   and U18775 ( n15810,n17479,n16260,n15567 );
   not U18776 ( n17479,n15942 );
   nand U18777 ( n19273,n19293,n19294,n18456 );
   nand U18778 ( n19295,n19296,n19297 );
   nand U18779 ( n19297,n15805,n15803 );
   nor U18780 ( n15803,n15576,n15946 );
   not U18781 ( n15805,n19291 );
   nand U18782 ( n19291,n15572,n15582,n15566 );
   nand U18783 ( n19296,n15804,n19292 );
   nand U18784 ( n19292,n19298,n17695,n16634,n16172 );
   nand U18785 ( n16172,n15579,n16257 );
   not U18786 ( n15578,n15580 );
   nand U18787 ( n15580,n15946,n15809 );
   nand U18788 ( n17695,n16705,n15809 );
   not U18789 ( n16705,n16630 );
   not U18790 ( n16260,n15941 );
   nand U18791 ( n15941,n15577,n15943 );
   or U18792 ( n19298,n15576,n16264 );
   nand U18793 ( n15576,n17480,n15809,n15943 );
   nand U18794 ( n19294,n19299,n18497,n19300 );
   xor U18795 ( n19300,n19301,n15264 );
   nand U18796 ( n19299,n18498,n18496 );
   not U18797 ( n18498,n18494 );
   nand U18798 ( n19293,n18976,n19302,n18972 );
   and U18799 ( n18972,n18978,n18496 );
   nand U18800 ( n18496,n18495,n16741 );
   not U18801 ( n16741,n15267 );
   nand U18802 ( n18978,n19301,n15507 );
   not U18803 ( n15507,n15264 );
   nand U18804 ( n19302,n18494,n18497 );
   nand U18805 ( n18497,n19303,n15267 );
   nand U18806 ( n15267,n19304,n19305,n19306,n19307 );
   nand U18807 ( n19307,p3_reg2_reg_6_,n17590 );
   nand U18808 ( n19306,p3_reg1_reg_6_,n17591 );
   nand U18809 ( n19305,p3_reg0_reg_6_,n17592 );
   nand U18810 ( n19304,n18768,n16769 );
   nand U18811 ( n16769,n19308,n19309 );
   nand U18812 ( n19309,p3_reg3_reg_6_,n19310 );
   not U18813 ( n19303,n18495 );
   xor U18814 ( n18495,n17569,n18755 );
   not U18815 ( n17569,n15509 );
   nand U18816 ( n15509,n19311,n19312,n19313 );
   nand U18817 ( n19313,si_6_,n17643 );
   nand U18818 ( n19312,n18211,n18921 );
   not U18819 ( n18211,n18187 );
   nand U18820 ( n18187,n19314,n19315 );
   or U18821 ( n19315,p3_ir_reg_31_,p3_ir_reg_6_ );
   nand U18822 ( n19314,p3_ir_reg_31_,n19316 );
   nand U18823 ( n19316,n16367,n16366 );
   nand U18824 ( n16366,p3_ir_reg_6_,n19317 );
   nand U18825 ( n19311,n17640,n16368 );
   nand U18826 ( n16368,n19318,n19319,n19320 );
   nand U18827 ( n19320,n19321,n19322 );
   nand U18828 ( n19319,n19323,p1_datao_reg_6_,p2_datao_reg_6_ );
   nand U18829 ( n19318,n19324,n19325 );
   xor U18830 ( n19324,n19323,p1_datao_reg_6_ );
   not U18831 ( n19323,n19322 );
   nand U18832 ( n19322,n19326,n19327 );
   nand U18833 ( n19327,n19328,n19329 );
   nand U18834 ( n19328,n19330,n19331 );
   nand U18835 ( n19326,p1_datao_reg_5_,n19332 );
   nand U18836 ( n18494,n18973,n19333 );
   nand U18837 ( n19333,n19334,n18656 );
   nand U18838 ( n18656,n19335,n19336 );
   nand U18839 ( n19336,n19337,n18613 );
   nand U18840 ( n18613,n19338,n18791 );
   nand U18841 ( n18791,n19339,n15783 );
   not U18842 ( n15783,n15276 );
   xor U18843 ( n19339,n16707,n18755 );
   nand U18844 ( n19338,n18788,n18790 );
   nand U18845 ( n18790,n19340,n15276 );
   nand U18846 ( n15276,n19341,n19342,n19343,n19344 );
   nand U18847 ( n19344,p3_reg2_reg_3_,n17590 );
   nand U18848 ( n19343,p3_reg1_reg_3_,n17591 );
   nand U18849 ( n19342,p3_reg0_reg_3_,n17592 );
   nand U18850 ( n19341,n18768,n16708 );
   xor U18851 ( n19340,n18859,n16707 );
   not U18852 ( n16707,n15528 );
   nand U18853 ( n15528,n19345,n19346,n19347 );
   nand U18854 ( n19347,si_3_,n17643 );
   nand U18855 ( n19346,n18326,n18921 );
   not U18856 ( n18326,n18301 );
   nand U18857 ( n18301,n19348,n19349,n19350 );
   nand U18858 ( n19349,n16578,n16344 );
   nand U18859 ( n19348,p3_ir_reg_31_,n16343,p3_ir_reg_3_ );
   nand U18860 ( n19345,n17640,n16345 );
   nand U18861 ( n16345,n19351,n19352,n19353 );
   nand U18862 ( n19353,n19354,n19355 );
   not U18863 ( n19354,n19356 );
   or U18864 ( n19352,n19355,n19357,n19358 );
   nand U18865 ( n19351,n19359,n19358 );
   xor U18866 ( n19359,n19355,n19357 );
   nand U18867 ( n19355,n19360,n19361 );
   nand U18868 ( n19361,n19362,n19363 );
   and U18869 ( n18788,n18795,n19364 );
   nand U18870 ( n19364,n18793,n18523 );
   nand U18871 ( n18523,n18720,n19365 );
   nand U18872 ( n19365,n18719,n18721 );
   nand U18873 ( n18721,n19366,n15796 );
   not U18874 ( n15796,n15282 );
   xor U18875 ( n19366,n16639,n18755 );
   nand U18876 ( n18719,n16610,n19367 );
   nand U18877 ( n19367,n16170,n18755 );
   not U18878 ( n16170,n15561 );
   nand U18879 ( n16610,n15561,n15285 );
   nand U18880 ( n15285,n19368,n19369,n19370,n19371 );
   nand U18881 ( n19371,p3_reg2_reg_0_,n17590 );
   nand U18882 ( n19370,p3_reg1_reg_0_,n17591 );
   nand U18883 ( n19369,p3_reg0_reg_0_,n17592 );
   nand U18884 ( n19368,p3_reg3_reg_0_,n18768 );
   nand U18885 ( n15561,n19372,n19373,n19374 );
   nand U18886 ( n19374,p3_ir_reg_0_,n18921 );
   nand U18887 ( n19373,n17640,n16318 );
   nand U18888 ( n16318,n19375,n19376 );
   nand U18889 ( n19376,p1_datao_reg_0_,n19377 );
   nand U18890 ( n19372,si_0_,n17643 );
   nand U18891 ( n18720,n19378,n15282 );
   nand U18892 ( n15282,n19379,n19380,n19381,n19382 );
   nand U18893 ( n19382,p3_reg2_reg_1_,n17590 );
   nand U18894 ( n19381,p3_reg1_reg_1_,n17591 );
   nand U18895 ( n19380,p3_reg0_reg_1_,n17592 );
   nand U18896 ( n19379,p3_reg3_reg_1_,n18768 );
   xor U18897 ( n19378,n18859,n16639 );
   not U18898 ( n16639,n15548 );
   nand U18899 ( n15548,n19383,n19384,n19385 );
   nand U18900 ( n19385,si_1_,n17643 );
   nand U18901 ( n19384,n18378,n18921 );
   not U18902 ( n18378,n18381 );
   nand U18903 ( n18381,n19386,n19387,n19388 );
   nand U18904 ( n19387,n16327,n16578 );
   nand U18905 ( n19386,p3_ir_reg_1_,p3_ir_reg_0_,p3_ir_reg_31_ );
   nand U18906 ( n19383,n17640,n16328 );
   xor U18907 ( n16328,n19389,n19390 );
   xor U18908 ( n19389,p2_datao_reg_1_,p1_datao_reg_1_ );
   not U18909 ( n18793,n18522 );
   nor U18910 ( n18522,n18524,n15279 );
   nand U18911 ( n18795,n18524,n15279 );
   nand U18912 ( n15279,n19391,n19392,n19393,n19394 );
   nand U18913 ( n19394,p3_reg2_reg_2_,n17590 );
   nand U18914 ( n19393,p3_reg1_reg_2_,n17591 );
   nand U18915 ( n19392,p3_reg0_reg_2_,n17592 );
   nand U18916 ( n19391,p3_reg3_reg_2_,n18768 );
   xor U18917 ( n18524,n15538,n18755 );
   nand U18918 ( n15538,n19395,n19396,n19397 );
   nand U18919 ( n19397,si_2_,n17643 );
   nand U18920 ( n19396,n18355,n18921 );
   not U18921 ( n18355,n18342 );
   nand U18922 ( n18342,n19398,n19399 );
   or U18923 ( n19399,p3_ir_reg_2_,p3_ir_reg_31_ );
   nand U18924 ( n19398,p3_ir_reg_31_,n16334 );
   nand U18925 ( n16334,n16343,n19400 );
   nand U18926 ( n19400,p3_ir_reg_2_,n19388 );
   not U18927 ( n16343,n16342 );
   nand U18928 ( n19395,n17640,n16335 );
   nand U18929 ( n16335,n19401,n19402,n19403 );
   nand U18930 ( n19403,n19404,n19363 );
   or U18931 ( n19402,n19363,p1_datao_reg_2_,p2_datao_reg_2_ );
   nand U18932 ( n19401,n19405,p2_datao_reg_2_ );
   xor U18933 ( n19405,p1_datao_reg_2_,n19363 );
   or U18934 ( n19337,n18612,n17571 );
   nand U18935 ( n19335,n18612,n17571 );
   not U18936 ( n17571,n15273 );
   nand U18937 ( n15273,n19406,n19407,n19408,n19409 );
   nand U18938 ( n19409,n16719,n18768 );
   xor U18939 ( n16719,n16708,p3_reg3_reg_4_ );
   not U18940 ( n16708,p3_reg3_reg_3_ );
   nand U18941 ( n19408,p3_reg2_reg_4_,n17590 );
   nand U18942 ( n19407,p3_reg1_reg_4_,n17591 );
   nand U18943 ( n19406,p3_reg0_reg_4_,n17592 );
   xor U18944 ( n18612,n17568,n18755 );
   not U18945 ( n17568,n15522 );
   nand U18946 ( n15522,n19410,n19411,n19412 );
   nand U18947 ( n19412,si_4_,n17643 );
   nand U18948 ( n19411,n18264,n18921 );
   not U18949 ( n18264,n18267 );
   nand U18950 ( n18267,n19413,n19414 );
   or U18951 ( n19414,p3_ir_reg_31_,p3_ir_reg_4_ );
   nand U18952 ( n19413,p3_ir_reg_31_,n19415 );
   nand U18953 ( n19415,n16351,n16350 );
   nand U18954 ( n16350,p3_ir_reg_4_,n19350 );
   nand U18955 ( n19410,n17640,n16352 );
   xor U18956 ( n16352,n19416,n19417 );
   xor U18957 ( n19416,p2_datao_reg_4_,n19418 );
   nand U18958 ( n19334,n18655,n15270 );
   not U18959 ( n18973,n18653 );
   nor U18960 ( n18653,n18655,n15270 );
   nand U18961 ( n15270,n19419,n19420,n19421,n19422 );
   nand U18962 ( n19422,n18768,n16742 );
   nand U18963 ( n16742,n19310,n19423 );
   nand U18964 ( n19423,p3_reg3_reg_5_,n19424 );
   nand U18965 ( n19421,p3_reg2_reg_5_,n17590 );
   nand U18966 ( n19420,p3_reg1_reg_5_,n17591 );
   nand U18967 ( n19419,p3_reg0_reg_5_,n17592 );
   xor U18968 ( n18655,n15516,n18755 );
   nand U18969 ( n15516,n19425,n19426,n19427 );
   nand U18970 ( n19427,si_5_,n17643 );
   nand U18971 ( n19426,n18247,n18921 );
   not U18972 ( n18247,n18220 );
   nand U18973 ( n18220,n19428,n19429,n19317 );
   nand U18974 ( n19429,n16578,n16360 );
   nand U18975 ( n19428,p3_ir_reg_31_,n16351,p3_ir_reg_5_ );
   not U18976 ( n16351,n16359 );
   nand U18977 ( n19425,n17640,n16361 );
   xor U18978 ( n16361,n19430,n19330 );
   not U18979 ( n19330,n19332 );
   xor U18980 ( n19430,p2_datao_reg_5_,p1_datao_reg_5_ );
   nand U18981 ( n18976,n19431,n15264 );
   nand U18982 ( n15264,n19432,n19433,n19434,n19435 );
   nand U18983 ( n19435,n18768,n16798 );
   nand U18984 ( n16798,n19271,n19436 );
   nand U18985 ( n19436,p3_reg3_reg_7_,n19308 );
   not U18986 ( n19271,n18996 );
   nor U18987 ( n18996,n19308,p3_reg3_reg_7_ );
   or U18988 ( n19308,n19310,p3_reg3_reg_6_ );
   or U18989 ( n19310,n19424,p3_reg3_reg_5_ );
   or U18990 ( n19424,p3_reg3_reg_4_,p3_reg3_reg_3_ );
   nand U18991 ( n19434,p3_reg2_reg_7_,n17590 );
   nand U18992 ( n19433,p3_reg1_reg_7_,n17591 );
   not U18993 ( n19439,n19437 );
   nand U18994 ( n19432,p3_reg0_reg_7_,n17592 );
   nand U18995 ( n19437,n19440,n19441 );
   nand U18996 ( n19441,p3_ir_reg_29_,n16578 );
   nand U18997 ( n19440,p3_ir_reg_31_,n16560 );
   nand U18998 ( n16560,p3_ir_reg_29_,n16577 );
   xor U18999 ( n19438,n16578,n16570 );
   not U19000 ( n16570,p3_ir_reg_30_ );
   not U19001 ( n19431,n19301 );
   xor U19002 ( n19301,n17578,n18755 );
   nand U19003 ( n19442,n16264,n15809,n15570 );
   nand U19004 ( n15942,n15946,n16257 );
   nand U19005 ( n17522,n15946,n15577 );
   not U19006 ( n17578,n15496 );
   nand U19007 ( n19272,n18499,n15496 );
   nand U19008 ( n15496,n19443,n19444,n19445 );
   nand U19009 ( n19445,si_7_,n17643 );
   nand U19010 ( n19444,n18146,n18921 );
   not U19011 ( n18146,n18158 );
   nand U19012 ( n18158,n19446,n19447,n18988 );
   nand U19013 ( n19447,n16578,n16376 );
   nand U19014 ( n19446,p3_ir_reg_31_,n16367,p3_ir_reg_7_ );
   not U19015 ( n16367,n16375 );
   nand U19016 ( n19443,n17640,n16377 );
   nand U19017 ( n16377,n19448,n19449,n19450 );
   nand U19018 ( n19450,n19262,n19451 );
   nor U19019 ( n19262,n19266,p1_datao_reg_7_ );
   or U19020 ( n19449,n19451,n19452,n19266 );
   nand U19021 ( n19448,n19453,n19266 );
   not U19022 ( n19266,p2_datao_reg_7_ );
   xor U19023 ( n19453,n19451,n19452 );
   nand U19024 ( n19451,n19265,n19264 );
   nand U19025 ( n19264,n19332,n19454,n19455 );
   nand U19026 ( n19455,p2_datao_reg_5_,n19331 );
   nand U19027 ( n19332,n19456,n19457 );
   nand U19028 ( n19457,n19458,n19459 );
   not U19029 ( n19459,p2_datao_reg_4_ );
   or U19030 ( n19458,n19417,p1_datao_reg_4_ );
   nand U19031 ( n19456,p1_datao_reg_4_,n19417 );
   nand U19032 ( n19417,n19460,n19461 );
   nand U19033 ( n19461,n19462,n19356 );
   nand U19034 ( n19462,n19360,n19463 );
   nand U19035 ( n19463,p1_datao_reg_3_,n19358 );
   not U19036 ( n19360,n19404 );
   nor U19037 ( n19404,n19464,p2_datao_reg_2_ );
   nand U19038 ( n19460,n19363,n19356,n19362 );
   nand U19039 ( n19362,p2_datao_reg_2_,n19464 );
   nand U19040 ( n19356,p2_datao_reg_3_,n19357 );
   nand U19041 ( n19363,n19465,n19466 );
   nand U19042 ( n19466,n19467,n19468 );
   nand U19043 ( n19467,n19390,n19469 );
   nand U19044 ( n19465,p1_datao_reg_1_,n19375 );
   not U19045 ( n19375,n19390 );
   nor U19046 ( n19390,n19377,p1_datao_reg_0_ );
   not U19047 ( n19377,p2_datao_reg_0_ );
   and U19048 ( n19265,n19470,n19471 );
   nand U19049 ( n19471,n19454,n19329,p1_datao_reg_5_ );
   not U19050 ( n19454,n19321 );
   nor U19051 ( n19321,n19325,p1_datao_reg_6_ );
   nand U19052 ( n19470,p1_datao_reg_6_,n19325 );
   nand U19053 ( n18453,n15567,n19472 );
   nand U19054 ( n19472,n17662,n19473 );
   nand U19055 ( n19473,n17685,n15804 );
   not U19056 ( n15804,n19285 );
   nand U19057 ( n19285,n15570,n15583,n15566 );
   and U19058 ( n15566,n19474,n19475,n19476,n19477 );
   nor U19059 ( n19477,n19478,n19479,n19480,n19481 );
   nor U19060 ( n19481,n16590,n16581 );
   not U19061 ( n16581,p3_d_reg_6_ );
   nor U19062 ( n19480,n16590,n16583 );
   not U19063 ( n16583,p3_d_reg_13_ );
   nor U19064 ( n19479,n16590,n16585 );
   not U19065 ( n16585,p3_d_reg_17_ );
   nor U19066 ( n19478,n19482,n16590 );
   nor U19067 ( n19482,p3_d_reg_22_,p3_d_reg_24_,p3_d_reg_23_ );
   nor U19068 ( n19476,n19483,n19484,n19485,n19486 );
   nor U19069 ( n19486,n16590,n16587 );
   not U19070 ( n16587,p3_d_reg_19_ );
   nor U19071 ( n19485,n16590,n16584 );
   not U19072 ( n16584,p3_d_reg_16_ );
   nor U19073 ( n19484,n19487,n16590 );
   nor U19074 ( n19487,p3_d_reg_7_,p3_d_reg_9_,p3_d_reg_8_ );
   nor U19075 ( n19483,n16590,n16582 );
   not U19076 ( n16582,p3_d_reg_10_ );
   nor U19077 ( n19475,n19488,n19489,n19490,n19491 );
   nor U19078 ( n19491,n16590,n16589 );
   not U19079 ( n16589,p3_d_reg_29_ );
   nor U19080 ( n19490,n16590,n16580 );
   not U19081 ( n16580,p3_d_reg_2_ );
   nor U19082 ( n19489,n16590,n16588 );
   not U19083 ( n16588,p3_d_reg_27_ );
   nor U19084 ( n19488,n16590,n16586 );
   not U19085 ( n16586,p3_d_reg_18_ );
   nor U19086 ( n19474,n19492,n19493,n19494,n19495 );
   nor U19087 ( n19495,n19496,n16590 );
   nor U19088 ( n19496,p3_d_reg_5_,p3_d_reg_4_,p3_d_reg_3_,p3_d_reg_30_ );
   nor U19089 ( n19494,n19497,n16590 );
   nor U19090 ( n19497,p3_d_reg_20_,p3_d_reg_26_,p3_d_reg_25_ );
   nor U19091 ( n19493,n19498,n16590 );
   nor U19092 ( n19498,p3_d_reg_15_,p3_d_reg_14_,p3_d_reg_12_,p3_d_reg_11_ );
   nor U19093 ( n19492,n19499,n16590 );
   nor U19094 ( n19499,p3_d_reg_21_,p3_d_reg_31_,p3_d_reg_28_ );
   not U19095 ( n15583,n15572 );
   nand U19096 ( n15572,n15815,n19500 );
   or U19097 ( n19500,n16590,p3_d_reg_1_ );
   nand U19098 ( n15815,n19501,n19502 );
   not U19099 ( n15570,n15582 );
   nand U19100 ( n15582,n15818,n19503 );
   or U19101 ( n19503,n16590,p3_d_reg_0_ );
   and U19102 ( n19504,n19505,n19502 );
   xor U19103 ( n19505,n19506,n17660 );
   not U19104 ( n17660,p3_b_reg );
   nand U19105 ( n15818,n19506,n19501 );
   and U19106 ( n17685,n19507,n15562 );
   nor U19107 ( n15562,n15943,n16257 );
   nand U19108 ( n19507,n15946,n17480 );
   not U19109 ( n15946,n16264 );
   nand U19110 ( n17662,n15558,n15809 );
   nor U19111 ( n15558,n15577,n15943,n16264 );
   nand U19112 ( n16264,n19508,n19509 );
   nand U19113 ( n19509,p3_ir_reg_20_,n16578 );
   nand U19114 ( n19508,n16483,n16484,p3_ir_reg_31_ );
   nand U19115 ( n16483,p3_ir_reg_20_,n16477 );
   not U19116 ( n15577,n17480 );
   nand U19117 ( n17480,n19510,n19511 );
   nand U19118 ( n19511,p3_ir_reg_19_,n16578 );
   nand U19119 ( n19510,n16476,n16477,p3_ir_reg_31_ );
   nand U19120 ( n16476,p3_ir_reg_19_,n19116 );
   nand U19121 ( p3_u3150,n18443,n19512 );
   nand U19122 ( n19512,n16262,n15938,n17657 );
   not U19123 ( n15938,n18437 );
   nor U19124 ( n18437,n19501,n19506,n19502 );
   nand U19125 ( n19502,n19513,n19514,n19515 );
   nand U19126 ( n19514,n16527,n16578 );
   nand U19127 ( n19513,p3_ir_reg_25_,n16526,p3_ir_reg_31_ );
   nand U19128 ( n19506,n19516,n19517 );
   or U19129 ( n19517,p3_ir_reg_24_,p3_ir_reg_31_ );
   nand U19130 ( n19516,p3_ir_reg_31_,n16517 );
   nand U19131 ( n16517,n16526,n19518 );
   nand U19132 ( n19518,p3_ir_reg_24_,n19519 );
   not U19133 ( n16526,n16525 );
   nand U19134 ( n19501,n19520,n19521 );
   or U19135 ( n19521,p3_ir_reg_26_,p3_ir_reg_31_ );
   nand U19136 ( n19520,p3_ir_reg_31_,n16534 );
   nand U19137 ( n16534,n16543,n19522 );
   nand U19138 ( n19522,p3_ir_reg_26_,n19515 );
   nand U19139 ( n16262,n15943,n16257 );
   not U19140 ( n16257,n15809 );
   nand U19141 ( n15809,n19523,n19524,n19525 );
   nand U19142 ( n19524,n16493,n16578 );
   nand U19143 ( n19523,p3_ir_reg_21_,n16484,p3_ir_reg_31_ );
   not U19144 ( n16484,n16492 );
   not U19145 ( n15943,n15579 );
   nand U19146 ( n15579,n19526,n19527 );
   or U19147 ( n19527,p3_ir_reg_22_,p3_ir_reg_31_ );
   nand U19148 ( n19526,p3_ir_reg_31_,n16500 );
   nand U19149 ( n16500,n16509,n19528 );
   nand U19150 ( n19528,p3_ir_reg_22_,n19525 );
   and U19151 ( n18443,n19529,p3_state_reg );
   nand U19152 ( n19529,n15944,n17657 );
   nand U19153 ( n17657,n15937,n18431 );
   nand U19154 ( n18431,n19530,n19531,n16577 );
   nand U19155 ( n16577,n16552,n16554 );
   not U19156 ( n16552,n16553 );
   nand U19157 ( n19531,n16554,n16578 );
   not U19158 ( n16554,p3_ir_reg_28_ );
   nand U19159 ( n19530,p3_ir_reg_28_,n16553,p3_ir_reg_31_ );
   nand U19160 ( n16553,n16542,n16544 );
   nand U19161 ( n19533,n16544,n16578 );
   not U19162 ( n16544,p3_ir_reg_27_ );
   nand U19163 ( n19532,p3_ir_reg_27_,n16543,p3_ir_reg_31_ );
   not U19164 ( n16543,n16542 );
   nor U19165 ( n16542,n19515,p3_ir_reg_26_ );
   nand U19166 ( n19515,n16525,n16527 );
   not U19167 ( n16527,p3_ir_reg_25_ );
   nor U19168 ( n16525,n19519,p3_ir_reg_24_ );
   not U19169 ( n15944,n15824 );
   nand U19170 ( n15824,n19534,n19535,n19519 );
   nand U19171 ( n19519,n16508,n16510 );
   nand U19172 ( n19535,n16510,n16578 );
   not U19173 ( n16578,p3_ir_reg_31_ );
   not U19174 ( n16510,p3_ir_reg_23_ );
   nand U19175 ( n19534,p3_ir_reg_23_,n16509,p3_ir_reg_31_ );
   not U19176 ( n16509,n16508 );
   nor U19177 ( n16508,n19525,p3_ir_reg_22_ );
   nand U19178 ( n19525,n16492,n16493 );
   not U19179 ( n16493,p3_ir_reg_21_ );
   nor U19180 ( n16492,n16477,p3_ir_reg_20_ );
   or U19181 ( n16477,n19116,p3_ir_reg_19_ );
   nand U19182 ( n19116,n16468,n16470 );
   not U19183 ( n16470,p3_ir_reg_18_ );
   not U19184 ( n16468,n16469 );
   nand U19185 ( n16469,n16458,n16460 );
   not U19186 ( n16460,p3_ir_reg_17_ );
   nor U19187 ( n16458,n18935,p3_ir_reg_16_ );
   nand U19188 ( n18935,n16441,n16443 );
   not U19189 ( n16443,p3_ir_reg_15_ );
   nor U19190 ( n16441,n19067,p3_ir_reg_14_ );
   nand U19191 ( n19067,n16424,n16426 );
   not U19192 ( n16426,p3_ir_reg_13_ );
   nor U19193 ( n16424,n19052,p3_ir_reg_12_ );
   nand U19194 ( n19052,n16407,n16409 );
   not U19195 ( n16409,p3_ir_reg_11_ );
   nor U19196 ( n16407,n19002,p3_ir_reg_10_ );
   nand U19197 ( n19002,n16391,n16392 );
   not U19198 ( n16392,p3_ir_reg_9_ );
   nor U19199 ( n16391,n18988,p3_ir_reg_8_ );
   nand U19200 ( n18988,n16375,n16376 );
   not U19201 ( n16376,p3_ir_reg_7_ );
   nor U19202 ( n16375,n19317,p3_ir_reg_6_ );
   nand U19203 ( n19317,n16359,n16360 );
   not U19204 ( n16360,p3_ir_reg_5_ );
   nor U19205 ( n16359,n19350,p3_ir_reg_4_ );
   nand U19206 ( n19350,n16342,n16344 );
   not U19207 ( n16344,p3_ir_reg_3_ );
   nor U19208 ( n16342,n19388,p3_ir_reg_2_ );
   nand U19209 ( n19388,n16326,n16327 );
   not U19210 ( n16327,p3_ir_reg_1_ );
   not U19211 ( n16326,p3_ir_reg_0_ );
   nand U19212 ( p2_u3562,n19536,n19537 );
   nand U19213 ( n19537,p2_datao_reg_31_,n19538 );
   nand U19214 ( n19536,p2_u3947,n19539 );
   nand U19215 ( p2_u3561,n19540,n19541 );
   nand U19216 ( n19541,p2_datao_reg_30_,n19538 );
   nand U19217 ( n19540,p2_u3947,n19542 );
   nand U19218 ( p2_u3560,n19543,n19544 );
   nand U19219 ( n19544,p2_datao_reg_29_,n19538 );
   nand U19220 ( n19543,p2_u3947,n19545 );
   nand U19221 ( p2_u3559,n19546,n19547 );
   nand U19222 ( n19547,p2_datao_reg_28_,n19538 );
   nand U19223 ( n19546,p2_u3947,n19548 );
   nand U19224 ( p2_u3558,n19549,n19550 );
   nand U19225 ( n19550,p2_datao_reg_27_,n19538 );
   nand U19226 ( n19549,p2_u3947,n19551 );
   nand U19227 ( p2_u3557,n19552,n19553 );
   nand U19228 ( n19553,p2_datao_reg_26_,n19538 );
   nand U19229 ( n19552,p2_u3947,n19554 );
   nand U19230 ( p2_u3556,n19555,n19556 );
   nand U19231 ( n19556,p2_datao_reg_25_,n19538 );
   nand U19232 ( n19555,p2_u3947,n19557 );
   nand U19233 ( p2_u3555,n19558,n19559 );
   nand U19234 ( n19559,p2_datao_reg_24_,n19538 );
   nand U19235 ( n19558,p2_u3947,n19560 );
   nand U19236 ( p2_u3554,n19561,n19562 );
   nand U19237 ( n19562,p2_datao_reg_23_,n19538 );
   nand U19238 ( n19561,p2_u3947,n19563 );
   nand U19239 ( p2_u3553,n19564,n19565 );
   nand U19240 ( n19565,p2_datao_reg_22_,n19538 );
   nand U19241 ( n19564,p2_u3947,n19566 );
   nand U19242 ( p2_u3552,n19567,n19568 );
   nand U19243 ( n19568,p2_datao_reg_21_,n19538 );
   nand U19244 ( n19567,p2_u3947,n19569 );
   nand U19245 ( p2_u3551,n19570,n19571 );
   nand U19246 ( n19571,p2_datao_reg_20_,n19538 );
   nand U19247 ( n19570,p2_u3947,n19572 );
   nand U19248 ( p2_u3550,n19573,n19574 );
   nand U19249 ( n19574,p2_datao_reg_19_,n19538 );
   nand U19250 ( n19573,p2_u3947,n19575 );
   nand U19251 ( p2_u3549,n19576,n19577 );
   nand U19252 ( n19577,p2_datao_reg_18_,n19538 );
   nand U19253 ( n19576,p2_u3947,n19578 );
   nand U19254 ( p2_u3548,n19579,n19580 );
   nand U19255 ( n19580,p2_datao_reg_17_,n19538 );
   nand U19256 ( n19579,p2_u3947,n19581 );
   nand U19257 ( p2_u3547,n19582,n19583 );
   nand U19258 ( n19583,p2_datao_reg_16_,n19538 );
   nand U19259 ( n19582,p2_u3947,n19584 );
   nand U19260 ( p2_u3546,n19585,n19586 );
   nand U19261 ( n19586,p2_datao_reg_15_,n19538 );
   nand U19262 ( n19585,p2_u3947,n19587 );
   nand U19263 ( p2_u3545,n19588,n19589 );
   nand U19264 ( n19589,p2_datao_reg_14_,n19538 );
   nand U19265 ( n19588,p2_u3947,n19590 );
   nand U19266 ( p2_u3544,n19591,n19592 );
   nand U19267 ( n19592,p2_datao_reg_13_,n19538 );
   nand U19268 ( n19591,p2_u3947,n19593 );
   nand U19269 ( p2_u3543,n19594,n19595 );
   nand U19270 ( n19595,p2_datao_reg_12_,n19538 );
   nand U19271 ( n19594,p2_u3947,n19596 );
   nand U19272 ( p2_u3542,n19597,n19598 );
   nand U19273 ( n19598,p2_datao_reg_11_,n19538 );
   nand U19274 ( n19597,p2_u3947,n19599 );
   nand U19275 ( p2_u3541,n19600,n19601 );
   nand U19276 ( n19601,p2_datao_reg_10_,n19538 );
   nand U19277 ( n19600,p2_u3947,n19602 );
   nand U19278 ( p2_u3540,n19603,n19604 );
   nand U19279 ( n19604,p2_datao_reg_9_,n19538 );
   nand U19280 ( n19603,p2_u3947,n19605 );
   nand U19281 ( p2_u3539,n19606,n19607 );
   nand U19282 ( n19607,p2_datao_reg_8_,n19538 );
   nand U19283 ( n19606,p2_u3947,n19608 );
   nand U19284 ( p2_u3538,n19609,n19610 );
   nand U19285 ( n19610,p2_datao_reg_7_,n19538 );
   nand U19286 ( n19609,p2_u3947,n19611 );
   nand U19287 ( p2_u3537,n19612,n19613 );
   nand U19288 ( n19613,p2_datao_reg_6_,n19538 );
   nand U19289 ( n19612,p2_u3947,n19614 );
   nand U19290 ( p2_u3536,n19615,n19616 );
   nand U19291 ( n19616,p2_datao_reg_5_,n19538 );
   nand U19292 ( n19615,p2_u3947,n19617 );
   nand U19293 ( p2_u3535,n19618,n19619 );
   nand U19294 ( n19619,p2_datao_reg_4_,n19538 );
   nand U19295 ( n19618,p2_u3947,n19620 );
   nand U19296 ( p2_u3534,n19621,n19622 );
   nand U19297 ( n19622,p2_datao_reg_3_,n19538 );
   nand U19298 ( n19621,p2_u3947,n19623 );
   nand U19299 ( p2_u3533,n19624,n19625 );
   nand U19300 ( n19625,p2_datao_reg_2_,n19538 );
   nand U19301 ( n19624,p2_u3947,n19626 );
   nand U19302 ( p2_u3532,n19627,n19628 );
   nand U19303 ( n19628,p2_datao_reg_1_,n19538 );
   nand U19304 ( n19627,p2_u3947,n19629 );
   nand U19305 ( p2_u3531,n19630,n19631 );
   nand U19306 ( n19631,p2_datao_reg_0_,n19538 );
   nand U19307 ( n19630,p2_u3947,n19632 );
   nand U19308 ( p2_u3530,n19633,n19634 );
   nand U19309 ( n19634,n19635,n19636 );
   nand U19310 ( n19633,p2_reg1_reg_31_,n19637 );
   nand U19311 ( p2_u3529,n19638,n19639 );
   nand U19312 ( n19639,p2_reg1_reg_30_,n19637 );
   nand U19313 ( n19638,n19635,n19640 );
   nand U19314 ( p2_u3528,n19641,n19642 );
   nand U19315 ( n19642,p2_reg1_reg_29_,n19637 );
   nand U19316 ( n19641,n19635,n19643 );
   nand U19317 ( p2_u3527,n19644,n19645 );
   nand U19318 ( n19645,p2_reg1_reg_28_,n19637 );
   nand U19319 ( n19644,n19635,n19646 );
   nand U19320 ( p2_u3526,n19647,n19648 );
   nand U19321 ( n19648,p2_reg1_reg_27_,n19637 );
   nand U19322 ( n19647,n19635,n19649 );
   nand U19323 ( p2_u3525,n19650,n19651 );
   nand U19324 ( n19651,p2_reg1_reg_26_,n19637 );
   nand U19325 ( n19650,n19635,n19652 );
   nand U19326 ( p2_u3524,n19653,n19654 );
   nand U19327 ( n19654,p2_reg1_reg_25_,n19637 );
   nand U19328 ( n19653,n19635,n19655 );
   nand U19329 ( p2_u3523,n19656,n19657 );
   nand U19330 ( n19657,p2_reg1_reg_24_,n19637 );
   nand U19331 ( n19656,n19635,n19658 );
   nand U19332 ( p2_u3522,n19659,n19660 );
   nand U19333 ( n19660,p2_reg1_reg_23_,n19637 );
   nand U19334 ( n19659,n19635,n19661 );
   nand U19335 ( p2_u3521,n19662,n19663 );
   nand U19336 ( n19663,p2_reg1_reg_22_,n19637 );
   nand U19337 ( n19662,n19635,n19664 );
   nand U19338 ( p2_u3520,n19665,n19666 );
   nand U19339 ( n19666,p2_reg1_reg_21_,n19637 );
   nand U19340 ( n19665,n19635,n19667 );
   nand U19341 ( p2_u3519,n19668,n19669 );
   nand U19342 ( n19669,p2_reg1_reg_20_,n19637 );
   nand U19343 ( n19668,n19635,n19670 );
   nand U19344 ( p2_u3518,n19671,n19672 );
   nand U19345 ( n19672,p2_reg1_reg_19_,n19637 );
   nand U19346 ( n19671,n19635,n19673 );
   nand U19347 ( p2_u3517,n19674,n19675 );
   nand U19348 ( n19675,p2_reg1_reg_18_,n19637 );
   nand U19349 ( n19674,n19635,n19676 );
   nand U19350 ( p2_u3516,n19677,n19678 );
   nand U19351 ( n19678,p2_reg1_reg_17_,n19637 );
   nand U19352 ( n19677,n19635,n19679 );
   nand U19353 ( p2_u3515,n19680,n19681 );
   nand U19354 ( n19681,p2_reg1_reg_16_,n19637 );
   nand U19355 ( n19680,n19635,n19682 );
   nand U19356 ( p2_u3514,n19683,n19684 );
   nand U19357 ( n19684,p2_reg1_reg_15_,n19637 );
   nand U19358 ( n19683,n19635,n19685 );
   nand U19359 ( p2_u3513,n19686,n19687 );
   nand U19360 ( n19687,p2_reg1_reg_14_,n19637 );
   nand U19361 ( n19686,n19635,n19688 );
   nand U19362 ( p2_u3512,n19689,n19690 );
   nand U19363 ( n19690,p2_reg1_reg_13_,n19637 );
   nand U19364 ( n19689,n19635,n19691 );
   nand U19365 ( p2_u3511,n19692,n19693 );
   nand U19366 ( n19693,p2_reg1_reg_12_,n19637 );
   nand U19367 ( n19692,n19635,n19694 );
   nand U19368 ( p2_u3510,n19695,n19696 );
   nand U19369 ( n19696,p2_reg1_reg_11_,n19637 );
   nand U19370 ( n19695,n19635,n19697 );
   nand U19371 ( p2_u3509,n19698,n19699 );
   nand U19372 ( n19699,p2_reg1_reg_10_,n19637 );
   nand U19373 ( n19698,n19635,n19700 );
   nand U19374 ( p2_u3508,n19701,n19702 );
   nand U19375 ( n19702,p2_reg1_reg_9_,n19637 );
   nand U19376 ( n19701,n19635,n19703 );
   nand U19377 ( p2_u3507,n19704,n19705 );
   nand U19378 ( n19705,p2_reg1_reg_8_,n19637 );
   nand U19379 ( n19704,n19635,n19706 );
   nand U19380 ( p2_u3506,n19707,n19708 );
   nand U19381 ( n19708,p2_reg1_reg_7_,n19637 );
   nand U19382 ( n19707,n19635,n19709 );
   nand U19383 ( p2_u3505,n19710,n19711 );
   nand U19384 ( n19711,p2_reg1_reg_6_,n19637 );
   nand U19385 ( n19710,n19635,n19712 );
   nand U19386 ( p2_u3504,n19713,n19714 );
   nand U19387 ( n19714,p2_reg1_reg_5_,n19637 );
   nand U19388 ( n19713,n19635,n19715 );
   nand U19389 ( p2_u3503,n19716,n19717 );
   nand U19390 ( n19717,p2_reg1_reg_4_,n19637 );
   nand U19391 ( n19716,n19635,n19718 );
   nand U19392 ( p2_u3502,n19719,n19720 );
   nand U19393 ( n19720,p2_reg1_reg_3_,n19637 );
   nand U19394 ( n19719,n19635,n19721 );
   nand U19395 ( p2_u3501,n19722,n19723 );
   nand U19396 ( n19723,p2_reg1_reg_2_,n19637 );
   nand U19397 ( n19722,n19635,n19724 );
   nand U19398 ( p2_u3500,n19725,n19726 );
   nand U19399 ( n19726,p2_reg1_reg_1_,n19637 );
   nand U19400 ( n19725,n19635,n19727 );
   nand U19401 ( p2_u3499,n19728,n19729 );
   nand U19402 ( n19729,p2_reg1_reg_0_,n19637 );
   nand U19403 ( n19728,n19635,n19730 );
   nand U19404 ( p2_u3498,n19733,n19734 );
   nand U19405 ( n19734,n19735,n19636 );
   nand U19406 ( n19636,n19736,n19737,n19738 );
   nand U19407 ( n19738,n19739,n19740 );
   nand U19408 ( n19736,n19741,n19742 );
   nand U19409 ( n19733,p2_reg0_reg_31_,n19743 );
   nand U19410 ( p2_u3497,n19744,n19745 );
   nand U19411 ( n19745,n19735,n19640 );
   nand U19412 ( n19640,n19746,n19737,n19747 );
   nand U19413 ( n19747,n19748,n19739 );
   not U19414 ( n19737,n19749 );
   nand U19415 ( n19746,n19750,n19751,n19741 );
   nand U19416 ( n19744,p2_reg0_reg_30_,n19743 );
   nand U19417 ( p2_u3496,n19752,n19753 );
   nand U19418 ( n19753,n19735,n19643 );
   nand U19419 ( n19643,n19754,n19755,n19756,n19757 );
   or U19420 ( n19757,n19758,n19759 );
   or U19421 ( n19756,n19760,n19761 );
   nand U19422 ( n19755,n19762,n19739 );
   not U19423 ( n19754,n19763 );
   nand U19424 ( n19752,p2_reg0_reg_29_,n19743 );
   nand U19425 ( p2_u3495,n19764,n19765 );
   nand U19426 ( n19765,n19735,n19646 );
   nand U19427 ( n19646,n19766,n19767,n19768,n19769 );
   nor U19428 ( n19769,n19770,n19771,n19772 );
   nor U19429 ( n19772,n19773,n19774 );
   nor U19430 ( n19771,n19775,n19776 );
   nor U19431 ( n19770,n19777,n19778 );
   nand U19432 ( n19768,n19779,n19741 );
   or U19433 ( n19766,n19780,n19781 );
   nand U19434 ( n19764,p2_reg0_reg_28_,n19743 );
   nand U19435 ( p2_u3494,n19782,n19783 );
   nand U19436 ( n19783,n19735,n19649 );
   nand U19437 ( n19649,n19784,n19785,n19786 );
   nor U19438 ( n19786,n19787,n19788,n19789 );
   nor U19439 ( n19789,n19760,n19790 );
   nor U19440 ( n19788,n19759,n19791 );
   nor U19441 ( n19787,n19792,n19774 );
   nand U19442 ( n19785,n19793,n19739 );
   nand U19443 ( n19782,p2_reg0_reg_27_,n19743 );
   nand U19444 ( p2_u3493,n19794,n19795 );
   nand U19445 ( n19795,n19735,n19652 );
   nand U19446 ( n19652,n19796,n19797,n19798 );
   nor U19447 ( n19798,n19799,n19800,n19801 );
   nor U19448 ( n19801,n19759,n19802 );
   nor U19449 ( n19800,n19760,n19803 );
   nor U19450 ( n19799,n19775,n19774 );
   nand U19451 ( n19797,n19804,n19739 );
   nand U19452 ( n19794,p2_reg0_reg_26_,n19743 );
   nand U19453 ( p2_u3492,n19805,n19806 );
   nand U19454 ( n19806,n19735,n19655 );
   nand U19455 ( n19655,n19807,n19808,n19809,n19810 );
   nor U19456 ( n19810,n19811,n19812,n19813 );
   nor U19457 ( n19813,n19814,n19774 );
   nor U19458 ( n19812,n19815,n19776 );
   nor U19459 ( n19811,n19777,n19816 );
   nand U19460 ( n19809,n19817,n19818 );
   nand U19461 ( n19808,n19819,n19741 );
   nand U19462 ( n19807,n19820,n19821 );
   nand U19463 ( n19805,p2_reg0_reg_25_,n19743 );
   nand U19464 ( p2_u3491,n19822,n19823 );
   nand U19465 ( n19823,n19735,n19658 );
   nand U19466 ( n19658,n19824,n19825,n19826,n19827 );
   nor U19467 ( n19827,n19828,n19829,n19830 );
   nor U19468 ( n19830,n19831,n19774 );
   nor U19469 ( n19829,n19832,n19776 );
   nor U19470 ( n19828,n19777,n19833 );
   or U19471 ( n19826,n19834,n19759 );
   nand U19472 ( n19825,n19835,n19821 );
   nand U19473 ( n19824,n19836,n19818 );
   nand U19474 ( n19822,p2_reg0_reg_24_,n19743 );
   nand U19475 ( p2_u3490,n19837,n19838 );
   nand U19476 ( n19838,n19735,n19661 );
   nand U19477 ( n19661,n19839,n19840,n19841 );
   nor U19478 ( n19841,n19842,n19843,n19844 );
   nor U19479 ( n19844,n19760,n19845 );
   nor U19480 ( n19843,n19759,n19846 );
   nor U19481 ( n19842,n19815,n19774 );
   nand U19482 ( n19840,n19847,n19739 );
   nand U19483 ( n19837,p2_reg0_reg_23_,n19743 );
   nand U19484 ( p2_u3489,n19848,n19849 );
   nand U19485 ( n19849,n19735,n19664 );
   nand U19486 ( n19664,n19850,n19851,n19852,n19853 );
   nor U19487 ( n19853,n19854,n19855,n19856 );
   nor U19488 ( n19856,n19832,n19774 );
   nor U19489 ( n19855,n19857,n19776 );
   nor U19490 ( n19854,n19777,n19858 );
   or U19491 ( n19852,n19859,n19759 );
   nand U19492 ( n19850,n19860,n19821 );
   nand U19493 ( n19848,p2_reg0_reg_22_,n19743 );
   nand U19494 ( p2_u3488,n19861,n19862 );
   nand U19495 ( n19862,n19735,n19667 );
   nand U19496 ( n19667,n19863,n19864,n19865 );
   nor U19497 ( n19865,n19866,n19867,n19868 );
   nor U19498 ( n19868,n19760,n19869 );
   nor U19499 ( n19867,n19759,n19870 );
   nor U19500 ( n19866,n19871,n19774 );
   nand U19501 ( n19864,n19872,n19739 );
   nand U19502 ( n19861,p2_reg0_reg_21_,n19743 );
   nand U19503 ( p2_u3487,n19873,n19874 );
   nand U19504 ( n19874,n19735,n19670 );
   nand U19505 ( n19670,n19875,n19876,n19877 );
   nor U19506 ( n19877,n19878,n19879,n19880 );
   nor U19507 ( n19880,n19759,n19881 );
   nor U19508 ( n19879,n19760,n19882 );
   nor U19509 ( n19878,n19857,n19774 );
   nand U19510 ( n19876,n19883,n19739 );
   nand U19511 ( n19873,p2_reg0_reg_20_,n19743 );
   nand U19512 ( p2_u3486,n19884,n19885 );
   nand U19513 ( n19885,n19735,n19673 );
   nand U19514 ( n19673,n19886,n19887,n19888,n19889 );
   nor U19515 ( n19889,n19890,n19891 );
   nor U19516 ( n19890,n19777,n19892 );
   nand U19517 ( n19888,n19893,n19572 );
   nand U19518 ( n19887,n19894,n19741 );
   nand U19519 ( n19886,n19895,n19896 );
   nand U19520 ( n19884,p2_reg0_reg_19_,n19743 );
   nand U19521 ( p2_u3484,n19897,n19898 );
   nand U19522 ( n19898,n19735,n19676 );
   nand U19523 ( n19676,n19899,n19900,n19901,n19902 );
   nor U19524 ( n19902,n19903,n19904,n19905 );
   nor U19525 ( n19905,n19906,n19774 );
   nor U19526 ( n19904,n19907,n19776 );
   nor U19527 ( n19903,n19777,n19908 );
   or U19528 ( n19901,n19909,n19759 );
   or U19529 ( n19900,n19910,n19781 );
   nand U19530 ( n19899,n19911,n19818 );
   nand U19531 ( n19897,p2_reg0_reg_18_,n19743 );
   nand U19532 ( p2_u3481,n19912,n19913 );
   nand U19533 ( n19913,n19735,n19679 );
   nand U19534 ( n19679,n19914,n19915,n19916 );
   nor U19535 ( n19916,n19917,n19918,n19919 );
   nor U19536 ( n19919,n19760,n19920 );
   nor U19537 ( n19918,n19759,n19921 );
   nor U19538 ( n19917,n19922,n19774 );
   nand U19539 ( n19915,n19923,n19739 );
   nand U19540 ( n19912,p2_reg0_reg_17_,n19743 );
   nand U19541 ( p2_u3478,n19924,n19925 );
   nand U19542 ( n19925,n19735,n19682 );
   nand U19543 ( n19682,n19926,n19927,n19928 );
   nor U19544 ( n19928,n19929,n19930,n19931 );
   nor U19545 ( n19931,n19759,n19932 );
   nor U19546 ( n19930,n19933,n19760 );
   nor U19547 ( n19929,n19907,n19774 );
   nand U19548 ( n19927,n19934,n19739 );
   nand U19549 ( n19924,p2_reg0_reg_16_,n19743 );
   nand U19550 ( p2_u3475,n19935,n19936 );
   nand U19551 ( n19936,n19735,n19685 );
   nand U19552 ( n19685,n19937,n19938,n19939,n19940 );
   nor U19553 ( n19940,n19941,n19942,n19943 );
   nor U19554 ( n19943,n19944,n19774 );
   nor U19555 ( n19942,n19945,n19776 );
   nor U19556 ( n19941,n19946,n19777 );
   nand U19557 ( n19939,n19947,n19821 );
   nand U19558 ( n19937,n19741,n19948 );
   nand U19559 ( n19935,p2_reg0_reg_15_,n19743 );
   nand U19560 ( p2_u3472,n19949,n19950 );
   nand U19561 ( n19950,n19735,n19688 );
   nand U19562 ( n19688,n19951,n19952,n19953,n19954 );
   nor U19563 ( n19954,n19955,n19956,n19957 );
   nor U19564 ( n19957,n19958,n19777 );
   nor U19565 ( n19956,n19959,n19774 );
   nand U19566 ( n19953,n19960,n19593 );
   or U19567 ( n19952,n19961,n19781 );
   or U19568 ( n19951,n19962,n19759 );
   nand U19569 ( n19949,p2_reg0_reg_14_,n19743 );
   nand U19570 ( p2_u3469,n19963,n19964 );
   nand U19571 ( n19964,n19735,n19691 );
   nand U19572 ( n19691,n19965,n19966,n19967 );
   nor U19573 ( n19967,n19968,n19969,n19970 );
   nor U19574 ( n19970,n19760,n19971 );
   nor U19575 ( n19969,n19759,n19972 );
   nor U19576 ( n19968,n19945,n19774 );
   nand U19577 ( n19966,n19973,n19739 );
   nand U19578 ( n19963,p2_reg0_reg_13_,n19743 );
   nand U19579 ( p2_u3466,n19974,n19975 );
   nand U19580 ( n19975,n19735,n19694 );
   nand U19581 ( n19694,n19976,n19977,n19978,n19979 );
   nor U19582 ( n19979,n19980,n19981,n19982 );
   nor U19583 ( n19982,n19983,n19774 );
   nor U19584 ( n19981,n19984,n19776 );
   nor U19585 ( n19980,n19777,n19985 );
   or U19586 ( n19978,n19986,n19759 );
   or U19587 ( n19977,n19987,n19781 );
   nand U19588 ( n19976,n19988,n19818 );
   nand U19589 ( n19974,p2_reg0_reg_12_,n19743 );
   nand U19590 ( p2_u3463,n19989,n19990 );
   nand U19591 ( n19990,n19735,n19697 );
   nand U19592 ( n19697,n19991,n19992,n19993 );
   nor U19593 ( n19993,n19994,n19995,n19996 );
   nor U19594 ( n19996,n19760,n19997 );
   nor U19595 ( n19995,n19759,n19998 );
   nor U19596 ( n19994,n19999,n19774 );
   nand U19597 ( n19992,n20000,n19739 );
   nand U19598 ( n19989,p2_reg0_reg_11_,n19743 );
   nand U19599 ( p2_u3460,n20001,n20002 );
   nand U19600 ( n20002,n19735,n19700 );
   nand U19601 ( n19700,n20003,n20004,n20005 );
   nor U19602 ( n20005,n20006,n20007,n20008 );
   nor U19603 ( n20008,n19759,n20009 );
   nor U19604 ( n20007,n19760,n20010 );
   nor U19605 ( n20006,n19984,n19774 );
   nand U19606 ( n20004,n19739,n20011 );
   nand U19607 ( n20001,p2_reg0_reg_10_,n19743 );
   nand U19608 ( p2_u3457,n20012,n20013 );
   nand U19609 ( n20013,n19735,n19703 );
   nand U19610 ( n19703,n20014,n20015,n20016,n20017 );
   nor U19611 ( n20017,n20018,n20019,n20020 );
   nor U19612 ( n20020,n20021,n19774 );
   nor U19613 ( n20019,n20022,n19776 );
   nor U19614 ( n20018,n19777,n20023 );
   nand U19615 ( n20016,n20024,n19818 );
   nand U19616 ( n20015,n20025,n19741 );
   or U19617 ( n20014,n20026,n19781 );
   nand U19618 ( n20012,p2_reg0_reg_9_,n19743 );
   nand U19619 ( p2_u3454,n20027,n20028 );
   nand U19620 ( n20028,n19735,n19706 );
   nand U19621 ( n19706,n20029,n20030,n20031 );
   nor U19622 ( n20031,n20032,n20033,n20034 );
   nor U19623 ( n20034,n19759,n20035 );
   nor U19624 ( n20033,n20036,n19760 );
   nor U19625 ( n20032,n20037,n19774 );
   nand U19626 ( n20030,n20038,n19739 );
   nand U19627 ( n20027,p2_reg0_reg_8_,n19743 );
   nand U19628 ( p2_u3451,n20039,n20040 );
   nand U19629 ( n20040,n19735,n19709 );
   nand U19630 ( n19709,n20041,n20042,n20043 );
   nor U19631 ( n20043,n20044,n20045,n20046 );
   nor U19632 ( n20046,n19760,n20047 );
   nor U19633 ( n20045,n19759,n20048 );
   nor U19634 ( n20044,n20022,n19774 );
   nand U19635 ( n20042,n20049,n19739 );
   nand U19636 ( n20039,p2_reg0_reg_7_,n19743 );
   nand U19637 ( p2_u3448,n20050,n20051 );
   nand U19638 ( n20051,n19735,n19712 );
   nand U19639 ( n19712,n20052,n20053,n20054 );
   nor U19640 ( n20054,n20055,n20056,n20057 );
   nor U19641 ( n20057,n19759,n20058 );
   nor U19642 ( n20056,n20059,n19760 );
   nor U19643 ( n20055,n20060,n19774 );
   nand U19644 ( n20053,n19739,n20061 );
   nand U19645 ( n20050,p2_reg0_reg_6_,n19743 );
   nand U19646 ( p2_u3445,n20062,n20063 );
   nand U19647 ( n20063,n19735,n19715 );
   nand U19648 ( n19715,n20064,n20065,n20066,n20067 );
   nand U19649 ( n20067,n19893,n19614 );
   nor U19650 ( n20066,n20068,n20069 );
   nor U19651 ( n20069,n20070,n19760 );
   nor U19652 ( n20068,n19759,n20071 );
   nand U19653 ( n20065,n20072,n19739 );
   nand U19654 ( n20062,p2_reg0_reg_5_,n19743 );
   nand U19655 ( p2_u3442,n20073,n20074 );
   nand U19656 ( n20074,n19735,n19718 );
   nand U19657 ( n19718,n20075,n20076,n20077,n20078 );
   nor U19658 ( n20078,n20079,n20080,n20081 );
   nor U19659 ( n20081,n20082,n19774 );
   nor U19660 ( n20080,n20083,n19776 );
   nor U19661 ( n20079,n19777,n20084 );
   or U19662 ( n20077,n20085,n19759 );
   nand U19663 ( n20076,n20086,n19821 );
   nand U19664 ( n20075,n20087,n19818 );
   nand U19665 ( n20073,p2_reg0_reg_4_,n19743 );
   nand U19666 ( p2_u3439,n20088,n20089 );
   nand U19667 ( n20089,n19735,n19721 );
   nand U19668 ( n19721,n20090,n20091,n20092,n20093 );
   nor U19669 ( n20093,n20094,n20095,n20096 );
   nor U19670 ( n20096,n19781,n20097 );
   nor U19671 ( n20095,n19759,n20098 );
   nor U19672 ( n20094,n20099,n19776 );
   nand U19673 ( n20091,n19893,n19620 );
   nand U19674 ( n20090,n20100,n19739 );
   nand U19675 ( n20088,p2_reg0_reg_3_,n19743 );
   nand U19676 ( p2_u3436,n20101,n20102 );
   nand U19677 ( n20102,n19735,n19724 );
   nand U19678 ( n19724,n20103,n20104,n20105,n20106 );
   nor U19679 ( n20106,n20107,n20108,n20109 );
   nor U19680 ( n20109,n20110,n19777 );
   nor U19681 ( n20108,n20083,n19774 );
   nand U19682 ( n20105,n19960,n19629 );
   or U19683 ( n20104,n20111,n19781 );
   not U19684 ( n19781,n19821 );
   or U19685 ( n20103,n20112,n19759 );
   nand U19686 ( n20101,p2_reg0_reg_2_,n19743 );
   nand U19687 ( p2_u3433,n20113,n20114 );
   nand U19688 ( n20114,n19735,n19727 );
   nand U19689 ( n19727,n20115,n20116,n20117,n20118 );
   nor U19690 ( n20118,n20119,n20120,n20121 );
   nor U19691 ( n20121,n20099,n19774 );
   nor U19692 ( n20120,n20122,n19776 );
   nor U19693 ( n20119,n20123,n19777 );
   nand U19694 ( n20117,n20124,n19818 );
   nand U19695 ( n20116,n19741,n20125 );
   nand U19696 ( n20115,n20126,n19821 );
   nand U19697 ( n19821,n20127,n19760 );
   nand U19698 ( n20113,p2_reg0_reg_1_,n19743 );
   nand U19699 ( p2_u3430,n20128,n20129 );
   nand U19700 ( n20129,n19735,n19730 );
   nand U19701 ( n19730,n20130,n20131,n20132,n20133 );
   nand U19702 ( n20133,n20134,n20135 );
   nand U19703 ( n20134,n19759,n19777 );
   nand U19704 ( n20132,n20136,n19896 );
   not U19705 ( n19896,n19760 );
   nand U19706 ( n20131,n19893,n19629 );
   nand U19707 ( n20128,p2_reg0_reg_0_,n19743 );
   and U19708 ( n19732,n20141,n20142,n20143,n20144 );
   nand U19709 ( n20142,n20145,n20146,n20147 );
   or U19710 ( n20147,n20148,n20149 );
   nand U19711 ( p2_u3417,n20150,n20151 );
   nand U19712 ( n20151,p2_d_reg_1_,n20152 );
   nand U19713 ( n20150,n20153,n20154 );
   nand U19714 ( p2_u3416,n20155,n20156 );
   nand U19715 ( n20156,p2_d_reg_0_,n20152 );
   nand U19716 ( n20155,n20153,n20157 );
   nor U19717 ( p2_u3328,n20158,n20159 );
   nor U19718 ( n20159,n20160,n20161 );
   nor U19719 ( n20158,n20162,n20161,n20163,n20164 );
   nor U19720 ( n20164,n20165,n20166 );
   and U19721 ( n20163,n20165,n20167,n20168 );
   nand U19722 ( n20165,n20169,n20170,n20171,n20172 );
   nor U19723 ( n20172,n20173,n20174,n20175,n20176 );
   nand U19724 ( n20176,n20177,n20178,n20179,n20180 );
   nand U19725 ( n20175,n20181,n20182,n20183,n20184 );
   nand U19726 ( n20174,n20185,n20186,n20187,n20188 );
   nand U19727 ( n20173,n20189,n20190,n20191,n20192 );
   nor U19728 ( n20171,n20193,n20194,n20195,n20196 );
   nand U19729 ( n20194,n20197,n20198 );
   nand U19730 ( n20193,n20199,n20200,n20201,n20202 );
   nor U19731 ( n20170,n20203,n20204,n20205,n20206 );
   nor U19732 ( n20169,n20207,n20208,n20209,n20210 );
   xor U19733 ( n20208,n19740,n19539 );
   xor U19734 ( n20207,n20211,n20212 );
   and U19735 ( n20161,n20213,n20214,p2_b_reg );
   or U19736 ( n20214,n20215,n20216,n20217 );
   nand U19737 ( n20213,n20160,n20138 );
   not U19738 ( n20160,n20218 );
   nand U19739 ( n20162,n20219,n20220 );
   nand U19740 ( n20220,n20221,n20222 );
   nand U19741 ( n20221,n20223,n20224 );
   nand U19742 ( n20224,n20168,n20137 );
   nand U19743 ( n20219,n20225,n20226 );
   nand U19744 ( n20226,n20146,n20227 );
   nand U19745 ( n20227,n20228,n20229 );
   nand U19746 ( n20229,n20139,n20230 );
   nand U19747 ( n20230,n20137,n20138 );
   not U19748 ( n20225,n20222 );
   nand U19749 ( n20222,n20231,n20232,n20233,n20234 );
   nor U19750 ( n20234,n20235,n20236,n20237,n20238 );
   nor U19751 ( n20238,n20239,n20240 );
   not U19752 ( n20240,n20241 );
   nor U19753 ( n20239,n20242,n20243 );
   nor U19754 ( n20243,n20244,n20245 );
   nor U19755 ( n20244,n20246,n20247,n20248 );
   nor U19756 ( n20248,n20249,n20250,n20251 );
   not U19757 ( n20250,n20252 );
   nor U19758 ( n20247,n20253,n20254,n20255 );
   nor U19759 ( n20246,n20256,n20257 );
   nor U19760 ( n20242,n20258,n20259 );
   nor U19761 ( n20259,n20260,n20261 );
   nor U19762 ( n20261,n20262,n20263 );
   nor U19763 ( n20260,n20264,n20265 );
   nor U19764 ( n20265,n20266,n20267 );
   nor U19765 ( n20267,n20268,n20269 );
   nor U19766 ( n20266,n20270,n20271,n20272 );
   not U19767 ( n20271,n20273 );
   not U19768 ( n20264,n20274 );
   not U19769 ( n20258,n20275 );
   nor U19770 ( n20237,n20276,n20277,n20278 );
   nor U19771 ( n20236,n20279,n20280 );
   nor U19772 ( n20279,n20281,n20282 );
   nor U19773 ( n20282,n20283,n20284 );
   nor U19774 ( n20281,n20285,n20245,n20286,n20253 );
   nand U19775 ( n20253,n20287,n20252 );
   nand U19776 ( n20252,n20256,n20257 );
   nand U19777 ( n20257,n20288,n20289 );
   nand U19778 ( n20289,n20100,n20290 );
   nand U19779 ( n20288,n20291,n19623 );
   and U19780 ( n20256,n20292,n20293 );
   nand U19781 ( n20293,n20294,n19623 );
   nand U19782 ( n20292,n20291,n20100 );
   nand U19783 ( n20287,n20251,n20249 );
   nand U19784 ( n20249,n20295,n20296 );
   nand U19785 ( n20296,n20290,n20297 );
   nand U19786 ( n20295,n20291,n19626 );
   and U19787 ( n20251,n20298,n20299 );
   nand U19788 ( n20299,n20294,n19626 );
   nand U19789 ( n20298,n20291,n20297 );
   nand U19790 ( n20245,n20300,n20275,n20274,n20273 );
   nand U19791 ( n20273,n20268,n20269 );
   nand U19792 ( n20269,n20301,n20302 );
   nand U19793 ( n20302,n20072,n20290 );
   nand U19794 ( n20301,n20291,n19617 );
   and U19795 ( n20268,n20303,n20304 );
   nand U19796 ( n20304,n20294,n19617 );
   nand U19797 ( n20303,n20291,n20072 );
   nand U19798 ( n20274,n20262,n20263 );
   nand U19799 ( n20263,n20305,n20306 );
   nand U19800 ( n20306,n20290,n20061 );
   nand U19801 ( n20305,n20291,n19614 );
   and U19802 ( n20262,n20307,n20308 );
   nand U19803 ( n20308,n20294,n19614 );
   nand U19804 ( n20307,n20291,n20061 );
   nand U19805 ( n20275,n20309,n20310,n20311 );
   not U19806 ( n20311,n20312 );
   nand U19807 ( n20310,n20313,n20314 );
   nand U19808 ( n20309,n20315,n20060 );
   nand U19809 ( n20300,n20272,n20270 );
   nand U19810 ( n20270,n20316,n20317 );
   nand U19811 ( n20317,n20318,n20290 );
   nand U19812 ( n20316,n20291,n19620 );
   and U19813 ( n20272,n20319,n20320 );
   nand U19814 ( n20320,n20294,n19620 );
   nand U19815 ( n20319,n20291,n20318 );
   nand U19816 ( n20285,n20321,n20322,n20323,n20324 );
   nand U19817 ( n20324,n20325,n20326 );
   nand U19818 ( n20322,n20327,n20328 );
   or U19819 ( n20328,n20326,n20325 );
   and U19820 ( n20325,n20329,n20330 );
   nand U19821 ( n20330,n20294,n19632 );
   nand U19822 ( n20329,n20291,n20135 );
   nand U19823 ( n20326,n20331,n20332 );
   nand U19824 ( n20332,n20148,n20137 );
   not U19825 ( n20331,n20333 );
   nand U19826 ( n20327,n20334,n20335 );
   nand U19827 ( n20335,n20290,n20135 );
   nand U19828 ( n20334,n20291,n19632 );
   nand U19829 ( n20321,n20254,n20255 );
   nand U19830 ( n20255,n20336,n20337 );
   nand U19831 ( n20337,n20290,n20338 );
   nand U19832 ( n20336,n20291,n19629 );
   and U19833 ( n20254,n20339,n20340 );
   nand U19834 ( n20340,n20294,n19629 );
   nand U19835 ( n20339,n20291,n20338 );
   nand U19836 ( n20235,n20341,n20342,n20343 );
   nand U19837 ( n20343,n20241,n20344,n20313,n20312 );
   nand U19838 ( n20312,n20345,n20346 );
   nand U19839 ( n20346,n20294,n19611 );
   nand U19840 ( n20345,n20291,n20049 );
   nand U19841 ( n20313,n20049,n20290 );
   nand U19842 ( n20344,n20291,n19611 );
   nor U19843 ( n20241,n20286,n20278 );
   nand U19844 ( n20286,n20347,n20348,n20349,n20350 );
   nor U19845 ( n20350,n20351,n20352 );
   nand U19846 ( n20349,n20353,n20354 );
   nand U19847 ( n20342,n20355,n20356,n20357,n20358 );
   nand U19848 ( n20356,n20291,n19596 );
   nand U19849 ( n20341,n20359,n20360,n20361,n20362 );
   not U19850 ( n20360,n20278 );
   nor U19851 ( n20233,n20363,n20364,n20365 );
   nor U19852 ( n20365,n20366,n20367 );
   not U19853 ( n20367,n20355 );
   nor U19854 ( n20355,n20351,n20278 );
   nand U19855 ( n20278,n20368,n20323 );
   nand U19856 ( n20323,n20283,n20284 );
   nand U19857 ( n20284,n20369,n20370 );
   nand U19858 ( n20370,n20290,n20371 );
   nand U19859 ( n20369,n20291,n19587 );
   and U19860 ( n20283,n20372,n20373 );
   nand U19861 ( n20373,n20294,n19587 );
   nand U19862 ( n20372,n20291,n20371 );
   not U19863 ( n20368,n20280 );
   nand U19864 ( n20280,n20374,n20375,n20376,n20377 );
   nor U19865 ( n20377,n20378,n20379 );
   or U19866 ( n20374,n20380,n20381 );
   nand U19867 ( n20351,n20361,n20382 );
   or U19868 ( n20382,n20362,n20359 );
   and U19869 ( n20359,n20383,n20384 );
   nand U19870 ( n20384,n19973,n20290 );
   nand U19871 ( n20383,n20291,n19593 );
   nand U19872 ( n20362,n20385,n20386 );
   nand U19873 ( n20386,n20294,n19593 );
   nand U19874 ( n20385,n20291,n19973 );
   nand U19875 ( n20361,n20277,n20276 );
   nand U19876 ( n20276,n20387,n20388 );
   nand U19877 ( n20388,n20290,n20389 );
   nand U19878 ( n20387,n20291,n19590 );
   and U19879 ( n20277,n20390,n20391 );
   nand U19880 ( n20391,n20294,n19590 );
   nand U19881 ( n20390,n20291,n20389 );
   nor U19882 ( n20366,n20392,n20393 );
   nor U19883 ( n20393,n20394,n20352 );
   nand U19884 ( n20352,n20395,n20396 );
   nand U19885 ( n20396,n20397,n20398 );
   nor U19886 ( n20394,n20399,n20400 );
   nor U19887 ( n20400,n20401,n20402 );
   nor U19888 ( n20399,n20403,n20404 );
   nor U19889 ( n20404,n20405,n20406 );
   nor U19890 ( n20406,n20407,n20408 );
   nor U19891 ( n20405,n20354,n20409,n20353 );
   and U19892 ( n20353,n20410,n20411 );
   nand U19893 ( n20411,n20294,n19608 );
   nand U19894 ( n20410,n20291,n20038 );
   not U19895 ( n20409,n20347 );
   nand U19896 ( n20347,n20407,n20408 );
   nand U19897 ( n20408,n20412,n20413 );
   nand U19898 ( n20413,n20414,n20290 );
   nand U19899 ( n20412,n20291,n19605 );
   and U19900 ( n20407,n20415,n20416 );
   nand U19901 ( n20416,n20294,n19605 );
   nand U19902 ( n20415,n20291,n20414 );
   nand U19903 ( n20354,n20417,n20418 );
   nand U19904 ( n20418,n20038,n20290 );
   nand U19905 ( n20417,n20291,n19608 );
   not U19906 ( n20403,n20348 );
   nand U19907 ( n20348,n20401,n20402 );
   nand U19908 ( n20402,n20419,n20420 );
   nand U19909 ( n20420,n20290,n20011 );
   nand U19910 ( n20419,n20291,n19602 );
   and U19911 ( n20401,n20421,n20422 );
   nand U19912 ( n20422,n20294,n19602 );
   nand U19913 ( n20421,n20291,n20011 );
   nor U19914 ( n20392,n20398,n20397,n20423 );
   not U19915 ( n20423,n20395 );
   nand U19916 ( n20395,n20424,n20425,n20426 );
   not U19917 ( n20426,n20358 );
   nand U19918 ( n20358,n20427,n20428 );
   nand U19919 ( n20428,n20294,n19596 );
   nand U19920 ( n20427,n20291,n20429 );
   nand U19921 ( n20425,n20357,n20314 );
   nand U19922 ( n20357,n20429,n20290 );
   nand U19923 ( n20424,n20315,n19999 );
   and U19924 ( n20397,n20430,n20431 );
   nand U19925 ( n20431,n20294,n19599 );
   nand U19926 ( n20430,n20291,n20000 );
   nand U19927 ( n20398,n20432,n20433 );
   nand U19928 ( n20433,n20000,n20290 );
   nand U19929 ( n20432,n20291,n19599 );
   nor U19930 ( n20364,n20434,n20435 );
   nor U19931 ( n20435,n20436,n20437 );
   nor U19932 ( n20437,n20438,n20439 );
   nor U19933 ( n20436,n20440,n20441 );
   nor U19934 ( n20441,n20442,n20443 );
   nor U19935 ( n20443,n20444,n20445 );
   nor U19936 ( n20442,n20446,n20379 );
   nor U19937 ( n20446,n20447,n20448,n20449 );
   nor U19938 ( n20449,n20450,n20451 );
   nor U19939 ( n20448,n20452,n20453,n20454 );
   not U19940 ( n20453,n20455 );
   nor U19941 ( n20447,n20456,n20457 );
   not U19942 ( n20434,n20458 );
   nor U19943 ( n20363,n20459,n20460,n20461 );
   nor U19944 ( n20461,n20462,n20463,n20464 );
   nor U19945 ( n20464,n20465,n20466 );
   nor U19946 ( n20465,n20467,n20468 );
   nor U19947 ( n20468,n20469,n20470 );
   nor U19948 ( n20467,n20471,n20472,n20473 );
   not U19949 ( n20472,n20474 );
   nor U19950 ( n20463,n20475,n20476 );
   nor U19951 ( n20476,n20477,n20478 );
   nor U19952 ( n20478,n20479,n20480 );
   nor U19953 ( n20477,n20481,n20482,n20483 );
   not U19954 ( n20483,n20484 );
   not U19955 ( n20475,n20485 );
   nor U19956 ( n20462,n20486,n20487 );
   nor U19957 ( n20460,n20488,n20489 );
   not U19958 ( n20459,n20490 );
   nand U19959 ( n20232,n20490,n20491 );
   nand U19960 ( n20491,n20492,n20493,n20494 );
   nand U19961 ( n20494,n20488,n20489 );
   nand U19962 ( n20493,n20376,n20380,n20381 );
   and U19963 ( n20381,n20495,n20496 );
   nand U19964 ( n20496,n19934,n20290 );
   nand U19965 ( n20495,n20291,n19584 );
   nand U19966 ( n20380,n20497,n20498 );
   nand U19967 ( n20498,n20294,n19584 );
   nand U19968 ( n20497,n20291,n19934 );
   and U19969 ( n20376,n20499,n20500,n20501,n20502 );
   or U19970 ( n20500,n20503,n20504 );
   nand U19971 ( n20492,n20499,n20505 );
   nand U19972 ( n20505,n20506,n20507 );
   nand U19973 ( n20507,n20508,n20502 );
   nand U19974 ( n20502,n20509,n20510 );
   nand U19975 ( n20508,n20511,n20512 );
   nand U19976 ( n20512,n20501,n20503,n20504 );
   and U19977 ( n20504,n20513,n20514 );
   nand U19978 ( n20514,n19923,n20290 );
   nand U19979 ( n20513,n20291,n19581 );
   nand U19980 ( n20503,n20515,n20516,n20517 );
   nand U19981 ( n20517,n20518,n19581 );
   nand U19982 ( n20516,n20519,n19581 );
   nand U19983 ( n20515,n20291,n19923 );
   nand U19984 ( n20501,n20520,n20521 );
   or U19985 ( n20511,n20521,n20520 );
   and U19986 ( n20520,n20522,n20523,n20524 );
   nand U19987 ( n20524,n20518,n19578 );
   nand U19988 ( n20523,n20519,n19578 );
   nand U19989 ( n20522,n20291,n20525 );
   nand U19990 ( n20521,n20526,n20527 );
   nand U19991 ( n20527,n20525,n20290 );
   nand U19992 ( n20526,n20291,n19578 );
   or U19993 ( n20506,n20510,n20509 );
   and U19994 ( n20509,n20528,n20529 );
   nand U19995 ( n20529,n20294,n19575 );
   nand U19996 ( n20528,n20291,n20530 );
   nand U19997 ( n20510,n20531,n20532 );
   nand U19998 ( n20532,n20530,n20290 );
   nand U19999 ( n20531,n20291,n19575 );
   and U20000 ( n20499,n20533,n20534,n20535,n20474 );
   nand U20001 ( n20474,n20469,n20470 );
   nand U20002 ( n20470,n20536,n20537 );
   nand U20003 ( n20537,n19872,n20290 );
   nand U20004 ( n20536,n20291,n19569 );
   and U20005 ( n20469,n20538,n20539 );
   nand U20006 ( n20539,n20294,n19569 );
   nand U20007 ( n20538,n20291,n19872 );
   nand U20008 ( n20535,n20473,n20471 );
   nand U20009 ( n20471,n20540,n20541 );
   nand U20010 ( n20541,n19883,n20290 );
   nand U20011 ( n20540,n20291,n19572 );
   and U20012 ( n20473,n20542,n20543 );
   nand U20013 ( n20543,n20294,n19572 );
   nand U20014 ( n20542,n20291,n19883 );
   or U20015 ( n20534,n20489,n20488 );
   and U20016 ( n20488,n20544,n20545 );
   nand U20017 ( n20545,n20546,n20290 );
   nand U20018 ( n20544,n20291,n19557 );
   nand U20019 ( n20489,n20547,n20548 );
   nand U20020 ( n20548,n20294,n19557 );
   nand U20021 ( n20547,n20291,n20546 );
   not U20022 ( n20533,n20466 );
   nand U20023 ( n20466,n20549,n20485,n20484 );
   nand U20024 ( n20484,n20479,n20480 );
   nand U20025 ( n20480,n20550,n20551 );
   nand U20026 ( n20551,n19847,n20290 );
   nand U20027 ( n20550,n20291,n19563 );
   and U20028 ( n20479,n20552,n20553,n20554 );
   nand U20029 ( n20554,n20518,n19563 );
   nand U20030 ( n20553,n20519,n19563 );
   nand U20031 ( n20552,n20291,n19847 );
   nand U20032 ( n20485,n20486,n20487 );
   nand U20033 ( n20487,n20555,n20556 );
   nand U20034 ( n20556,n20557,n20290 );
   nand U20035 ( n20555,n20291,n19560 );
   and U20036 ( n20486,n20558,n20559 );
   nand U20037 ( n20559,n20294,n19560 );
   nand U20038 ( n20558,n20291,n20557 );
   nand U20039 ( n20549,n20482,n20481 );
   nand U20040 ( n20481,n20560,n20561 );
   nand U20041 ( n20561,n20562,n20290 );
   nand U20042 ( n20560,n20291,n19566 );
   and U20043 ( n20482,n20563,n20564,n20565 );
   nand U20044 ( n20565,n20518,n19566 );
   not U20045 ( n20518,n20566 );
   nand U20046 ( n20564,n20519,n19566 );
   nand U20047 ( n20563,n20291,n20562 );
   nor U20048 ( n20490,n20378,n20440,n20379 );
   nand U20049 ( n20379,n20567,n20568 );
   nand U20050 ( n20568,n20444,n20445 );
   nand U20051 ( n20445,n20569,n20570 );
   nand U20052 ( n20570,n19762,n20290 );
   nand U20053 ( n20569,n20291,n19545 );
   and U20054 ( n20444,n20571,n20572 );
   nand U20055 ( n20572,n20294,n19545 );
   nand U20056 ( n20571,n20291,n19762 );
   nand U20057 ( n20567,n20456,n20457 );
   nand U20058 ( n20457,n20573,n20574 );
   nand U20059 ( n20574,n20575,n20290 );
   nand U20060 ( n20573,n20291,n19548 );
   and U20061 ( n20456,n20576,n20577 );
   nand U20062 ( n20577,n20294,n19548 );
   nand U20063 ( n20576,n20291,n20575 );
   not U20064 ( n20440,n20375 );
   nand U20065 ( n20375,n20438,n20439 );
   nand U20066 ( n20439,n20578,n20579 );
   nand U20067 ( n20579,n19748,n20290 );
   nand U20068 ( n20578,n20291,n19542 );
   and U20069 ( n20438,n20580,n20581 );
   nand U20070 ( n20581,n20519,n19542 );
   nand U20071 ( n20580,n20291,n19748 );
   nand U20072 ( n20378,n20458,n20455,n20582 );
   nand U20073 ( n20582,n20454,n20452 );
   nand U20074 ( n20452,n20583,n20584 );
   nand U20075 ( n20584,n19804,n20290 );
   nand U20076 ( n20583,n20291,n19554 );
   and U20077 ( n20454,n20585,n20586 );
   nand U20078 ( n20586,n20294,n19554 );
   nand U20079 ( n20585,n20291,n19804 );
   nand U20080 ( n20455,n20450,n20451 );
   nand U20081 ( n20451,n20587,n20588 );
   nand U20082 ( n20588,n19793,n20290 );
   nand U20083 ( n20587,n20291,n19551 );
   and U20084 ( n20450,n20589,n20590 );
   nand U20085 ( n20590,n20294,n19551 );
   nand U20086 ( n20566,n19542,n20592,n20593 );
   nand U20087 ( n20589,n20291,n19793 );
   nand U20088 ( n20458,n20594,n20595 );
   nand U20089 ( n20231,n20594,n20596 );
   nand U20090 ( n20594,n20596,n20595 );
   nand U20091 ( n20595,n20597,n20598 );
   nand U20092 ( n20598,n20519,n19539 );
   not U20093 ( n20519,n20591 );
   nand U20094 ( n20591,n20290,n20599 );
   nand U20095 ( n20599,n20600,n19542,n20593,n20601 );
   nor U20096 ( n20601,n20602,n20603,n20149 );
   nand U20097 ( n20597,n20291,n19740 );
   nand U20098 ( n20596,n20604,n20605 );
   nand U20099 ( n20605,n19740,n20290 );
   nor U20100 ( n20315,n20149,n20603,n20602,n20606 );
   or U20101 ( n20606,n20607,n20592 );
   nand U20102 ( n20592,n20608,n20145,n20609 );
   nand U20103 ( n20604,n20291,n19539 );
   nand U20104 ( p2_u3327,n20610,n20611,n20612 );
   nand U20105 ( n20612,n20613,p1_datao_reg_0_ );
   nand U20106 ( n20611,p2_ir_reg_0_,n20614 );
   or U20107 ( n20614,n20615,n20616 );
   nand U20108 ( n20610,n20617,n20618 );
   nand U20109 ( p2_u3326,n20619,n20620,n20621,n20622 );
   nand U20110 ( n20622,p2_ir_reg_1_,n20623 );
   nand U20111 ( n20623,n20624,n20625 );
   nand U20112 ( n20625,n20616,n20626 );
   nand U20113 ( n20621,n20616,p2_ir_reg_0_,n20627 );
   nand U20114 ( n20620,n20617,n20628 );
   nand U20115 ( n20619,n20613,p1_datao_reg_1_ );
   nand U20116 ( p2_u3325,n20629,n20630,n20631,n20632 );
   nand U20117 ( n20632,n20633,n20616 );
   not U20118 ( n20633,n20634 );
   nand U20119 ( n20631,n20617,n20635 );
   nand U20120 ( n20630,n20613,p1_datao_reg_2_ );
   nand U20121 ( n20629,n20615,p2_ir_reg_2_ );
   nand U20122 ( p2_u3324,n20636,n20637,n20638,n20639 );
   nand U20123 ( n20639,p2_ir_reg_3_,n20640 );
   nand U20124 ( n20640,n20624,n20641 );
   nand U20125 ( n20641,n20616,n20642 );
   nand U20126 ( n20638,n20616,n20643,n20644 );
   nand U20127 ( n20637,n20645,n20617 );
   nand U20128 ( n20636,n20613,p1_datao_reg_3_ );
   nand U20129 ( p2_u3323,n20646,n20647,n20648,n20649 );
   nand U20130 ( n20649,n20650,n20651,n20616 );
   nand U20131 ( n20648,n20652,n20617 );
   nand U20132 ( n20647,n20613,p1_datao_reg_4_ );
   nand U20133 ( n20646,n20615,p2_ir_reg_4_ );
   nand U20134 ( p2_u3322,n20653,n20654,n20655,n20656 );
   nand U20135 ( n20656,p2_ir_reg_5_,n20657 );
   nand U20136 ( n20657,n20624,n20658 );
   nand U20137 ( n20658,n20616,n20659 );
   nand U20138 ( n20655,n20616,n20651,n20660 );
   nand U20139 ( n20654,n20661,n20617 );
   nand U20140 ( n20653,n20613,p1_datao_reg_5_ );
   nand U20141 ( p2_u3321,n20662,n20663,n20664,n20665 );
   nand U20142 ( n20665,n20666,n20667,n20616 );
   nand U20143 ( n20664,n20617,n20668 );
   nand U20144 ( n20663,n20613,p1_datao_reg_6_ );
   nand U20145 ( n20662,n20615,p2_ir_reg_6_ );
   nand U20146 ( p2_u3320,n20669,n20670,n20671,n20672 );
   nand U20147 ( n20672,p2_ir_reg_7_,n20673 );
   nand U20148 ( n20673,n20624,n20674 );
   nand U20149 ( n20674,n20616,n20675 );
   nand U20150 ( n20671,n20616,n20667,n20676 );
   nand U20151 ( n20670,n20677,n20617 );
   nand U20152 ( n20669,n20613,p1_datao_reg_7_ );
   nand U20153 ( p2_u3319,n20678,n20679,n20680,n20681 );
   nand U20154 ( n20681,n20682,n20683,n20616 );
   nand U20155 ( n20680,n20684,n20617 );
   nand U20156 ( n20679,n20613,p1_datao_reg_8_ );
   nand U20157 ( n20678,n20615,p2_ir_reg_8_ );
   nand U20158 ( p2_u3318,n20685,n20686,n20687,n20688 );
   nand U20159 ( n20688,p2_ir_reg_9_,n20689 );
   nand U20160 ( n20689,n20624,n20690 );
   nand U20161 ( n20690,n20616,n20691 );
   nand U20162 ( n20687,n20616,n20683,n20692 );
   nand U20163 ( n20686,n20693,n20617 );
   nand U20164 ( n20685,n20613,p1_datao_reg_9_ );
   nand U20165 ( p2_u3317,n20694,n20695,n20696,n20697 );
   nand U20166 ( n20697,n20698,n20616 );
   not U20167 ( n20698,n20699 );
   nand U20168 ( n20696,n20617,n20700 );
   nand U20169 ( n20695,n20613,p1_datao_reg_10_ );
   nand U20170 ( n20694,n20615,p2_ir_reg_10_ );
   nand U20171 ( p2_u3316,n20701,n20702,n20703,n20704 );
   nand U20172 ( n20704,p2_ir_reg_11_,n20705 );
   nand U20173 ( n20705,n20624,n20706 );
   nand U20174 ( n20706,n20616,n20707 );
   nand U20175 ( n20703,n20616,n20708,n20709 );
   nand U20176 ( n20702,n20710,n20617 );
   nand U20177 ( n20701,n20613,p1_datao_reg_11_ );
   nand U20178 ( p2_u3315,n20711,n20712,n20713,n20714 );
   nand U20179 ( n20714,n20715,n20616 );
   not U20180 ( n20715,n20716 );
   nand U20181 ( n20713,n20717,n20617 );
   nand U20182 ( n20712,n20613,p1_datao_reg_12_ );
   nand U20183 ( n20711,n20615,p2_ir_reg_12_ );
   nand U20184 ( p2_u3314,n20718,n20719,n20720,n20721 );
   nand U20185 ( n20721,p2_ir_reg_13_,n20722 );
   nand U20186 ( n20722,n20624,n20723 );
   nand U20187 ( n20723,n20616,n20724 );
   nand U20188 ( n20720,n20616,n20725,n20726 );
   nand U20189 ( n20719,n20727,n20617 );
   nand U20190 ( n20718,n20613,p1_datao_reg_13_ );
   nand U20191 ( p2_u3313,n20728,n20729,n20730,n20731 );
   nand U20192 ( n20731,n20732,n20616 );
   not U20193 ( n20732,n20733 );
   nand U20194 ( n20730,n20617,n20734 );
   nand U20195 ( n20729,n20613,p1_datao_reg_14_ );
   nand U20196 ( n20728,n20615,p2_ir_reg_14_ );
   nand U20197 ( p2_u3312,n20735,n20736,n20737,n20738 );
   nand U20198 ( n20738,p2_ir_reg_15_,n20739 );
   nand U20199 ( n20739,n20624,n20740 );
   nand U20200 ( n20740,n20616,n20741 );
   nand U20201 ( n20737,n20616,n20742,n20743 );
   nand U20202 ( n20736,n20617,n20744 );
   nand U20203 ( n20735,n20613,p1_datao_reg_15_ );
   nand U20204 ( p2_u3311,n20745,n20746,n20747,n20748 );
   nand U20205 ( n20748,n20749,n20616 );
   not U20206 ( n20749,n20750 );
   nand U20207 ( n20747,n20751,n20617 );
   nand U20208 ( n20746,n20613,p1_datao_reg_16_ );
   nand U20209 ( n20745,n20615,p2_ir_reg_16_ );
   nand U20210 ( p2_u3310,n20752,n20753,n20754,n20755 );
   nand U20211 ( n20755,p2_ir_reg_17_,n20756 );
   nand U20212 ( n20756,n20624,n20757 );
   nand U20213 ( n20757,n20616,n20758 );
   nand U20214 ( n20754,n20616,n20759,n20760 );
   nand U20215 ( n20753,n20761,n20617 );
   nand U20216 ( n20752,n20613,p1_datao_reg_17_ );
   nand U20217 ( p2_u3309,n20762,n20763,n20764,n20765 );
   nand U20218 ( n20765,n20766,n20616 );
   not U20219 ( n20766,n20767 );
   nand U20220 ( n20764,n20768,n20617 );
   nand U20221 ( n20763,n20613,p1_datao_reg_18_ );
   nand U20222 ( n20762,n20615,p2_ir_reg_18_ );
   nand U20223 ( p2_u3308,n20769,n20770,n20771,n20772 );
   nand U20224 ( n20772,p2_ir_reg_19_,n20773 );
   nand U20225 ( n20773,n20624,n20774 );
   nand U20226 ( n20774,n20616,n20775 );
   nand U20227 ( n20771,n20616,n20776,n20777 );
   nand U20228 ( n20770,n20778,n20617 );
   nand U20229 ( n20769,n20613,p1_datao_reg_19_ );
   nand U20230 ( p2_u3307,n20779,n20780,n20781,n20782 );
   nand U20231 ( n20782,n20783,n20784,n20616 );
   nand U20232 ( n20781,n20785,n20617 );
   nand U20233 ( n20780,n20613,p1_datao_reg_20_ );
   nand U20234 ( n20779,n20615,p2_ir_reg_20_ );
   nand U20235 ( p2_u3306,n20786,n20787,n20788,n20789 );
   nand U20236 ( n20789,p2_ir_reg_21_,n20790 );
   nand U20237 ( n20790,n20624,n20791 );
   nand U20238 ( n20791,n20616,n20792 );
   nand U20239 ( n20788,n20616,n20784,n20793 );
   nand U20240 ( n20787,n20794,n20617 );
   nand U20241 ( n20786,n20613,p1_datao_reg_21_ );
   nand U20242 ( p2_u3305,n20795,n20796,n20797,n20798 );
   nand U20243 ( n20798,p2_ir_reg_22_,n20799 );
   nand U20244 ( n20799,n20624,n20800 );
   nand U20245 ( n20800,n20616,n20801 );
   nand U20246 ( n20797,n20616,n20802,n20803 );
   nand U20247 ( n20796,n20804,n20617 );
   nand U20248 ( n20795,n20613,p1_datao_reg_22_ );
   nand U20249 ( p2_u3304,n20805,n20806,n20807,n20808 );
   nand U20250 ( n20808,n20809,n20810,n20616 );
   nand U20251 ( n20807,n20811,n20617 );
   nand U20252 ( n20806,n20613,p1_datao_reg_23_ );
   nand U20253 ( n20805,n20615,p2_ir_reg_23_ );
   nand U20254 ( p2_u3303,n20812,n20813,n20814,n20815 );
   nand U20255 ( n20815,n20816,n20817,n20616 );
   nand U20256 ( n20814,n20818,n20617 );
   nand U20257 ( n20813,n20613,p1_datao_reg_24_ );
   nand U20258 ( n20812,n20615,p2_ir_reg_24_ );
   nand U20259 ( p2_u3302,n20819,n20820,n20821,n20822 );
   nand U20260 ( n20822,p2_ir_reg_25_,n20823 );
   nand U20261 ( n20823,n20624,n20824 );
   nand U20262 ( n20824,n20616,n20825 );
   nand U20263 ( n20821,n20616,n20817,n20826 );
   nand U20264 ( n20820,n20827,n20617 );
   nand U20265 ( n20819,n20613,p1_datao_reg_25_ );
   nand U20266 ( p2_u3301,n20828,n20829,n20830,n20831 );
   nand U20267 ( n20831,n20832,n20833,n20616 );
   nand U20268 ( n20830,n20834,n20617 );
   nand U20269 ( n20829,n20613,p1_datao_reg_26_ );
   nand U20270 ( n20828,n20615,p2_ir_reg_26_ );
   nand U20271 ( p2_u3300,n20835,n20836,n20837,n20838 );
   nand U20272 ( n20838,p2_ir_reg_27_,n20839 );
   nand U20273 ( n20839,n20624,n20840 );
   nand U20274 ( n20840,n20616,n20841 );
   nand U20275 ( n20837,n20616,n20833,n20842 );
   nand U20276 ( n20836,n20843,n20617 );
   nand U20277 ( n20835,n20613,p1_datao_reg_27_ );
   nand U20278 ( p2_u3299,n20844,n20845,n20846,n20847 );
   nand U20279 ( n20847,p2_ir_reg_28_,n20848 );
   nand U20280 ( n20848,n20624,n20849 );
   nand U20281 ( n20849,n20616,n20850 );
   nand U20282 ( n20846,n20616,n20851,n20852 );
   nand U20283 ( n20845,n20853,n20617 );
   nand U20284 ( n20844,n20613,p1_datao_reg_28_ );
   nand U20285 ( p2_u3298,n20854,n20855,n20856,n20857 );
   nand U20286 ( n20857,n20858,n20859,n20616 );
   nand U20287 ( n20856,n20860,n20617 );
   nand U20288 ( n20855,n20613,p1_datao_reg_29_ );
   nand U20289 ( n20854,n20615,p2_ir_reg_29_ );
   nand U20290 ( p2_u3297,n20861,n20862,n20863,n20864 );
   nand U20291 ( n20864,p2_ir_reg_30_,n20865 );
   nand U20292 ( n20865,n20624,n20866 );
   nand U20293 ( n20866,n20867,n20616 );
   nand U20294 ( n20863,n20616,n20859,n20868 );
   not U20295 ( n20859,n20867 );
   nand U20296 ( n20862,n20617,n20869 );
   nand U20297 ( n20861,n20613,p1_datao_reg_30_ );
   nand U20298 ( p2_u3296,n20870,n20871 );
   nand U20299 ( n20871,n20616,n20868,n20867 );
   nor U20300 ( n20867,n20872,p2_ir_reg_29_ );
   not U20301 ( n20615,n20624 );
   nand U20302 ( n20624,p2_state_reg,n20873 );
   nand U20303 ( n20870,n20874,p2_u3088 );
   nor U20304 ( p2_u3295,n20153,n20875 );
   nor U20305 ( p2_u3294,n20153,n20876 );
   nor U20306 ( p2_u3293,n20153,n20877 );
   nor U20307 ( p2_u3292,n20153,n20878 );
   nor U20308 ( p2_u3291,n20153,n20879 );
   nor U20309 ( p2_u3290,n20153,n20880 );
   nor U20310 ( p2_u3289,n20153,n20881 );
   nor U20311 ( p2_u3288,n20153,n20882 );
   and U20312 ( p2_u3287,n20152,p2_d_reg_10_ );
   and U20313 ( p2_u3286,n20152,p2_d_reg_11_ );
   and U20314 ( p2_u3285,n20152,p2_d_reg_12_ );
   nor U20315 ( p2_u3284,n20153,n20883 );
   nor U20316 ( p2_u3283,n20153,n20884 );
   nor U20317 ( p2_u3282,n20153,n20885 );
   nor U20318 ( p2_u3281,n20153,n20886 );
   and U20319 ( p2_u3280,n20152,p2_d_reg_17_ );
   and U20320 ( p2_u3279,n20152,p2_d_reg_18_ );
   and U20321 ( p2_u3278,n20152,p2_d_reg_19_ );
   and U20322 ( p2_u3277,n20152,p2_d_reg_20_ );
   and U20323 ( p2_u3276,n20152,p2_d_reg_21_ );
   and U20324 ( p2_u3275,n20152,p2_d_reg_22_ );
   and U20325 ( p2_u3274,n20152,p2_d_reg_23_ );
   and U20326 ( p2_u3273,n20152,p2_d_reg_24_ );
   nor U20327 ( p2_u3272,n20153,n20887 );
   nor U20328 ( p2_u3271,n20153,n20888 );
   nor U20329 ( p2_u3270,n20153,n20889 );
   nor U20330 ( p2_u3269,n20153,n20890 );
   nor U20331 ( p2_u3268,n20153,n20891 );
   nor U20332 ( p2_u3267,n20153,n20892 );
   nor U20333 ( p2_u3266,n20153,n20893 );
   nand U20334 ( n20152,n20141,n20894 );
   nand U20335 ( p2_u3265,n20895,n20896,n20897,n20898 );
   nor U20336 ( n20898,n20899,n20900,n20901 );
   nor U20337 ( n20901,n20130,n20902 );
   and U20338 ( n20130,n20903,n20904 );
   nand U20339 ( n20904,n20905,n19818 );
   nand U20340 ( n20905,n20906,n20907 );
   nand U20341 ( n20907,n20908,n19632 );
   nand U20342 ( n20903,n20136,n20909 );
   nor U20343 ( n20900,n20910,n20911 );
   and U20344 ( n20899,p2_reg3_reg_0_,n20912 );
   nand U20345 ( n20897,n20913,n19629 );
   nand U20346 ( n20896,n20914,n20135 );
   nand U20347 ( n20914,n20915,n20916 );
   nand U20348 ( n20895,n20917,n20136 );
   not U20349 ( n20136,n20189 );
   nand U20350 ( n20189,n20918,n20919 );
   nand U20351 ( n20918,n20122,n20908 );
   nand U20352 ( p2_u3264,n20920,n20921,n20922,n20923 );
   nor U20353 ( n20923,n20924,n20925,n20926,n20927 );
   nor U20354 ( n20927,n20910,n20928 );
   nor U20355 ( n20926,n20123,n20915 );
   and U20356 ( n20925,p2_reg3_reg_1_,n20912 );
   nor U20357 ( n20924,n20099,n20929 );
   nor U20358 ( n20922,n20930,n20931 );
   and U20359 ( n20931,n20125,n20932 );
   xor U20360 ( n20125,n20338,n20135 );
   and U20361 ( n20930,n20124,n20933 );
   xor U20362 ( n20124,n20934,n20195 );
   nand U20363 ( n20921,n20935,n19632 );
   nand U20364 ( n20920,n20126,n20936 );
   xor U20365 ( n20126,n20937,n20195 );
   nor U20366 ( n20195,n20938,n20939 );
   not U20367 ( n20937,n20919 );
   nand U20368 ( p2_u3263,n20940,n20941,n20942,n20943 );
   nor U20369 ( n20943,n20944,n20945,n20946,n20947 );
   nor U20370 ( n20947,n20083,n20929 );
   nor U20371 ( n20946,n20112,n20916 );
   nand U20372 ( n20112,n20948,n20949 );
   nand U20373 ( n20949,n20950,n20297 );
   nand U20374 ( n20950,n20123,n20908 );
   nor U20375 ( n20945,n20951,n20111 );
   nand U20376 ( n20111,n20952,n20953 );
   or U20377 ( n20953,n20197,n20954 );
   nand U20378 ( n20952,n20955,n20956,n20954 );
   nor U20379 ( n20954,n20957,n20938 );
   nor U20380 ( n20944,n20958,n20959 );
   nor U20381 ( n20942,n20960,n20961 );
   nor U20382 ( n20961,n20110,n20915 );
   and U20383 ( n20960,p2_reg3_reg_2_,n20912 );
   nand U20384 ( n20941,p2_reg2_reg_2_,n20902 );
   nand U20385 ( n20940,n20910,n20107 );
   nand U20386 ( n20107,n20962,n20963,n20964,n20965 );
   nand U20387 ( n20965,n20966,n20967 );
   nand U20388 ( n20964,n20966,n20607 );
   nand U20389 ( n20963,n20966,n20968 );
   nand U20390 ( n20962,n20966,n20969 );
   and U20391 ( n20966,n20970,n20971 );
   or U20392 ( n20971,n20197,n20972 );
   nand U20393 ( n20197,n20973,n20974 );
   nand U20394 ( n20970,n20955,n20956,n20972 );
   nand U20395 ( p2_u3262,n20975,n20976,n20977,n20978 );
   nor U20396 ( n20978,n20979,n20980,n20981,n20982 );
   nor U20397 ( n20982,n20983,n20929 );
   nor U20398 ( n20981,n20951,n20097 );
   xor U20399 ( n20097,n20984,n20985 );
   nand U20400 ( n20985,n20986,n20987 );
   nand U20401 ( n20987,n20957,n20973 );
   nor U20402 ( n20980,n20099,n20959 );
   nor U20403 ( n20979,n20098,n20916 );
   xor U20404 ( n20098,n20100,n20988 );
   nor U20405 ( n20977,n20989,n20990 );
   nor U20406 ( n20990,n20092,n20902 );
   and U20407 ( n20092,n20991,n20992 );
   nand U20408 ( n20992,n20967,n20993 );
   nand U20409 ( n20991,n20994,n20993 );
   nand U20410 ( n20993,n20995,n20996 );
   nand U20411 ( n20996,n20997,n20956 );
   and U20412 ( n20997,n20206,n20998 );
   nand U20413 ( n20998,n20999,n20955 );
   nand U20414 ( n20995,n21000,n20984 );
   not U20415 ( n20984,n20206 );
   xor U20416 ( n20206,n20100,n19623 );
   nor U20417 ( n20989,n20910,n21001 );
   nand U20418 ( n20976,n20912,n21002 );
   nand U20419 ( n20975,n21003,n20100 );
   nand U20420 ( p2_u3261,n21004,n21005,n21006,n21007 );
   nor U20421 ( n21007,n21008,n21009,n21010,n21011 );
   and U20422 ( n21011,n20902,p2_reg2_reg_4_ );
   nor U20423 ( n21010,n20084,n20915 );
   nor U20424 ( n21009,n20082,n20929 );
   nor U20425 ( n21008,n20085,n20916 );
   nand U20426 ( n20085,n21012,n21013 );
   nand U20427 ( n21013,n20318,n21014 );
   nand U20428 ( n21014,n20988,n21015 );
   nor U20429 ( n21006,n21016,n21017 );
   and U20430 ( n21017,n20936,n20086 );
   xor U20431 ( n20086,n20205,n21018 );
   nor U20432 ( n21016,n20083,n20959 );
   nand U20433 ( n21005,n20933,n20087 );
   xor U20434 ( n20087,n21019,n21020 );
   not U20435 ( n21019,n20205 );
   xor U20436 ( n20205,n20318,n19620 );
   nand U20437 ( n21004,n20912,n21021 );
   nand U20438 ( p2_u3260,n21022,n21023,n21024,n21025 );
   nor U20439 ( n21025,n21026,n21027,n21028,n21029 );
   nor U20440 ( n21029,n21030,n20915 );
   and U20441 ( n21028,n21031,n20912 );
   nor U20442 ( n21027,n20064,n20902 );
   and U20443 ( n20064,n21032,n21033,n21034,n21035 );
   nor U20444 ( n21035,n21036,n21037,n21038,n21039 );
   nor U20445 ( n21039,n20983,n19776 );
   nor U20446 ( n21038,n21040,n21041 );
   nor U20447 ( n21037,n21042,n21041 );
   nor U20448 ( n21036,n20070,n21043 );
   not U20449 ( n20070,n21044 );
   nor U20450 ( n21034,n21045,n21046 );
   nor U20451 ( n21046,n20609,n21041 );
   nor U20452 ( n21045,n20600,n21041 );
   nand U20453 ( n21041,n21047,n21048 );
   nand U20454 ( n21048,n21049,n21050,n21051 );
   or U20455 ( n21047,n20198,n21051 );
   nand U20456 ( n21033,n21052,n21044 );
   nand U20457 ( n21032,n21053,n21044 );
   nor U20458 ( n21026,n20910,n21054 );
   nand U20459 ( n21024,n20913,n19614 );
   or U20460 ( n21023,n20916,n20071 );
   xor U20461 ( n20071,n21030,n21012 );
   nand U20462 ( n21022,n20917,n21044 );
   xor U20463 ( n21044,n20198,n21055 );
   nand U20464 ( n20198,n21056,n21057 );
   nand U20465 ( p2_u3259,n21058,n21059,n21060,n21061 );
   nor U20466 ( n21061,n21062,n21063,n21064,n21065 );
   nor U20467 ( n21065,n21066,n20915 );
   nor U20468 ( n21064,n21067,n21068 );
   nor U20469 ( n21063,n20052,n20902 );
   and U20470 ( n20052,n21069,n21070,n21071,n21072 );
   nor U20471 ( n21072,n21073,n21074,n21075,n21076 );
   nor U20472 ( n21076,n21077,n21040 );
   nor U20473 ( n21075,n20059,n21078 );
   nor U20474 ( n21074,n21077,n21042 );
   nor U20475 ( n21073,n20059,n20608 );
   nand U20476 ( n21071,n20602,n21079 );
   nand U20477 ( n21070,n21080,n21081 );
   not U20478 ( n21080,n21077 );
   nor U20479 ( n21077,n21082,n21083 );
   nand U20480 ( n21083,n21084,n21085 );
   nand U20481 ( n21085,n21086,n21050,n20199 );
   or U20482 ( n21084,n21086,n20199 );
   nor U20483 ( n21082,n20199,n21050 );
   nand U20484 ( n21069,n19960,n19617 );
   and U20485 ( n21062,n20902,p2_reg2_reg_6_ );
   nand U20486 ( n21060,n20913,n19611 );
   nand U20487 ( n21059,n20917,n21079 );
   not U20488 ( n21079,n20059 );
   xor U20489 ( n20059,n20199,n21087 );
   nand U20490 ( n20199,n21088,n21089 );
   or U20491 ( n21058,n20916,n20058 );
   nand U20492 ( n20058,n21090,n21091 );
   nand U20493 ( n21091,n21092,n20061 );
   nand U20494 ( n21092,n21093,n21030 );
   nand U20495 ( p2_u3258,n21094,n21095,n21096,n21097 );
   nor U20496 ( n21097,n21098,n21099,n21100,n21101 );
   nor U20497 ( n21101,n21102,n20915 );
   and U20498 ( n21100,n21103,n20912 );
   nor U20499 ( n21099,n20041,n20902 );
   and U20500 ( n20041,n21104,n21105,n21106,n21107 );
   nor U20501 ( n21107,n21108,n21109,n21110,n21111 );
   nor U20502 ( n21111,n21040,n21112 );
   nor U20503 ( n21110,n20609,n21112 );
   nor U20504 ( n21109,n21113,n19776 );
   nor U20505 ( n21108,n20600,n21112 );
   nor U20506 ( n21106,n21114,n21115 );
   nor U20507 ( n21115,n20608,n20047 );
   nor U20508 ( n21114,n21042,n21112 );
   nand U20509 ( n21112,n21116,n21117 );
   nand U20510 ( n21117,n21118,n21119 );
   nand U20511 ( n21116,n21120,n21121 );
   nand U20512 ( n21105,n21122,n20602 );
   nand U20513 ( n21104,n21122,n21053 );
   nor U20514 ( n21098,n20910,n21123 );
   nand U20515 ( n21096,n20913,n19608 );
   or U20516 ( n21095,n20916,n20048 );
   xor U20517 ( n20048,n21102,n21090 );
   nand U20518 ( n21094,n20917,n21122 );
   not U20519 ( n21122,n20047 );
   nand U20520 ( n20047,n21124,n21125 );
   nand U20521 ( n21125,n21126,n21088,n20200 );
   nand U20522 ( n21124,n21127,n21089,n21118 );
   not U20523 ( n21118,n20200 );
   nand U20524 ( n20200,n21128,n21129 );
   nand U20525 ( n21127,n21130,n21088 );
   nand U20526 ( p2_u3257,n21131,n21132,n21133,n21134 );
   nor U20527 ( n21134,n21135,n21136,n21137,n21138 );
   nor U20528 ( n21138,n21139,n20915 );
   nor U20529 ( n21137,n21140,n21068 );
   nor U20530 ( n21136,n20029,n20902 );
   and U20531 ( n20029,n21141,n21142,n21143,n21144 );
   nor U20532 ( n21144,n21145,n21146,n21147,n21148 );
   nor U20533 ( n21148,n21149,n21040 );
   xor U20534 ( n21149,n21150,n20201 );
   nor U20535 ( n21147,n21151,n21042 );
   nor U20536 ( n21151,n21152,n21153 );
   not U20537 ( n21153,n21154 );
   nor U20538 ( n21152,n21150,n20201 );
   nor U20539 ( n21146,n20036,n20608 );
   nor U20540 ( n21145,n20060,n19776 );
   nand U20541 ( n21143,n21053,n21155 );
   nand U20542 ( n21142,n21081,n21156 );
   nand U20543 ( n21156,n21157,n21154 );
   nand U20544 ( n21154,n21150,n20201 );
   nand U20545 ( n21157,n21158,n21159 );
   not U20546 ( n21158,n20201 );
   nand U20547 ( n21081,n20600,n20609 );
   nand U20548 ( n21141,n20602,n21155 );
   nor U20549 ( n21135,n20910,n21160 );
   nand U20550 ( n21133,n20913,n19605 );
   or U20551 ( n21132,n20916,n20035 );
   nand U20552 ( n20035,n21161,n21162 );
   nand U20553 ( n21162,n20038,n21163 );
   nand U20554 ( n21163,n21164,n21102 );
   nand U20555 ( n21131,n20917,n21155 );
   not U20556 ( n21155,n20036 );
   xor U20557 ( n20036,n21165,n20201 );
   nand U20558 ( n20201,n21166,n21167 );
   nand U20559 ( p2_u3256,n21168,n21169,n21170,n21171 );
   nor U20560 ( n21171,n21172,n21173,n21174,n21175 );
   and U20561 ( n21175,n20902,p2_reg2_reg_9_ );
   nor U20562 ( n21174,n20023,n20915 );
   and U20563 ( n21173,n21176,n20912 );
   nor U20564 ( n21172,n20021,n20929 );
   nor U20565 ( n21170,n21177,n21178 );
   nor U20566 ( n21178,n20951,n20026 );
   xor U20567 ( n20026,n20190,n21179 );
   nor U20568 ( n21177,n20022,n20959 );
   nand U20569 ( n21169,n20933,n20024 );
   nand U20570 ( n20024,n21180,n21181 );
   nand U20571 ( n21181,n21182,n20190 );
   nand U20572 ( n20190,n21183,n21184 );
   not U20573 ( n21182,n21185 );
   nand U20574 ( n21180,n21186,n21185 );
   nand U20575 ( n21186,n21187,n21188 );
   nand U20576 ( n21168,n20932,n20025 );
   xor U20577 ( n20025,n20414,n21161 );
   nand U20578 ( p2_u3255,n21189,n21190,n21191,n21192 );
   nor U20579 ( n21192,n21193,n21194,n21195,n21196 );
   nor U20580 ( n21196,n21197,n20915 );
   nor U20581 ( n21195,n21198,n21068 );
   nor U20582 ( n21194,n20003,n20902 );
   and U20583 ( n20003,n21199,n21200,n21201,n21202 );
   nor U20584 ( n21202,n21203,n21204,n21205,n21206 );
   nor U20585 ( n21206,n20600,n21207 );
   nor U20586 ( n21205,n21078,n20010 );
   nor U20587 ( n21204,n21043,n20010 );
   nor U20588 ( n21203,n20608,n20010 );
   nand U20589 ( n21201,n21208,n20968 );
   nand U20590 ( n21200,n21208,n21209 );
   nand U20591 ( n21209,n21040,n21042 );
   not U20592 ( n21208,n21207 );
   nand U20593 ( n21207,n21210,n21211 );
   nand U20594 ( n21211,n21212,n21213,n21214 );
   nand U20595 ( n21210,n21215,n21216 );
   nand U20596 ( n21199,n19960,n19605 );
   nor U20597 ( n21193,n20910,n21217 );
   nand U20598 ( n21191,n20913,n19599 );
   or U20599 ( n21190,n20916,n20009 );
   nand U20600 ( n20009,n21218,n21219 );
   nand U20601 ( n21219,n21220,n20011 );
   nand U20602 ( n21220,n21221,n20023 );
   or U20603 ( n21189,n21222,n20010 );
   nand U20604 ( n20010,n21223,n21224 );
   nand U20605 ( n21224,n21225,n21183,n20202 );
   nand U20606 ( n21223,n21226,n21184,n21215 );
   not U20607 ( n21215,n20202 );
   nand U20608 ( n20202,n21227,n21228 );
   nand U20609 ( n21226,n21229,n21183 );
   not U20610 ( n21229,n21179 );
   nand U20611 ( p2_u3254,n21230,n21231,n21232,n21233 );
   nor U20612 ( n21233,n21234,n21235,n21236,n21237 );
   nor U20613 ( n21237,n21238,n20915 );
   nor U20614 ( n21236,n21239,n21068 );
   nor U20615 ( n21235,n19991,n20902 );
   and U20616 ( n19991,n21240,n21241 );
   nor U20617 ( n21241,n21242,n21243,n21244,n21245 );
   nor U20618 ( n21245,n21246,n21042 );
   nor U20619 ( n21244,n20608,n19997 );
   nor U20620 ( n21243,n20021,n19776 );
   nor U20621 ( n21242,n21246,n20609 );
   nor U20622 ( n21240,n21247,n21248,n21249,n21250 );
   nor U20623 ( n21250,n21246,n20600 );
   and U20624 ( n21246,n21251,n21252,n21253 );
   not U20625 ( n21253,n21254 );
   nand U20626 ( n21252,n21255,n21214 );
   nand U20627 ( n21251,n21216,n21256 );
   nor U20628 ( n21249,n21078,n19997 );
   nor U20629 ( n21248,n21043,n19997 );
   nor U20630 ( n21247,n21257,n21040 );
   nor U20631 ( n21257,n21254,n21258,n21259 );
   nor U20632 ( n21259,n21260,n21214 );
   and U20633 ( n21258,n21214,n21255 );
   not U20634 ( n21214,n21216 );
   nor U20635 ( n21216,n21261,n21262 );
   nand U20636 ( n21254,n21263,n21264 );
   nand U20637 ( n21264,n21265,n21255 );
   nor U20638 ( n21255,n20177,n21266 );
   not U20639 ( n21265,n21212 );
   nand U20640 ( n21263,n21266,n21256 );
   not U20641 ( n21256,n21260 );
   nand U20642 ( n21260,n21267,n21268 );
   not U20643 ( n21266,n21213 );
   nor U20644 ( n21234,n20910,n21269 );
   nand U20645 ( n21232,n20913,n19596 );
   or U20646 ( n21231,n20916,n19998 );
   xor U20647 ( n19998,n21238,n21218 );
   or U20648 ( n21230,n21222,n19997 );
   xor U20649 ( n19997,n20177,n21270 );
   or U20650 ( n20177,n21271,n21272 );
   nor U20651 ( n21272,n19599,n20000 );
   nand U20652 ( p2_u3253,n21273,n21274,n21275,n21276 );
   nor U20653 ( n21276,n21277,n21278,n21279,n21280 );
   and U20654 ( n21280,n20902,p2_reg2_reg_12_ );
   nor U20655 ( n21279,n19985,n20915 );
   nor U20656 ( n21278,n21281,n21068 );
   nor U20657 ( n21277,n19983,n20929 );
   nor U20658 ( n21275,n21282,n21283 );
   nor U20659 ( n21283,n19986,n20916 );
   nand U20660 ( n19986,n21284,n21285 );
   nand U20661 ( n21285,n20429,n21286 );
   nand U20662 ( n21286,n21287,n21238 );
   nor U20663 ( n21282,n20951,n19987 );
   xor U20664 ( n19987,n20178,n21288 );
   nand U20665 ( n21274,n20933,n19988 );
   xor U20666 ( n19988,n21289,n20178 );
   nand U20667 ( n20178,n21290,n21291 );
   nand U20668 ( n21273,n20935,n19599 );
   nand U20669 ( p2_u3252,n21292,n21293,n21294,n21295 );
   nor U20670 ( n21295,n21296,n21297,n21298,n21299 );
   nor U20671 ( n21299,n21300,n20915 );
   and U20672 ( n21298,n21301,n20912 );
   nor U20673 ( n21297,n19965,n20902 );
   and U20674 ( n19965,n21302,n21303,n21304,n21305 );
   nor U20675 ( n21305,n21306,n21307,n21308,n21309 );
   nor U20676 ( n21309,n21078,n19971 );
   nor U20677 ( n21308,n21043,n19971 );
   nor U20678 ( n21307,n20608,n19971 );
   nor U20679 ( n21306,n21040,n21310 );
   nor U20680 ( n21304,n21311,n21312 );
   nor U20681 ( n21312,n19999,n19776 );
   nor U20682 ( n21311,n20600,n21310 );
   not U20683 ( n21310,n21313 );
   nand U20684 ( n21303,n21313,n20968 );
   nand U20685 ( n21302,n21313,n20967 );
   xor U20686 ( n21313,n21314,n20179 );
   nor U20687 ( n21296,n20910,n21315 );
   nand U20688 ( n21294,n20913,n19590 );
   or U20689 ( n21293,n20916,n19972 );
   xor U20690 ( n19972,n21300,n21284 );
   or U20691 ( n21292,n21222,n19971 );
   nand U20692 ( n19971,n21316,n21317 );
   nand U20693 ( n21317,n21318,n21291,n20179 );
   nand U20694 ( n21318,n21290,n21288 );
   not U20695 ( n21288,n21319 );
   nand U20696 ( n21316,n21320,n21290,n21321 );
   not U20697 ( n21321,n20179 );
   nand U20698 ( n20179,n21322,n21323 );
   nand U20699 ( n21320,n21319,n21291 );
   nor U20700 ( n21319,n21324,n21271 );
   nand U20701 ( p2_u3251,n21325,n21326,n21327,n21328 );
   nor U20702 ( n21328,n21329,n21330,n21331,n21332 );
   nor U20703 ( n21332,n19959,n20929 );
   nor U20704 ( n21331,n19962,n20916 );
   nand U20705 ( n19962,n21333,n21334 );
   nand U20706 ( n21334,n21335,n20389 );
   nand U20707 ( n21335,n21336,n21300 );
   nor U20708 ( n21330,n20951,n19961 );
   xor U20709 ( n19961,n21337,n20210 );
   nor U20710 ( n21329,n19983,n20959 );
   nor U20711 ( n21327,n21338,n21339 );
   nor U20712 ( n21339,n19958,n20915 );
   nor U20713 ( n21338,n21340,n21068 );
   nand U20714 ( n21326,p2_reg2_reg_14_,n20902 );
   nand U20715 ( n21325,n20910,n19955 );
   nand U20716 ( n19955,n21341,n21342 );
   nand U20717 ( n21342,n21343,n21344,n20968 );
   nand U20718 ( n21343,n21345,n21346 );
   nand U20719 ( n21341,n21347,n21344,n21348 );
   nand U20720 ( n21344,n20210,n21349 );
   xor U20721 ( n20210,n19590,n20389 );
   nand U20722 ( n21347,n21350,n21346,n21351 );
   nand U20723 ( p2_u3250,n21352,n21353,n21354,n21355 );
   nor U20724 ( n21355,n21356,n21357,n21358,n21359 );
   nor U20725 ( n21359,n19944,n20929 );
   and U20726 ( n21358,n20936,n19947 );
   xor U20727 ( n19947,n21360,n20209 );
   nor U20728 ( n21357,n19945,n20959 );
   and U20729 ( n21356,n19948,n20932 );
   xor U20730 ( n19948,n20371,n21333 );
   nor U20731 ( n21354,n21361,n21362 );
   nor U20732 ( n21362,n20902,n19938 );
   nand U20733 ( n19938,n21363,n21364,n19818 );
   nand U20734 ( n21364,n21365,n21366 );
   nand U20735 ( n21363,n21367,n20209 );
   xor U20736 ( n20209,n19587,n20371 );
   nor U20737 ( n21361,n20910,n21368 );
   nand U20738 ( n21353,n20912,n21369 );
   nand U20739 ( n21352,n21003,n20371 );
   nand U20740 ( p2_u3249,n21370,n21371,n21372,n21373 );
   nor U20741 ( n21373,n21374,n21375,n21376,n21377 );
   nor U20742 ( n21377,n21378,n20915 );
   nor U20743 ( n21376,n21379,n21068 );
   nor U20744 ( n21375,n19926,n20902 );
   and U20745 ( n19926,n21380,n21381 );
   nor U20746 ( n21381,n21382,n21383,n21384,n21385 );
   nor U20747 ( n21385,n21042,n21386,n21387 );
   nor U20748 ( n21387,n21388,n21389 );
   nor U20749 ( n21389,n20191,n21390,n21391 );
   and U20750 ( n21391,n21366,n21367 );
   and U20751 ( n21386,n20191,n21365 );
   nor U20752 ( n21384,n21392,n21040 );
   nor U20753 ( n21383,n19933,n21078 );
   nor U20754 ( n21382,n21392,n20609 );
   nor U20755 ( n21380,n21393,n21394,n21395,n21396 );
   nor U20756 ( n21396,n19933,n21043 );
   nor U20757 ( n21395,n19933,n20608 );
   nor U20758 ( n21394,n21392,n20600 );
   and U20759 ( n21392,n21397,n21398,n21399,n21400 );
   nand U20760 ( n21400,n21401,n21365 );
   nor U20761 ( n21365,n21367,n21390 );
   nand U20762 ( n21399,n21367,n21388 );
   nor U20763 ( n21367,n21345,n21402 );
   nand U20764 ( n21398,n21390,n21388 );
   and U20765 ( n21388,n21403,n21404 );
   not U20766 ( n21390,n21405 );
   or U20767 ( n21397,n21366,n20191 );
   nor U20768 ( n21393,n19959,n19776 );
   and U20769 ( n21374,n20902,p2_reg2_reg_16_ );
   nand U20770 ( n21372,n20913,n19581 );
   or U20771 ( n21371,n20916,n19932 );
   nand U20772 ( n19932,n21406,n21407 );
   nand U20773 ( n21407,n19934,n21408 );
   nand U20774 ( n21408,n21409,n19946 );
   or U20775 ( n21370,n21222,n19933 );
   xor U20776 ( n19933,n21401,n21410 );
   not U20777 ( n21401,n20191 );
   nand U20778 ( n20191,n21411,n21412 );
   nand U20779 ( p2_u3248,n21413,n21414,n21415,n21416 );
   nor U20780 ( n21416,n21417,n21418,n21419,n21420 );
   nor U20781 ( n21420,n21421,n20915 );
   nor U20782 ( n21419,n21422,n21068 );
   nor U20783 ( n21418,n19914,n20902 );
   and U20784 ( n19914,n21423,n21424,n21425,n21426 );
   nor U20785 ( n21426,n21427,n21428,n21429,n21430 );
   nor U20786 ( n21430,n21078,n19920 );
   nor U20787 ( n21429,n21043,n19920 );
   nor U20788 ( n21428,n20608,n19920 );
   nor U20789 ( n21427,n21431,n21040 );
   nor U20790 ( n21425,n21432,n21433 );
   nor U20791 ( n21433,n19944,n19776 );
   nor U20792 ( n21432,n21431,n20600 );
   nand U20793 ( n21424,n20968,n21434 );
   nand U20794 ( n21423,n20967,n21434 );
   not U20795 ( n21434,n21431 );
   xor U20796 ( n21431,n21435,n21436 );
   nor U20797 ( n21417,n20910,n21437 );
   nand U20798 ( n21415,n20913,n19578 );
   or U20799 ( n21414,n20916,n19921 );
   xor U20800 ( n19921,n21421,n21406 );
   or U20801 ( n21413,n21222,n19920 );
   nand U20802 ( n19920,n21438,n21439 );
   nand U20803 ( n21439,n21440,n21411,n20180 );
   nand U20804 ( n21438,n21441,n21412,n21435 );
   not U20805 ( n21435,n20180 );
   nand U20806 ( n20180,n21442,n21443 );
   nand U20807 ( n21441,n21410,n21411 );
   nand U20808 ( p2_u3247,n21444,n21445,n21446,n21447 );
   nor U20809 ( n21447,n21448,n21449,n21450,n21451 );
   nor U20810 ( n21451,n20910,n21452 );
   nor U20811 ( n21450,n19908,n20915 );
   nor U20812 ( n21449,n21453,n21068 );
   nor U20813 ( n21448,n19906,n20929 );
   nor U20814 ( n21446,n21454,n21455 );
   nor U20815 ( n21455,n19909,n20916 );
   nand U20816 ( n19909,n21456,n21457 );
   nand U20817 ( n21457,n20525,n21458 );
   nand U20818 ( n21458,n21459,n21421 );
   nor U20819 ( n21454,n20951,n19910 );
   xor U20820 ( n19910,n20181,n21460 );
   not U20821 ( n20181,n21461 );
   nand U20822 ( n21445,n20933,n19911 );
   xor U20823 ( n19911,n21461,n21462 );
   nor U20824 ( n21461,n21463,n21464 );
   nor U20825 ( n21464,n19578,n20525 );
   nand U20826 ( n21444,n20935,n19581 );
   nand U20827 ( p2_u3246,n21465,n21466,n21467,n21468 );
   nor U20828 ( n21468,n21469,n21470,n21471,n21472 );
   nor U20829 ( n21472,n19892,n20915 );
   nor U20830 ( n21471,n21473,n21068 );
   and U20831 ( n21470,n19891,n20910 );
   nand U20832 ( n19891,n21474,n21475,n21476 );
   nand U20833 ( n21476,n19960,n19578 );
   nand U20834 ( n21475,n21477,n19818 );
   xor U20835 ( n21477,n21478,n20182 );
   nand U20836 ( n21474,n19895,n20909 );
   and U20837 ( n21469,n20902,p2_reg2_reg_19_ );
   nand U20838 ( n21467,n20913,n19572 );
   nand U20839 ( n21466,n20932,n19894 );
   xor U20840 ( n19894,n20530,n21456 );
   nand U20841 ( n21465,n20917,n19895 );
   xor U20842 ( n19895,n20182,n21479 );
   nand U20843 ( n20182,n21480,n21481 );
   nand U20844 ( p2_u3245,n21482,n21483,n21484,n21485 );
   nor U20845 ( n21485,n21486,n21487,n21488,n21489 );
   nor U20846 ( n21489,n21490,n20915 );
   nor U20847 ( n21488,n21491,n21068 );
   nor U20848 ( n21487,n19875,n20902 );
   and U20849 ( n19875,n21492,n21493,n21494,n21495 );
   nor U20850 ( n21495,n21496,n21497,n21498,n21499 );
   nor U20851 ( n21499,n21078,n19882 );
   nor U20852 ( n21498,n21043,n19882 );
   nor U20853 ( n21497,n20608,n19882 );
   nor U20854 ( n21496,n21040,n21500 );
   nor U20855 ( n21494,n21501,n21502 );
   nor U20856 ( n21502,n19906,n19776 );
   nor U20857 ( n21501,n20600,n21500 );
   nand U20858 ( n21493,n21503,n20968 );
   nand U20859 ( n21492,n21503,n20967 );
   not U20860 ( n21503,n21500 );
   xor U20861 ( n21500,n20183,n21504 );
   and U20862 ( n21486,n20902,p2_reg2_reg_20_ );
   nand U20863 ( n21484,n20913,n19569 );
   or U20864 ( n21483,n20916,n19881 );
   nand U20865 ( n19881,n21505,n21506 );
   nand U20866 ( n21506,n19883,n21507 );
   nand U20867 ( n21507,n21508,n19892 );
   or U20868 ( n21482,n21222,n19882 );
   nand U20869 ( n19882,n21509,n21510 );
   nand U20870 ( n21510,n21511,n21512,n21513 );
   nand U20871 ( n21511,n21479,n21480 );
   nand U20872 ( n21509,n20183,n21480,n21514 );
   nand U20873 ( n21514,n21515,n21481 );
   nand U20874 ( n20183,n21512,n21516 );
   nand U20875 ( p2_u3244,n21517,n21518,n21519,n21520 );
   nor U20876 ( n21520,n21521,n21522,n21523,n21524 );
   nor U20877 ( n21524,n21525,n20915 );
   and U20878 ( n21523,n21526,n20912 );
   nor U20879 ( n21522,n19863,n20902 );
   and U20880 ( n19863,n21527,n21528,n21529,n21530 );
   nor U20881 ( n21530,n21531,n21532 );
   nor U20882 ( n21532,n21533,n19776 );
   nor U20883 ( n21531,n21534,n21535,n21536 );
   nor U20884 ( n21536,n21537,n21538,n21539 );
   and U20885 ( n21535,n21537,n21540 );
   nand U20886 ( n21529,n21541,n21542 );
   nand U20887 ( n21528,n21543,n21544,n20968 );
   not U20888 ( n20968,n20609 );
   nand U20889 ( n21544,n21540,n21537 );
   nand U20890 ( n21543,n21545,n21546 );
   nand U20891 ( n21527,n21053,n21547,n21548,n21549 );
   not U20892 ( n21053,n21078 );
   and U20893 ( n21521,n20902,p2_reg2_reg_21_ );
   nand U20894 ( n21519,n20913,n19566 );
   or U20895 ( n21518,n20916,n19870 );
   xor U20896 ( n19870,n21505,n21525 );
   nand U20897 ( n21517,n20917,n21541 );
   not U20898 ( n21541,n19869 );
   nand U20899 ( n19869,n21548,n21549,n21547 );
   nand U20900 ( n21547,n21513,n21515,n21540 );
   nand U20901 ( n21549,n21540,n21550 );
   not U20902 ( n21540,n20184 );
   nand U20903 ( n21548,n21551,n20184,n21552 );
   nand U20904 ( n20184,n21553,n21554 );
   nand U20905 ( n21551,n21513,n21515 );
   not U20906 ( n21515,n21479 );
   nor U20907 ( n21479,n21463,n21555 );
   nand U20908 ( p2_u3243,n21556,n21557,n21558,n21559 );
   nor U20909 ( n21559,n21560,n21561,n21562,n21563 );
   nor U20910 ( n21563,n19832,n20929 );
   nor U20911 ( n21562,n19859,n20916 );
   nand U20912 ( n19859,n21564,n21565 );
   nand U20913 ( n21565,n20562,n21566 );
   nand U20914 ( n21566,n21567,n21525 );
   and U20915 ( n21561,n20936,n19860 );
   xor U20916 ( n19860,n20204,n21568 );
   nor U20917 ( n21560,n19857,n20959 );
   nor U20918 ( n21558,n21569,n21570 );
   nor U20919 ( n21570,n20902,n19851 );
   nand U20920 ( n19851,n21571,n21572,n19818 );
   nand U20921 ( n21572,n20204,n21573 );
   xor U20922 ( n20204,n19566,n20562 );
   nand U20923 ( n21571,n21574,n21575,n21576 );
   and U20924 ( n21569,n20902,p2_reg2_reg_22_ );
   nand U20925 ( n21557,n20912,n21577 );
   nand U20926 ( n21556,n21003,n20562 );
   nand U20927 ( p2_u3242,n21578,n21579,n21580,n21581 );
   nor U20928 ( n21581,n21582,n21583,n21584,n21585 );
   nor U20929 ( n21585,n21586,n20915 );
   and U20930 ( n21584,n21587,n20912 );
   nor U20931 ( n21583,n19839,n20902 );
   and U20932 ( n19839,n21588,n21589,n21590,n21591 );
   nor U20933 ( n21591,n21592,n21593,n21594,n21595 );
   nor U20934 ( n21595,n19871,n19776 );
   nor U20935 ( n21594,n21078,n19845 );
   nor U20936 ( n21593,n20608,n19845 );
   not U20937 ( n19845,n21596 );
   nor U20938 ( n21592,n21597,n20609 );
   nor U20939 ( n21590,n21598,n21599 );
   nor U20940 ( n21599,n21597,n21040 );
   nor U20941 ( n21598,n21597,n20600 );
   and U20942 ( n21597,n21600,n21601 );
   nand U20943 ( n21600,n21602,n21603 );
   nand U20944 ( n21603,n21575,n21576 );
   not U20945 ( n21602,n21604 );
   nand U20946 ( n21589,n21596,n20602 );
   not U20947 ( n20602,n21043 );
   nand U20948 ( n21588,n21605,n21606,n20967 );
   not U20949 ( n20967,n21042 );
   nand U20950 ( n21606,n21576,n21575,n21607 );
   not U20951 ( n21576,n21573 );
   nand U20952 ( n21605,n21601,n21604 );
   nand U20953 ( n21604,n21607,n21574 );
   nand U20954 ( n21601,n21608,n21609 );
   nand U20955 ( n21609,n21573,n21574 );
   nor U20956 ( n21573,n21545,n21538 );
   and U20957 ( n21608,n20203,n21575 );
   and U20958 ( n21582,n20902,p2_reg2_reg_23_ );
   nand U20959 ( n21580,n20913,n19560 );
   or U20960 ( n21579,n20916,n19846 );
   xor U20961 ( n19846,n21564,n21586 );
   nand U20962 ( n21578,n20917,n21596 );
   xor U20963 ( n21596,n21607,n21610 );
   not U20964 ( n21607,n20203 );
   xor U20965 ( n20203,n19832,n21586 );
   not U20966 ( n20917,n21222 );
   nand U20967 ( p2_u3241,n21611,n21612,n21613,n21614 );
   nor U20968 ( n21614,n21615,n21616,n21617,n21618 );
   and U20969 ( n21618,n20902,p2_reg2_reg_24_ );
   nor U20970 ( n21617,n19833,n20915 );
   and U20971 ( n21616,n21619,n20912 );
   nor U20972 ( n21615,n19831,n20929 );
   nor U20973 ( n21613,n21620,n21621 );
   nor U20974 ( n21621,n19834,n20916 );
   nand U20975 ( n19834,n21622,n21623 );
   nand U20976 ( n21623,n20557,n21624 );
   nand U20977 ( n21624,n21625,n21586 );
   and U20978 ( n21620,n20936,n19835 );
   xor U20979 ( n19835,n21626,n20185 );
   nand U20980 ( n21612,n20933,n19836 );
   xor U20981 ( n19836,n20185,n21627 );
   nand U20982 ( n20185,n21628,n21629 );
   nand U20983 ( n21611,n20935,n19563 );
   not U20984 ( n20935,n20959 );
   nand U20985 ( p2_u3240,n21630,n21631,n21632,n21633 );
   nor U20986 ( n21633,n21634,n21635,n21636,n21637 );
   and U20987 ( n21637,n20902,p2_reg2_reg_25_ );
   nor U20988 ( n21636,n19816,n20915 );
   and U20989 ( n21635,n21638,n20912 );
   nor U20990 ( n21634,n19814,n20929 );
   nor U20991 ( n21632,n21639,n21640 );
   and U20992 ( n21640,n20936,n19820 );
   xor U20993 ( n19820,n20186,n21641 );
   nor U20994 ( n21639,n19815,n20959 );
   nand U20995 ( n21631,n20933,n19817 );
   xor U20996 ( n19817,n21642,n21643 );
   not U20997 ( n21642,n20186 );
   nand U20998 ( n20186,n21644,n21645 );
   nor U20999 ( n20933,n20902,n21646 );
   nand U21000 ( n21630,n20932,n19819 );
   xor U21001 ( n19819,n21647,n19816 );
   nand U21002 ( p2_u3239,n21648,n21649,n21650,n21651 );
   nor U21003 ( n21651,n21652,n21653,n21654,n21655 );
   nor U21004 ( n21655,n21656,n20915 );
   nor U21005 ( n21654,n21657,n21068 );
   nor U21006 ( n21653,n19796,n20902 );
   and U21007 ( n19796,n21658,n21659,n21660,n21661 );
   nor U21008 ( n21661,n21662,n21663,n21664,n21665 );
   nor U21009 ( n21665,n21078,n19803 );
   nor U21010 ( n21664,n21043,n19803 );
   nor U21011 ( n21663,n20608,n19803 );
   nor U21012 ( n21662,n21042,n21666,n21667 );
   nor U21013 ( n21660,n21668,n21669 );
   nor U21014 ( n21669,n20609,n21666,n21667 );
   nor U21015 ( n21668,n20600,n21666,n21667 );
   and U21016 ( n21667,n21670,n21671 );
   nor U21017 ( n21666,n20187,n21672 );
   nand U21018 ( n21659,n19960,n19557 );
   nand U21019 ( n21658,n21673,n21674,n20969 );
   nand U21020 ( n21674,n21675,n21676 );
   or U21021 ( n21673,n21677,n21678,n21676 );
   and U21022 ( n21652,n20902,p2_reg2_reg_26_ );
   nand U21023 ( n21650,n20913,n19551 );
   or U21024 ( n21649,n20916,n19802 );
   nand U21025 ( n19802,n21679,n21680 );
   nand U21026 ( n21680,n19804,n21681 );
   nand U21027 ( n21681,n21647,n19816 );
   or U21028 ( n21648,n21222,n19803 );
   nand U21029 ( n19803,n21682,n21683 );
   nand U21030 ( n21683,n21684,n21645,n20187 );
   nand U21031 ( n21684,n21685,n21644 );
   not U21032 ( n21685,n21641 );
   nand U21033 ( n21682,n21686,n21644,n21675 );
   not U21034 ( n21675,n20187 );
   nand U21035 ( n20187,n21687,n21688 );
   nand U21036 ( n21686,n21645,n21641 );
   nand U21037 ( n21641,n21628,n21689 );
   nand U21038 ( n21689,n21629,n21626 );
   nand U21039 ( p2_u3238,n21690,n21691,n21692,n21693 );
   nor U21040 ( n21693,n21694,n21695,n21696,n21697 );
   nor U21041 ( n21697,n21698,n20915 );
   and U21042 ( n21696,n21699,n20912 );
   nor U21043 ( n21695,n19784,n20902 );
   and U21044 ( n19784,n21700,n21701,n21702,n21703 );
   nor U21045 ( n21703,n21704,n21705,n21706,n21707 );
   nor U21046 ( n21707,n21708,n21042 );
   nor U21047 ( n21708,n21709,n21710 );
   nor U21048 ( n21710,n20188,n21677,n21711 );
   nor U21049 ( n21711,n21678,n21672 );
   not U21050 ( n21672,n21676 );
   not U21051 ( n21709,n21712 );
   nor U21052 ( n21706,n19790,n21043 );
   and U21053 ( n21705,n21713,n20969 );
   nor U21054 ( n21704,n19790,n21078 );
   nor U21055 ( n21702,n21714,n21715 );
   nor U21056 ( n21715,n19790,n20608 );
   nor U21057 ( n21714,n21716,n20609 );
   xor U21058 ( n21716,n21717,n20188 );
   nand U21059 ( n21701,n20607,n21713 );
   nand U21060 ( n21713,n21718,n21712 );
   nand U21061 ( n21712,n21717,n20188 );
   or U21062 ( n21718,n20188,n21717 );
   nor U21063 ( n21717,n21678,n21670 );
   nand U21064 ( n21700,n19960,n19554 );
   and U21065 ( n21694,n20902,p2_reg2_reg_27_ );
   nand U21066 ( n21692,n20913,n19548 );
   not U21067 ( n20913,n20929 );
   or U21068 ( n21691,n20916,n19791 );
   xor U21069 ( n19791,n21679,n21698 );
   or U21070 ( n21690,n21222,n19790 );
   xor U21071 ( n19790,n20188,n21719 );
   nand U21072 ( n21719,n21720,n21721,n21688 );
   nand U21073 ( n21688,n19804,n19554 );
   nand U21074 ( n21720,n21722,n21723 );
   nand U21075 ( n20188,n21724,n21725 );
   nand U21076 ( p2_u3237,n21726,n21727,n21728,n21729 );
   nor U21077 ( n21729,n21730,n21731,n21732,n21733 );
   and U21078 ( n21733,n19779,n20932 );
   nor U21079 ( n19779,n21734,n21735 );
   and U21080 ( n21735,n20575,n21736 );
   nand U21081 ( n21736,n21737,n21698 );
   not U21082 ( n21737,n21679 );
   nor U21083 ( n21732,n19773,n20929 );
   nand U21084 ( n20929,n20910,n19893 );
   not U21085 ( n19893,n19774 );
   nor U21086 ( n21731,n20951,n19780 );
   xor U21087 ( n19780,n21738,n21739 );
   nor U21088 ( n21738,n21740,n21741 );
   not U21089 ( n20951,n20936 );
   nand U21090 ( n20936,n21222,n21742 );
   nand U21091 ( n21742,n20910,n20909 );
   nor U21092 ( n21730,n19775,n20959 );
   nand U21093 ( n20959,n20910,n19960 );
   nor U21094 ( n21728,n21743,n21744 );
   nor U21095 ( n21744,n19778,n20915 );
   and U21096 ( n21743,n21745,n20912 );
   nand U21097 ( n21727,p2_reg2_reg_28_,n20902 );
   or U21098 ( n21726,n19767,n20902 );
   nand U21099 ( n19767,n21746,n21747 );
   xor U21100 ( n21746,n21748,n20192 );
   not U21101 ( n20192,n21739 );
   nor U21102 ( n21739,n21749,n21750 );
   nor U21103 ( n21749,n19548,n20575 );
   nand U21104 ( p2_u3236,n21751,n21752,n21753,n21754 );
   nor U21105 ( n21754,n21755,n21756,n21757 );
   nor U21106 ( n21757,n19758,n20916 );
   xor U21107 ( n19758,n21734,n19762 );
   and U21108 ( n21756,n21758,n20912 );
   not U21109 ( n20912,n21068 );
   nand U21110 ( n21068,n21759,n20910 );
   nor U21111 ( n21755,n19761,n21222 );
   nand U21112 ( n21753,n21003,n19762 );
   not U21113 ( n19762,n21761 );
   nand U21114 ( n21752,p2_reg2_reg_29_,n20902 );
   nand U21115 ( n21751,n20910,n19763 );
   nand U21116 ( n19763,n21762,n21763,n21764,n21765 );
   nor U21117 ( n21765,n21766,n21767 );
   nor U21118 ( n21767,n20127,n19761 );
   xor U21119 ( n19761,n20196,n21768 );
   nand U21120 ( n21768,n21769,n21770 );
   or U21121 ( n21770,n21740,n21750,n21741 );
   nand U21122 ( n21741,n21771,n21724,n21772 );
   nand U21123 ( n21772,n19554,n21725,n19804 );
   not U21124 ( n19804,n21656 );
   nand U21125 ( n21724,n19793,n19551 );
   nand U21126 ( n21771,n21723,n21725,n21722 );
   not U21127 ( n21725,n21773 );
   nand U21128 ( n21723,n21645,n21629 );
   nand U21129 ( n21629,n20557,n19560 );
   nand U21130 ( n21645,n20546,n19557 );
   nor U21131 ( n21740,n21721,n21773 );
   nor U21132 ( n21773,n19551,n19793 );
   nand U21133 ( n21721,n21722,n21628,n21774 );
   not U21134 ( n21774,n21626 );
   nand U21135 ( n21626,n21775,n21776 );
   nand U21136 ( n21776,n21777,n21586 );
   or U21137 ( n21777,n21610,n19832 );
   nand U21138 ( n21775,n19832,n21610 );
   nand U21139 ( n21610,n21778,n21779 );
   nand U21140 ( n21779,n21780,n19858 );
   nand U21141 ( n21780,n19566,n21568 );
   or U21142 ( n21778,n21568,n19566 );
   nand U21143 ( n21568,n21781,n21553,n21782 );
   nand U21144 ( n21782,n21554,n21783 );
   nand U21145 ( n21783,n21552,n21784 );
   nand U21146 ( n21784,n21463,n21513 );
   nor U21147 ( n21463,n19908,n19922 );
   not U21148 ( n21552,n21550 );
   nand U21149 ( n21550,n21512,n21785 );
   nand U21150 ( n21785,n21786,n21516 );
   not U21151 ( n21786,n21480 );
   nand U21152 ( n21480,n20530,n19575 );
   nand U21153 ( n21512,n19883,n19572 );
   nand U21154 ( n21553,n19872,n19569 );
   not U21155 ( n19872,n21525 );
   nand U21156 ( n21781,n21513,n21554,n21555 );
   and U21157 ( n21555,n21787,n21460 );
   nand U21158 ( n21460,n21443,n21788 );
   nand U21159 ( n21788,n21789,n21442 );
   nand U21160 ( n21442,n19907,n21421 );
   nand U21161 ( n21789,n21411,n21440 );
   nand U21162 ( n21440,n21790,n21412 );
   nand U21163 ( n21412,n19944,n21378 );
   not U21164 ( n21790,n21410 );
   nand U21165 ( n21410,n21791,n21792 );
   nand U21166 ( n21792,n19946,n21793 );
   nand U21167 ( n21793,n21360,n19587 );
   not U21168 ( n21360,n21794 );
   nand U21169 ( n21791,n19959,n21794 );
   nand U21170 ( n21794,n21795,n21796 );
   nand U21171 ( n21796,n19958,n21797 );
   nand U21172 ( n21797,n19590,n21798 );
   nand U21173 ( n21795,n21337,n19945 );
   not U21174 ( n21337,n21798 );
   nand U21175 ( n21798,n21799,n21800 );
   nand U21176 ( n21800,n21323,n21290,n21324 );
   and U21177 ( n21324,n21270,n21801 );
   nand U21178 ( n21801,n19984,n21238 );
   nand U21179 ( n21270,n21228,n21802 );
   nand U21180 ( n21802,n21803,n21227 );
   nand U21181 ( n21227,n20021,n21197 );
   nand U21182 ( n21803,n21183,n21225 );
   nand U21183 ( n21225,n21184,n21179 );
   nand U21184 ( n21179,n21804,n21166 );
   nand U21185 ( n21166,n20038,n19608 );
   nand U21186 ( n21804,n21165,n21167 );
   nand U21187 ( n21167,n20022,n21139 );
   and U21188 ( n21165,n21805,n21128 );
   nand U21189 ( n21128,n20060,n21102 );
   nand U21190 ( n21805,n21129,n21088,n21126 );
   nand U21191 ( n21126,n21087,n21089 );
   nand U21192 ( n21089,n21113,n21066 );
   not U21193 ( n21087,n21130 );
   nand U21194 ( n21130,n21806,n21056 );
   nand U21195 ( n21056,n20082,n21030 );
   nand U21196 ( n21806,n21055,n21057 );
   nand U21197 ( n21057,n20072,n19617 );
   nand U21198 ( n21055,n21807,n21808 );
   nand U21199 ( n21808,n21809,n20084 );
   nand U21200 ( n21809,n19620,n21018 );
   or U21201 ( n21807,n19620,n21018 );
   nand U21202 ( n21018,n21810,n21811,n21812 );
   nand U21203 ( n21812,n21813,n19623 );
   nand U21204 ( n21811,n21814,n20973,n20957 );
   nor U21205 ( n20957,n20919,n20939 );
   nor U21206 ( n20939,n19629,n20338 );
   nand U21207 ( n20919,n20135,n19632 );
   nand U21208 ( n21814,n20083,n21015 );
   nand U21209 ( n21810,n20100,n21815 );
   nand U21210 ( n21815,n20986,n20083 );
   not U21211 ( n20986,n21813 );
   nand U21212 ( n21813,n20974,n21816 );
   nand U21213 ( n21816,n20938,n20973 );
   nand U21214 ( n20973,n20099,n20110 );
   nor U21215 ( n20938,n20123,n20958 );
   nand U21216 ( n20974,n20297,n19626 );
   nand U21217 ( n21088,n20061,n19614 );
   nand U21218 ( n21129,n20049,n19611 );
   nand U21219 ( n21184,n20037,n20023 );
   nand U21220 ( n21183,n20414,n19605 );
   nand U21221 ( n21799,n21323,n21817 );
   nand U21222 ( n21817,n21322,n21291,n21818 );
   nand U21223 ( n21818,n21271,n21290 );
   nand U21224 ( n21290,n19999,n19985 );
   nor U21225 ( n21271,n21238,n19984 );
   nand U21226 ( n21291,n20429,n19596 );
   not U21227 ( n20429,n19985 );
   nand U21228 ( n21322,n19973,n19593 );
   nand U21229 ( n21323,n19983,n21300 );
   nand U21230 ( n21411,n19934,n19584 );
   nand U21231 ( n21443,n19923,n19581 );
   nand U21232 ( n21787,n19922,n19908 );
   nand U21233 ( n21554,n19857,n21525 );
   and U21234 ( n21513,n21481,n21516 );
   nand U21235 ( n21516,n21533,n21490 );
   nand U21236 ( n21481,n19906,n19892 );
   nand U21237 ( n21628,n19815,n19833 );
   and U21238 ( n21722,n21644,n21687 );
   nand U21239 ( n21687,n19814,n21656 );
   nand U21240 ( n21644,n19831,n19816 );
   nand U21241 ( n21769,n19792,n19778 );
   not U21242 ( n20127,n20909 );
   nand U21243 ( n20909,n21819,n21078 );
   nand U21244 ( n21078,n20603,n21820 );
   not U21245 ( n21819,n21542 );
   nand U21246 ( n21542,n21043,n20608 );
   nor U21247 ( n21766,n20211,n21821 );
   not U21248 ( n20211,n19542 );
   nand U21249 ( n19542,n21822,n21823,n21824 );
   nand U21250 ( n21824,p2_reg2_reg_30_,n21825 );
   nand U21251 ( n21823,p2_reg0_reg_30_,n21826 );
   nand U21252 ( n21822,p2_reg1_reg_30_,n21827 );
   nand U21253 ( n21764,n19960,n19548 );
   not U21254 ( n19960,n19776 );
   nand U21255 ( n21763,n20196,n21829 );
   nand U21256 ( n21829,n21830,n21831 );
   nand U21257 ( n21831,n21832,n21747 );
   nand U21258 ( n21747,n21833,n21042 );
   not U21259 ( n21833,n20994 );
   nand U21260 ( n20994,n20223,n20609 );
   not U21261 ( n21832,n21834 );
   or U21262 ( n21830,n21835,n21646 );
   nand U21263 ( n21762,n19818,n21834,n21835,n21836 );
   not U21264 ( n21836,n20196 );
   xor U21265 ( n20196,n19773,n21761 );
   not U21266 ( n19773,n19545 );
   nand U21267 ( n21835,n21837,n21748 );
   nand U21268 ( n21748,n21838,n21839 );
   nand U21269 ( n21839,n21840,n21841 );
   nand U21270 ( n21841,n19793,n21842 );
   nand U21271 ( n21842,n21678,n19551 );
   not U21272 ( n21678,n21671 );
   nand U21273 ( n21840,n19775,n21671 );
   nand U21274 ( n21671,n21656,n19554 );
   nand U21275 ( n21838,n21670,n21843 );
   nand U21276 ( n21843,n19775,n19793 );
   nor U21277 ( n21670,n21676,n21677 );
   nor U21278 ( n21677,n21656,n19554 );
   nand U21279 ( n21676,n21844,n21845 );
   nand U21280 ( n21845,n20546,n21846 );
   or U21281 ( n21846,n21643,n19831 );
   not U21282 ( n20546,n19816 );
   nand U21283 ( n21844,n19831,n21643 );
   nand U21284 ( n21643,n21847,n21848 );
   nand U21285 ( n21848,n20557,n21849 );
   nand U21286 ( n21849,n19560,n21627 );
   not U21287 ( n20557,n19833 );
   or U21288 ( n21847,n21627,n19560 );
   nand U21289 ( n21627,n21850,n21851 );
   nand U21290 ( n21851,n21852,n21575,n21545 );
   nor U21291 ( n21545,n21537,n21539 );
   nor U21292 ( n21539,n19569,n21525 );
   nand U21293 ( n21537,n21853,n21854 );
   nand U21294 ( n21854,n19883,n21855 );
   or U21295 ( n21855,n21504,n21533 );
   nand U21296 ( n21853,n21533,n21504 );
   nand U21297 ( n21504,n21856,n21857 );
   nand U21298 ( n21857,n19906,n21858 );
   nand U21299 ( n21858,n21478,n19892 );
   not U21300 ( n21478,n21859 );
   nand U21301 ( n21856,n20530,n21859 );
   nand U21302 ( n21859,n21860,n21861 );
   nand U21303 ( n21861,n20525,n21862 );
   or U21304 ( n21862,n21462,n19922 );
   nand U21305 ( n21860,n19922,n21462 );
   nand U21306 ( n21462,n21863,n21864 );
   nand U21307 ( n21864,n19923,n21865 );
   nand U21308 ( n21865,n19581,n21436 );
   not U21309 ( n19923,n21421 );
   or U21310 ( n21863,n21436,n19581 );
   nand U21311 ( n21436,n21866,n21867 );
   nand U21312 ( n21867,n21404,n21868 );
   nand U21313 ( n21868,n21403,n21869 );
   nand U21314 ( n21869,n21402,n21405 );
   not U21315 ( n21402,n21346 );
   nand U21316 ( n21346,n19958,n19590 );
   and U21317 ( n21403,n21366,n21870 );
   nand U21318 ( n21870,n21378,n19584 );
   nand U21319 ( n21366,n19946,n19587 );
   nand U21320 ( n21866,n21404,n21405,n21345 );
   and U21321 ( n21345,n21351,n21350 );
   nand U21322 ( n21350,n19945,n20389 );
   not U21323 ( n21351,n21349 );
   nand U21324 ( n21349,n21871,n21872 );
   nand U21325 ( n21872,n19973,n21873 );
   nand U21326 ( n21873,n21314,n19593 );
   not U21327 ( n21314,n21874 );
   nand U21328 ( n21871,n19983,n21874 );
   nand U21329 ( n21874,n21875,n21876 );
   nand U21330 ( n21876,n19999,n21877 );
   nand U21331 ( n21877,n19985,n21289 );
   or U21332 ( n21875,n21289,n19985 );
   nand U21333 ( n21289,n21878,n21879 );
   nand U21334 ( n21879,n21268,n21880 );
   nand U21335 ( n21880,n21267,n21881 );
   nand U21336 ( n21881,n21262,n21213 );
   not U21337 ( n21262,n21188 );
   nand U21338 ( n21188,n20023,n19605 );
   and U21339 ( n21267,n21212,n21882 );
   nand U21340 ( n21882,n21238,n19599 );
   nand U21341 ( n21878,n21268,n21213,n21261 );
   and U21342 ( n21261,n21185,n21187 );
   nand U21343 ( n21187,n20414,n20037 );
   not U21344 ( n20037,n19605 );
   nand U21345 ( n21185,n21883,n21884 );
   nand U21346 ( n21884,n21885,n19608 );
   nand U21347 ( n21885,n21150,n20038 );
   nand U21348 ( n21883,n21159,n21139 );
   not U21349 ( n21159,n21150 );
   nor U21350 ( n21150,n21886,n21120 );
   nor U21351 ( n21120,n21119,n21887 );
   nor U21352 ( n21887,n21102,n19611 );
   nand U21353 ( n21119,n21888,n21889 );
   nand U21354 ( n21889,n21086,n21050,n21890 );
   nand U21355 ( n21890,n21066,n19614 );
   nand U21356 ( n21050,n21030,n19617 );
   nand U21357 ( n21086,n21049,n21051 );
   nand U21358 ( n21051,n21891,n21892 );
   nand U21359 ( n21892,n21893,n21020 );
   nand U21360 ( n21020,n21894,n21895 );
   nand U21361 ( n21895,n21896,n21015 );
   nand U21362 ( n21896,n21000,n20083 );
   not U21363 ( n21000,n21897 );
   nand U21364 ( n21894,n21897,n19623 );
   nand U21365 ( n21897,n20955,n21898 );
   nand U21366 ( n21898,n20972,n20956 );
   nand U21367 ( n20956,n20099,n20297 );
   not U21368 ( n20972,n20999 );
   nand U21369 ( n20999,n21899,n21900 );
   nand U21370 ( n21900,n21901,n20338 );
   nand U21371 ( n21901,n19629,n20906 );
   nand U21372 ( n21899,n20934,n20958 );
   not U21373 ( n20934,n20906 );
   nand U21374 ( n20906,n20122,n20135 );
   not U21375 ( n20122,n19632 );
   nand U21376 ( n20955,n20110,n19626 );
   nand U21377 ( n21893,n20318,n20983 );
   nand U21378 ( n21891,n20084,n19620 );
   nand U21379 ( n21049,n20072,n20082 );
   nand U21380 ( n21888,n21113,n20061 );
   not U21381 ( n21886,n21121 );
   nand U21382 ( n21121,n21102,n19611 );
   nand U21383 ( n21213,n20021,n20011 );
   nand U21384 ( n21268,n20000,n19984 );
   not U21385 ( n19983,n19593 );
   nand U21386 ( n21405,n19959,n20371 );
   not U21387 ( n19959,n19587 );
   nand U21388 ( n21404,n19934,n19944 );
   not U21389 ( n19922,n19578 );
   not U21390 ( n20530,n19892 );
   nand U21391 ( n21850,n21902,n21852 );
   nand U21392 ( n21852,n19847,n19832 );
   not U21393 ( n19832,n19563 );
   not U21394 ( n19847,n21586 );
   nand U21395 ( n21902,n21903,n21574,n21904 );
   nand U21396 ( n21904,n21586,n19563 );
   nand U21397 ( n21574,n19858,n19566 );
   nand U21398 ( n21903,n21538,n21575 );
   nand U21399 ( n21575,n20562,n19871 );
   not U21400 ( n19871,n19566 );
   not U21401 ( n20562,n19858 );
   not U21402 ( n21538,n21546 );
   nand U21403 ( n21546,n21525,n19569 );
   nand U21404 ( p2_u3235,n21905,n21906,n21907,n21908 );
   nand U21405 ( n21908,p2_reg2_reg_30_,n20902 );
   nand U21406 ( n21906,n19750,n19751,n20932 );
   nand U21407 ( n19750,n19748,n21909 );
   nand U21408 ( n21909,n21734,n21761 );
   nand U21409 ( n21905,n21003,n19748 );
   not U21410 ( n19748,n20212 );
   nand U21411 ( p2_u3234,n21910,n21911,n21907,n21912 );
   nand U21412 ( n21912,p2_reg2_reg_31_,n20902 );
   nand U21413 ( n21907,n19749,n20910 );
   nor U21414 ( n19749,n21821,n20593 );
   not U21415 ( n20593,n19539 );
   nand U21416 ( n19539,n21913,n21914,n21915 );
   nand U21417 ( n21915,p2_reg2_reg_31_,n21825 );
   nand U21418 ( n21914,p2_reg0_reg_31_,n21826 );
   nand U21419 ( n21913,p2_reg1_reg_31_,n21827 );
   and U21420 ( n21821,n21916,n21917 );
   or U21421 ( n21917,n19774,p2_b_reg );
   nand U21422 ( n21916,n21918,n20148 );
   nand U21423 ( n21911,n20932,n19742 );
   xor U21424 ( n19742,n19740,n19751 );
   nand U21425 ( n19751,n21761,n20212,n21734 );
   nor U21426 ( n21734,n20575,n19793,n21679 );
   nand U21427 ( n21679,n19816,n21656,n21647 );
   not U21428 ( n21647,n21622 );
   nand U21429 ( n21622,n21586,n19833,n21625 );
   not U21430 ( n21625,n21564 );
   nand U21431 ( n21564,n19858,n21525,n21567 );
   not U21432 ( n21567,n21505 );
   nand U21433 ( n21505,n21490,n19892,n21508 );
   not U21434 ( n21508,n21456 );
   nand U21435 ( n21456,n19908,n21421,n21459 );
   not U21436 ( n21459,n21406 );
   nand U21437 ( n21406,n19946,n21378,n21409 );
   not U21438 ( n21409,n21333 );
   nand U21439 ( n21333,n19958,n21300,n21336 );
   not U21440 ( n21336,n21284 );
   nand U21441 ( n21284,n21238,n19985,n21287 );
   not U21442 ( n21287,n21218 );
   nand U21443 ( n21218,n21197,n20023,n21221 );
   not U21444 ( n21221,n21161 );
   nand U21445 ( n21161,n21139,n21102,n21164 );
   not U21446 ( n21164,n21090 );
   nand U21447 ( n21090,n21066,n21030,n21093 );
   not U21448 ( n21093,n21012 );
   nand U21449 ( n21012,n20084,n21015,n20988 );
   not U21450 ( n20988,n20948 );
   nand U21451 ( n20948,n20123,n20908,n20110 );
   not U21452 ( n20908,n20135 );
   not U21453 ( n19793,n21698 );
   nand U21454 ( n20212,n21919,n21920,n21921 );
   nand U21455 ( n21920,n16576,n17674 );
   not U21456 ( n17674,p1_datao_reg_30_ );
   or U21457 ( n21919,n20869,n16576 );
   nand U21458 ( n21761,n21922,n21923,n21921 );
   nand U21459 ( n21923,n16576,n17679 );
   or U21460 ( n21922,n20860,n16576 );
   nor U21461 ( n20932,n20902,n21924 );
   nand U21462 ( n21910,n21003,n19740 );
   and U21463 ( n19740,n20874,n21921 );
   and U21464 ( n20874,n21925,n21926 );
   nand U21465 ( n21926,n16576,n17669 );
   not U21466 ( n17669,p1_datao_reg_31_ );
   nand U21467 ( n21925,n21927,n16572 );
   not U21468 ( n21003,n20915 );
   nand U21469 ( n21928,n21929,n21930 );
   nand U21470 ( n21930,n21931,n21932,n20140,n20144 );
   nand U21471 ( p2_u3233,n21933,n21934,n21935 );
   nor U21472 ( n21935,n21936,n21937,n21938 );
   nor U21473 ( n21938,n21939,n21940 );
   xor U21474 ( n21940,n21941,n21942 );
   nand U21475 ( n21942,n21943,n21944 );
   nand U21476 ( n21944,p2_reg2_reg_18_,n21945 );
   or U21477 ( n21945,n21946,n21947 );
   nand U21478 ( n21943,n21947,n21946 );
   xor U21479 ( n21941,p2_reg2_reg_19_,n21948 );
   nor U21480 ( n21937,n21949,n21950 );
   xor U21481 ( n21950,n21951,n21952 );
   nand U21482 ( n21952,n21953,n21954 );
   nand U21483 ( n21954,p2_reg1_reg_18_,n21955 );
   or U21484 ( n21955,n21946,n21956 );
   nand U21485 ( n21953,n21956,n21946 );
   xor U21486 ( n21951,p2_reg1_reg_19_,n21948 );
   nor U21487 ( n21936,n21948,n21957 );
   nand U21488 ( n21934,n21958,p2_addr_reg_19_ );
   nand U21489 ( n21933,p2_reg3_reg_19_,p2_u3088 );
   nand U21490 ( p2_u3232,n21959,n21960,n21961,n21962 );
   nand U21491 ( n21962,n21963,n21964 );
   nand U21492 ( n21964,n21965,n21966 );
   nand U21493 ( n21966,n21967,n21968 );
   nand U21494 ( n21965,n21969,n21970 );
   xor U21495 ( n21970,n21947,p2_reg2_reg_18_ );
   nand U21496 ( n21961,n21946,n21971 );
   nand U21497 ( n21971,n21972,n21957,n21973 );
   nand U21498 ( n21973,n21974,n21969 );
   xor U21499 ( n21974,n21452,n21947 );
   nor U21500 ( n21947,n21975,n21976 );
   nor U21501 ( n21975,n21977,n21978 );
   not U21502 ( n21452,p2_reg2_reg_18_ );
   or U21503 ( n21972,n21968,n21949 );
   xor U21504 ( n21968,n21956,p2_reg1_reg_18_ );
   nor U21505 ( n21956,n21979,n21980 );
   nor U21506 ( n21979,n21981,n21982 );
   not U21507 ( n21946,n21963 );
   nand U21508 ( n21960,n21958,p2_addr_reg_18_ );
   nand U21509 ( n21959,p2_reg3_reg_18_,p2_u3088 );
   nand U21510 ( p2_u3231,n21983,n21984,n21985 );
   nor U21511 ( n21985,n21986,n21987,n21988 );
   nor U21512 ( n21988,n21939,n21989,n21990 );
   nor U21513 ( n21990,n21977,n21991 );
   xor U21514 ( n21991,n21992,n21437 );
   nand U21515 ( n21977,n21993,n21994 );
   or U21516 ( n21994,n21995,n21996 );
   nor U21517 ( n21989,n21996,n21978,n21997,n21976 );
   nor U21518 ( n21976,p2_reg2_reg_17_,n21998 );
   not U21519 ( n21997,n21999 );
   nor U21520 ( n21978,n21992,n21437 );
   not U21521 ( n21437,p2_reg2_reg_17_ );
   nor U21522 ( n21987,n21949,n22000,n22001 );
   nor U21523 ( n22001,n21981,n22002 );
   xor U21524 ( n22002,n21998,p2_reg1_reg_17_ );
   nand U21525 ( n21981,n22003,n22004 );
   or U21526 ( n22004,n22005,n22006 );
   nor U21527 ( n22000,n22006,n21982,n22007,n21980 );
   nor U21528 ( n21980,p2_reg1_reg_17_,n21998 );
   not U21529 ( n22007,n22008 );
   and U21530 ( n21982,n21998,p2_reg1_reg_17_ );
   not U21531 ( n21998,n21992 );
   nor U21532 ( n21986,n21992,n21957 );
   nand U21533 ( n21984,n21958,p2_addr_reg_17_ );
   nand U21534 ( n21983,p2_reg3_reg_17_,p2_u3088 );
   nand U21535 ( p2_u3230,n22009,n22010,n22011 );
   nor U21536 ( n22011,n22012,n22013,n22014 );
   nor U21537 ( n22014,n22015,n21939 );
   nor U21538 ( n22015,n22016,n22017 );
   nor U21539 ( n22017,n21996,n21999 );
   nand U21540 ( n21999,n21995,n21993 );
   nor U21541 ( n22016,n22018,n21995 );
   nand U21542 ( n21995,n22019,n22020 );
   nand U21543 ( n22020,n22021,n21368 );
   or U21544 ( n22021,n22022,n22023 );
   nand U21545 ( n22019,n22022,n22023 );
   nor U21546 ( n22018,n22024,n21996 );
   nor U21547 ( n21996,n22025,p2_reg2_reg_16_ );
   not U21548 ( n22024,n21993 );
   nand U21549 ( n21993,n22025,p2_reg2_reg_16_ );
   nor U21550 ( n22013,n22026,n21949 );
   nor U21551 ( n22026,n22027,n22028 );
   nor U21552 ( n22028,n22006,n22008 );
   nand U21553 ( n22008,n22005,n22003 );
   nor U21554 ( n22027,n22029,n22005 );
   nand U21555 ( n22005,n22030,n22031 );
   nand U21556 ( n22031,n22032,n22033 );
   or U21557 ( n22032,n22034,n22023 );
   nand U21558 ( n22030,n22034,n22023 );
   nor U21559 ( n22029,n22035,n22006 );
   nor U21560 ( n22006,n22025,p2_reg1_reg_16_ );
   not U21561 ( n22035,n22003 );
   nand U21562 ( n22003,n22025,p2_reg1_reg_16_ );
   not U21563 ( n22025,n22036 );
   nor U21564 ( n22012,n22036,n21957 );
   nand U21565 ( n22010,n21958,p2_addr_reg_16_ );
   nand U21566 ( n22009,p2_reg3_reg_16_,p2_u3088 );
   nand U21567 ( p2_u3229,n22037,n22038,n22039,n22040 );
   nand U21568 ( n22040,n22041,n22042 );
   nand U21569 ( n22042,n22043,n21957,n22044 );
   nand U21570 ( n22044,n22045,n21969 );
   xor U21571 ( n22045,p2_reg2_reg_15_,n22022 );
   nand U21572 ( n22043,n22046,n21967 );
   xor U21573 ( n22046,p2_reg1_reg_15_,n22034 );
   nand U21574 ( n22039,n22047,n22023 );
   nand U21575 ( n22047,n22048,n22049 );
   nand U21576 ( n22049,n21967,n22050 );
   xor U21577 ( n22050,n22034,n22033 );
   not U21578 ( n22033,p2_reg1_reg_15_ );
   nand U21579 ( n22034,n22051,n22052 );
   nand U21580 ( n22052,n22053,n22054 );
   nand U21581 ( n22053,n22055,n22056 );
   or U21582 ( n22051,n22056,n22055 );
   nand U21583 ( n22048,n21969,n22057 );
   xor U21584 ( n22057,n22022,n21368 );
   not U21585 ( n21368,p2_reg2_reg_15_ );
   nand U21586 ( n22022,n22058,n22059 );
   nand U21587 ( n22059,n22060,n22061 );
   nand U21588 ( n22060,n22055,n22062 );
   or U21589 ( n22058,n22062,n22055 );
   nand U21590 ( n22038,n21958,p2_addr_reg_15_ );
   nand U21591 ( n22037,p2_reg3_reg_15_,p2_u3088 );
   nand U21592 ( p2_u3228,n22063,n22064,n22065,n22066 );
   nand U21593 ( n22066,n22067,n22068 );
   nand U21594 ( n22068,n22069,n22070 );
   nand U21595 ( n22070,n22071,n21967 );
   xor U21596 ( n22071,n22056,p2_reg1_reg_14_ );
   nand U21597 ( n22069,n22072,n21969 );
   xor U21598 ( n22072,n22062,p2_reg2_reg_14_ );
   nand U21599 ( n22065,n22055,n22073 );
   nand U21600 ( n22073,n22074,n21957,n22075 );
   nand U21601 ( n22075,n21969,n22076 );
   xor U21602 ( n22076,n22061,n22062 );
   nand U21603 ( n22062,n22077,n22078 );
   nand U21604 ( n22078,n22079,n22080 );
   nand U21605 ( n22079,n22081,n22082,n22083 );
   nand U21606 ( n22083,n22084,n22085 );
   nand U21607 ( n22077,n22086,n22084 );
   not U21608 ( n22061,p2_reg2_reg_14_ );
   nand U21609 ( n22074,n21967,n22087 );
   xor U21610 ( n22087,n22054,n22056 );
   nand U21611 ( n22056,n22088,n22089 );
   nand U21612 ( n22089,n22090,n22091 );
   nand U21613 ( n22090,n22092,n22093,n22094 );
   nand U21614 ( n22094,n22095,n22096 );
   nand U21615 ( n22088,n22097,n22095 );
   not U21616 ( n22054,p2_reg1_reg_14_ );
   nand U21617 ( n22064,n21958,p2_addr_reg_14_ );
   nand U21618 ( n22063,p2_reg3_reg_14_,p2_u3088 );
   nand U21619 ( p2_u3227,n22098,n22099,n22100 );
   nor U21620 ( n22100,n22101,n22102,n22103 );
   nor U21621 ( n22103,n21939,n22104,n22105 );
   nor U21622 ( n22105,n22106,n22107,n22108 );
   nor U21623 ( n22108,n22109,n22110 );
   xor U21624 ( n22106,n22111,n21315 );
   and U21625 ( n22104,n22084,n22081,n22112 );
   or U21626 ( n22081,n22111,n21315 );
   nor U21627 ( n22084,n22113,n22110 );
   not U21628 ( n22113,n22080 );
   nand U21629 ( n22080,n21315,n22111 );
   not U21630 ( n21315,p2_reg2_reg_13_ );
   nor U21631 ( n22102,n21949,n22114,n22115 );
   nor U21632 ( n22115,n22116,n22117,n22118 );
   nor U21633 ( n22118,n22119,n22120 );
   xor U21634 ( n22116,n22111,n22121 );
   and U21635 ( n22114,n22095,n22092,n22122 );
   or U21636 ( n22092,n22111,n22121 );
   nor U21637 ( n22095,n22123,n22120 );
   not U21638 ( n22123,n22091 );
   nand U21639 ( n22091,n22121,n22111 );
   not U21640 ( n22121,p2_reg1_reg_13_ );
   nor U21641 ( n22101,n22111,n21957 );
   nand U21642 ( n22099,n21958,p2_addr_reg_13_ );
   nand U21643 ( n22098,p2_reg3_reg_13_,p2_u3088 );
   nand U21644 ( p2_u3226,n22124,n22125,n22126 );
   nor U21645 ( n22126,n22127,n22128,n22129 );
   nor U21646 ( n22129,n22130,n21939 );
   nor U21647 ( n22130,n22131,n22132 );
   nor U21648 ( n22132,n22110,n22112 );
   nand U21649 ( n22112,n22109,n22082 );
   nor U21650 ( n22131,n22109,n22133 );
   nor U21651 ( n22133,n22107,n22110 );
   nor U21652 ( n22110,n22134,p2_reg2_reg_12_ );
   not U21653 ( n22107,n22082 );
   nand U21654 ( n22082,n22134,p2_reg2_reg_12_ );
   nor U21655 ( n22109,n22086,n22085 );
   nor U21656 ( n22086,n22135,n22136 );
   nor U21657 ( n22128,n22137,n21949 );
   nor U21658 ( n22137,n22138,n22139 );
   nor U21659 ( n22139,n22120,n22122 );
   nand U21660 ( n22122,n22119,n22093 );
   nor U21661 ( n22138,n22119,n22140 );
   nor U21662 ( n22140,n22117,n22120 );
   nor U21663 ( n22120,n22134,p2_reg1_reg_12_ );
   not U21664 ( n22117,n22093 );
   nand U21665 ( n22093,n22134,p2_reg1_reg_12_ );
   not U21666 ( n22134,n22141 );
   nor U21667 ( n22119,n22097,n22096 );
   nor U21668 ( n22097,n22142,n22143 );
   nor U21669 ( n22127,n22141,n21957 );
   nand U21670 ( n22125,n21958,p2_addr_reg_12_ );
   nand U21671 ( n22124,p2_reg3_reg_12_,p2_u3088 );
   nand U21672 ( p2_u3225,n22144,n22145,n22146 );
   nor U21673 ( n22146,n22147,n22148,n22149 );
   nor U21674 ( n22149,n21939,n22150 );
   xor U21675 ( n22150,n22135,n22151 );
   nor U21676 ( n22151,n22085,n22136 );
   nor U21677 ( n22136,n22152,p2_reg2_reg_11_ );
   nor U21678 ( n22085,n22153,n21269 );
   not U21679 ( n21269,p2_reg2_reg_11_ );
   and U21680 ( n22135,n22154,n22155 );
   nand U21681 ( n22155,n22156,n22157,n22158 );
   nand U21682 ( n22157,n22159,n21160 );
   nand U21683 ( n22154,n22160,n22161 );
   nand U21684 ( n22161,n22162,n21217 );
   nand U21685 ( n22160,n22163,n22164,n22165 );
   nand U21686 ( n22165,n22166,p2_reg2_reg_8_,n22156 );
   nor U21687 ( n22148,n21949,n22167 );
   xor U21688 ( n22167,n22142,n22168 );
   nor U21689 ( n22168,n22096,n22143 );
   nor U21690 ( n22143,n22152,p2_reg1_reg_11_ );
   and U21691 ( n22096,n22152,p2_reg1_reg_11_ );
   not U21692 ( n22152,n22153 );
   and U21693 ( n22142,n22169,n22170 );
   nand U21694 ( n22170,n22171,n22172,n22173 );
   nand U21695 ( n22172,n22159,n22174 );
   nand U21696 ( n22169,n22175,n22176 );
   or U21697 ( n22176,n22177,p2_reg1_reg_10_ );
   nand U21698 ( n22175,n22178,n22179,n22180 );
   nand U21699 ( n22180,n22171,p2_reg1_reg_8_,n22166 );
   nor U21700 ( n22147,n22153,n21957 );
   nand U21701 ( n22145,n21958,p2_addr_reg_11_ );
   nand U21702 ( n22144,p2_reg3_reg_11_,p2_u3088 );
   nand U21703 ( p2_u3224,n22181,n22182,n22183 );
   nor U21704 ( n22183,n22184,n22185,n22186 );
   nor U21705 ( n22186,n21939,n22187,n22188 );
   nor U21706 ( n22188,n22189,n22190,n22191 );
   nor U21707 ( n22191,n22192,n22193 );
   xor U21708 ( n22189,n22162,n21217 );
   not U21709 ( n21217,p2_reg2_reg_10_ );
   and U21710 ( n22187,n22156,n22163,n22194 );
   nand U21711 ( n22163,n22177,p2_reg2_reg_10_ );
   nor U21712 ( n22156,n22192,n22195 );
   nor U21713 ( n22195,n22177,p2_reg2_reg_10_ );
   nor U21714 ( n22185,n21949,n22196,n22197 );
   nor U21715 ( n22197,n22198,n22199,n22200 );
   nor U21716 ( n22200,n22201,n22202 );
   xor U21717 ( n22198,n22177,p2_reg1_reg_10_ );
   and U21718 ( n22196,n22171,n22178,n22203 );
   nand U21719 ( n22178,n22177,p2_reg1_reg_10_ );
   nor U21720 ( n22171,n22201,n22204 );
   nor U21721 ( n22204,n22177,p2_reg1_reg_10_ );
   nor U21722 ( n22184,n22162,n21957 );
   nand U21723 ( n22182,n21958,p2_addr_reg_10_ );
   nand U21724 ( n22181,p2_reg3_reg_10_,p2_u3088 );
   nand U21725 ( p2_u3223,n22205,n22206,n22207 );
   nor U21726 ( n22207,n22208,n22209,n22210 );
   nor U21727 ( n22210,n22211,n21939 );
   nor U21728 ( n22211,n22212,n22213 );
   nor U21729 ( n22213,n22192,n22194 );
   nand U21730 ( n22194,n22193,n22164 );
   nor U21731 ( n22212,n22193,n22214 );
   nor U21732 ( n22214,n22192,n22190 );
   not U21733 ( n22190,n22164 );
   nand U21734 ( n22164,n22215,p2_reg2_reg_9_ );
   nor U21735 ( n22192,p2_reg2_reg_9_,n22215 );
   and U21736 ( n22193,n22216,n22217 );
   nand U21737 ( n22217,p2_reg2_reg_8_,n22218 );
   or U21738 ( n22218,n22166,n22158 );
   nand U21739 ( n22216,n22158,n22166 );
   nor U21740 ( n22209,n22219,n21949 );
   nor U21741 ( n22219,n22220,n22221 );
   nor U21742 ( n22221,n22201,n22203 );
   nand U21743 ( n22203,n22202,n22179 );
   nor U21744 ( n22220,n22202,n22222 );
   nor U21745 ( n22222,n22201,n22199 );
   not U21746 ( n22199,n22179 );
   nand U21747 ( n22179,n22215,p2_reg1_reg_9_ );
   nor U21748 ( n22201,p2_reg1_reg_9_,n22215 );
   not U21749 ( n22215,n22223 );
   and U21750 ( n22202,n22224,n22225 );
   nand U21751 ( n22225,p2_reg1_reg_8_,n22226 );
   or U21752 ( n22226,n22166,n22173 );
   nand U21753 ( n22224,n22166,n22173 );
   nor U21754 ( n22208,n22223,n21957 );
   nand U21755 ( n22206,n21958,p2_addr_reg_9_ );
   nand U21756 ( n22205,p2_reg3_reg_9_,p2_u3088 );
   nand U21757 ( p2_u3222,n22227,n22228,n22229,n22230 );
   nand U21758 ( n22230,n22159,n22231 );
   nand U21759 ( n22231,n22232,n22233 );
   nand U21760 ( n22233,n21967,n22234 );
   xor U21761 ( n22234,n22173,p2_reg1_reg_8_ );
   nand U21762 ( n22232,n21969,n22235 );
   xor U21763 ( n22235,n22158,p2_reg2_reg_8_ );
   nand U21764 ( n22229,n22166,n22236 );
   nand U21765 ( n22236,n22237,n21957,n22238 );
   nand U21766 ( n22238,n22239,n21969 );
   xor U21767 ( n22239,n21160,n22158 );
   nor U21768 ( n22158,n22240,n22241 );
   nor U21769 ( n22240,n22242,n22243 );
   not U21770 ( n21160,p2_reg2_reg_8_ );
   nand U21771 ( n22237,n22244,n21967 );
   not U21772 ( n21967,n21949 );
   xor U21773 ( n22244,n22174,n22173 );
   nor U21774 ( n22173,n22245,n22246 );
   nor U21775 ( n22245,n22247,n22248 );
   not U21776 ( n22174,p2_reg1_reg_8_ );
   not U21777 ( n22166,n22159 );
   nand U21778 ( n22228,n21958,p2_addr_reg_8_ );
   nand U21779 ( n22227,p2_reg3_reg_8_,p2_u3088 );
   nand U21780 ( p2_u3221,n22249,n22250,n22251 );
   nor U21781 ( n22251,n22252,n22253,n22254 );
   nor U21782 ( n22254,n21939,n22255,n22256 );
   nor U21783 ( n22256,n22242,n22257 );
   xor U21784 ( n22257,n22258,n21123 );
   nand U21785 ( n22242,n22259,n22260 );
   or U21786 ( n22260,n22261,n22262 );
   nor U21787 ( n22255,n22262,n22243,n22263,n22241 );
   nor U21788 ( n22241,p2_reg2_reg_7_,n22264 );
   not U21789 ( n22263,n22265 );
   nor U21790 ( n22243,n22258,n21123 );
   not U21791 ( n21123,p2_reg2_reg_7_ );
   nor U21792 ( n22253,n21949,n22266,n22267 );
   nor U21793 ( n22267,n22247,n22268 );
   xor U21794 ( n22268,n22264,p2_reg1_reg_7_ );
   nand U21795 ( n22247,n22269,n22270 );
   or U21796 ( n22270,n22271,n22272 );
   nor U21797 ( n22266,n22272,n22248,n22273,n22246 );
   nor U21798 ( n22246,p2_reg1_reg_7_,n22264 );
   not U21799 ( n22273,n22274 );
   and U21800 ( n22248,n22264,p2_reg1_reg_7_ );
   not U21801 ( n22264,n22258 );
   nor U21802 ( n22252,n22258,n21957 );
   nand U21803 ( n22250,n21958,p2_addr_reg_7_ );
   nand U21804 ( n22249,p2_reg3_reg_7_,p2_u3088 );
   nand U21805 ( p2_u3220,n22275,n22276,n22277 );
   nor U21806 ( n22277,n22278,n22279,n22280 );
   nor U21807 ( n22280,n22281,n21939 );
   nor U21808 ( n22281,n22282,n22283 );
   nor U21809 ( n22283,n22262,n22265 );
   nand U21810 ( n22265,n22261,n22259 );
   nor U21811 ( n22282,n22284,n22261 );
   or U21812 ( n22261,n22285,n22286 );
   nor U21813 ( n22285,n22287,n22288 );
   nor U21814 ( n22284,n22262,n22289 );
   not U21815 ( n22289,n22259 );
   nand U21816 ( n22259,n22290,p2_reg2_reg_6_ );
   nor U21817 ( n22262,n22290,p2_reg2_reg_6_ );
   nor U21818 ( n22279,n22291,n21949 );
   nor U21819 ( n22291,n22292,n22293 );
   nor U21820 ( n22293,n22272,n22274 );
   nand U21821 ( n22274,n22271,n22269 );
   nor U21822 ( n22292,n22294,n22271 );
   or U21823 ( n22271,n22295,n22296 );
   nor U21824 ( n22295,n22297,n22298 );
   nor U21825 ( n22294,n22272,n22299 );
   not U21826 ( n22299,n22269 );
   nand U21827 ( n22269,n22290,p2_reg1_reg_6_ );
   nor U21828 ( n22272,n22290,p2_reg1_reg_6_ );
   nor U21829 ( n22278,n22300,n21957 );
   nand U21830 ( n22276,n21958,p2_addr_reg_6_ );
   nand U21831 ( n22275,p2_reg3_reg_6_,p2_u3088 );
   nand U21832 ( p2_u3219,n22301,n22302,n22303 );
   nor U21833 ( n22303,n22304,n22305,n22306 );
   nor U21834 ( n22306,n21939,n22307,n22308 );
   nor U21835 ( n22308,n22287,n22309 );
   xor U21836 ( n22309,n22310,n21054 );
   nand U21837 ( n22287,n22311,n22312 );
   or U21838 ( n22312,n22313,n22314 );
   nor U21839 ( n22307,n22314,n22288,n22315,n22286 );
   nor U21840 ( n22286,p2_reg2_reg_5_,n22316 );
   not U21841 ( n22315,n22317 );
   nor U21842 ( n22288,n22310,n21054 );
   not U21843 ( n21054,p2_reg2_reg_5_ );
   nor U21844 ( n22305,n21949,n22318,n22319 );
   nor U21845 ( n22319,n22297,n22320 );
   xor U21846 ( n22320,n22316,p2_reg1_reg_5_ );
   nand U21847 ( n22297,n22321,n22322 );
   or U21848 ( n22322,n22323,n22324 );
   nor U21849 ( n22318,n22324,n22298,n22325,n22296 );
   nor U21850 ( n22296,p2_reg1_reg_5_,n22316 );
   not U21851 ( n22325,n22326 );
   and U21852 ( n22298,n22316,p2_reg1_reg_5_ );
   not U21853 ( n22316,n22310 );
   nor U21854 ( n22304,n22310,n21957 );
   nand U21855 ( n22302,n21958,p2_addr_reg_5_ );
   nand U21856 ( n22301,p2_reg3_reg_5_,p2_u3088 );
   nand U21857 ( p2_u3218,n22327,n22328,n22329 );
   nor U21858 ( n22329,n22330,n22331,n22332 );
   nor U21859 ( n22332,n22333,n21939 );
   nor U21860 ( n22333,n22334,n22335 );
   nor U21861 ( n22335,n22314,n22317 );
   nand U21862 ( n22317,n22313,n22311 );
   nor U21863 ( n22334,n22313,n22336 );
   nor U21864 ( n22336,n22314,n22337 );
   not U21865 ( n22337,n22311 );
   nand U21866 ( n22311,n22338,p2_reg2_reg_4_ );
   nor U21867 ( n22314,n22338,p2_reg2_reg_4_ );
   nor U21868 ( n22313,n22339,n22340 );
   nor U21869 ( n22340,n22341,n22342 );
   nor U21870 ( n22331,n22343,n21949 );
   nor U21871 ( n22343,n22344,n22345 );
   nor U21872 ( n22345,n22324,n22326 );
   nand U21873 ( n22326,n22323,n22321 );
   nor U21874 ( n22344,n22323,n22346 );
   nor U21875 ( n22346,n22324,n22347 );
   not U21876 ( n22347,n22321 );
   nand U21877 ( n22321,n22338,p2_reg1_reg_4_ );
   nor U21878 ( n22324,n22338,p2_reg1_reg_4_ );
   not U21879 ( n22338,n22348 );
   nor U21880 ( n22323,n22349,n22350 );
   nor U21881 ( n22350,n22351,n22352 );
   nor U21882 ( n22330,n22348,n21957 );
   nand U21883 ( n22328,n21958,p2_addr_reg_4_ );
   nand U21884 ( n22327,p2_reg3_reg_4_,p2_u3088 );
   nand U21885 ( p2_u3217,n22353,n22354,n22355 );
   nor U21886 ( n22355,n22356,n22357,n22358 );
   nor U21887 ( n22358,n21939,n22359 );
   xor U21888 ( n22359,n22342,n22360 );
   nor U21889 ( n22360,n22339,n22341 );
   nor U21890 ( n22341,p2_reg2_reg_3_,n22361 );
   nor U21891 ( n22339,n22362,n21001 );
   not U21892 ( n21001,p2_reg2_reg_3_ );
   and U21893 ( n22342,n22363,n22364,n22365 );
   nand U21894 ( n22365,n22366,n22367 );
   not U21895 ( n22366,n22368 );
   nand U21896 ( n22363,n22369,n22367 );
   nor U21897 ( n22357,n21949,n22370 );
   xor U21898 ( n22370,n22352,n22371 );
   nor U21899 ( n22371,n22349,n22351 );
   nor U21900 ( n22351,p2_reg1_reg_3_,n22361 );
   and U21901 ( n22349,n22361,p2_reg1_reg_3_ );
   not U21902 ( n22361,n22362 );
   and U21903 ( n22352,n22372,n22373,n22374 );
   nand U21904 ( n22374,n22375,n22376 );
   not U21905 ( n22375,n22377 );
   nand U21906 ( n22372,n22378,n22376 );
   nor U21907 ( n22356,n22362,n21957 );
   nand U21908 ( n22354,n21958,p2_addr_reg_3_ );
   nand U21909 ( n22353,p2_reg3_reg_3_,p2_u3088 );
   nand U21910 ( p2_u3216,n22379,n22380,n22381 );
   nor U21911 ( n22381,n22382,n22383,n22384 );
   nor U21912 ( n22384,n21939,n22385,n22386 );
   nor U21913 ( n22386,n22387,n22388 );
   xor U21914 ( n22388,n22389,p2_reg2_reg_2_ );
   and U21915 ( n22385,n22387,n22367,n22364 );
   nand U21916 ( n22364,n22389,p2_reg2_reg_2_ );
   or U21917 ( n22367,n22389,p2_reg2_reg_2_ );
   nand U21918 ( n22387,n22390,n22368 );
   nand U21919 ( n22368,n22391,n22392 );
   nor U21920 ( n22383,n21949,n22393,n22394 );
   nor U21921 ( n22394,n22395,n22396 );
   xor U21922 ( n22396,n22389,p2_reg1_reg_2_ );
   and U21923 ( n22393,n22395,n22376,n22373 );
   nand U21924 ( n22373,n22389,p2_reg1_reg_2_ );
   or U21925 ( n22376,n22389,p2_reg1_reg_2_ );
   nand U21926 ( n22395,n22397,n22377 );
   nand U21927 ( n22377,n22398,n22399 );
   nor U21928 ( n22382,n22400,n21957 );
   nand U21929 ( n22380,n21958,p2_addr_reg_2_ );
   nand U21930 ( n22379,p2_reg3_reg_2_,p2_u3088 );
   nand U21931 ( p2_u3215,n22401,n22402,n22403 );
   nor U21932 ( n22403,n22404,n22405,n22406 );
   nor U21933 ( n22406,n22407,n21939 );
   xor U21934 ( n22407,n22391,n22408 );
   nand U21935 ( n22408,n22390,n22392 );
   nand U21936 ( n22392,n20928,n22409 );
   not U21937 ( n22390,n22369 );
   nor U21938 ( n22369,n22409,n20928 );
   not U21939 ( n20928,p2_reg2_reg_1_ );
   nor U21940 ( n22405,n22410,n21949 );
   xor U21941 ( n22410,n22398,n22411 );
   nand U21942 ( n22411,n22397,n22399 );
   nand U21943 ( n22399,n22412,n22409 );
   not U21944 ( n22397,n22378 );
   nor U21945 ( n22378,n22409,n22412 );
   not U21946 ( n22412,p2_reg1_reg_1_ );
   nor U21947 ( n22404,n22409,n21957 );
   nand U21948 ( n22402,n21958,p2_addr_reg_1_ );
   nand U21949 ( n22401,p2_reg3_reg_1_,p2_u3088 );
   nand U21950 ( p2_u3214,n22414,n22415,n22416 );
   nor U21951 ( n22416,n22417,n22418,n22419 );
   nor U21952 ( n22419,n21939,n22391,n20911 );
   nor U21953 ( n22418,n21949,n22398,n22420 );
   nor U21954 ( n22417,n22421,n20626 );
   nor U21955 ( n22421,n22422,n22413,n22423 );
   nor U21956 ( n22423,n22398,n21949 );
   nand U21957 ( n22424,n22425,n22426 );
   nand U21958 ( n22425,n21828,p2_u3947 );
   nor U21959 ( n22398,n20626,n22420 );
   not U21960 ( n22420,p2_reg1_reg_0_ );
   nor U21961 ( n22413,n21828,n22427 );
   nor U21962 ( n22422,n22391,n21939 );
   nor U21963 ( n21969,n20216,n22427,n20217 );
   and U21964 ( n22427,n19538,n22426 );
   nand U21965 ( n22426,n22428,n22429 );
   nand U21966 ( n22428,n20218,n22430 );
   nand U21967 ( n22430,n20141,n22431 );
   nand U21968 ( n22431,n22432,n21924,n21646,n22433 );
   nor U21969 ( n22433,n21052,n19739,n21759 );
   not U21970 ( n21759,n21929 );
   not U21971 ( n21052,n20608 );
   not U21972 ( n21646,n19818 );
   nand U21973 ( n19818,n21534,n20609 );
   nand U21974 ( n20609,n20167,n22434,n20139 );
   not U21975 ( n21534,n21348 );
   nand U21976 ( n21348,n20223,n21042 );
   nor U21977 ( n20223,n20969,n20607 );
   not U21978 ( n20607,n20600 );
   nand U21979 ( n20600,n22434,n20137,n20139 );
   not U21980 ( n20969,n21040 );
   nand U21981 ( n20218,n22435,p2_state_reg );
   nor U21982 ( n22391,n20626,n20911 );
   not U21983 ( n20911,p2_reg2_reg_0_ );
   nand U21984 ( n22415,n21958,p2_addr_reg_0_ );
   nand U21985 ( n22429,n22438,n22439,n22440 );
   nand U21986 ( n22439,n21921,n22441 );
   nand U21987 ( n22438,n22437,n22436 );
   nand U21988 ( n22414,p2_reg3_reg_0_,p2_u3088 );
   nand U21989 ( p2_u3213,n22442,n22443,n22444,n22445 );
   nor U21990 ( n22445,n22446,n22447,n22448 );
   nor U21991 ( n22448,n19944,n22449 );
   not U21992 ( n19944,n19584 );
   nor U21993 ( n22447,n19946,n22450 );
   not U21994 ( n19946,n20371 );
   and U21995 ( n22446,p2_u3088,p2_reg3_reg_15_ );
   nand U21996 ( n22444,n22451,n19590 );
   or U21997 ( n22443,n22452,n22453 );
   xor U21998 ( n22453,n22454,n22455 );
   xor U21999 ( n22455,n22456,n22457 );
   nand U22000 ( n22442,n21369,n22458 );
   nand U22001 ( p2_u3212,n22459,n22460,n22461,n22462 );
   nor U22002 ( n22462,n22463,n22464,n22465 );
   nor U22003 ( n22465,n19775,n22449 );
   nor U22004 ( n22464,n21656,n22450 );
   nor U22005 ( n22463,p2_state_reg,n22466 );
   nand U22006 ( n22461,n22451,n19557 );
   nand U22007 ( n22460,n22467,n22468,n22469 );
   nand U22008 ( n22468,n22470,n22471,n22472 );
   nand U22009 ( n22467,n22473,n22474 );
   nand U22010 ( n22474,n22471,n22475 );
   nand U22011 ( n22473,n22476,n22470 );
   nand U22012 ( n22470,n22477,n22478 );
   nand U22013 ( n22459,n22479,n22480 );
   nand U22014 ( p2_u3211,n22481,n22482,n22483,n22484 );
   nor U22015 ( n22484,n22485,n22486,n22487 );
   nor U22016 ( n22487,n20082,n22488 );
   nor U22017 ( n22486,n20060,n22449 );
   nor U22018 ( n22485,p2_state_reg,n22489 );
   nand U22019 ( n22483,n22490,n22458 );
   nand U22020 ( n22482,n22491,n22492,n22469 );
   or U22021 ( n22492,n22493,n22494 );
   xor U22022 ( n22493,n22495,n22496 );
   nand U22023 ( n22491,n22497,n22498,n22494 );
   nand U22024 ( n22481,n22499,n20061 );
   nand U22025 ( p2_u3210,n22500,n22501,n22502,n22503 );
   nor U22026 ( n22503,n22504,n22505,n22506 );
   nor U22027 ( n22506,n19906,n22449 );
   nor U22028 ( n22505,n19907,n22488 );
   nor U22029 ( n22504,p2_state_reg,n22507 );
   nand U22030 ( n22502,n22499,n20525 );
   not U22031 ( n20525,n19908 );
   or U22032 ( n22501,n22508,n22452 );
   xor U22033 ( n22508,n22509,n22510 );
   xor U22034 ( n22509,n22511,n22512 );
   nand U22035 ( n22500,n22513,n22458 );
   nand U22036 ( p2_u3209,n22514,n22515,n22516,n22517 );
   nor U22037 ( n22517,n22518,n22519 );
   nor U22038 ( n22519,n20958,n22488 );
   not U22039 ( n20958,n19629 );
   nor U22040 ( n22518,n20083,n22449 );
   nand U22041 ( n22516,n22499,n20297 );
   nand U22042 ( n22515,n22520,n22521,n22469 );
   or U22043 ( n22521,n22522,n22523 );
   xor U22044 ( n22522,n22524,n22525 );
   nand U22045 ( n22520,n22526,n22527,n22523 );
   nand U22046 ( n22514,p2_reg3_reg_2_,n22528 );
   nand U22047 ( p2_u3208,n22529,n22530,n22531,n22532 );
   nor U22048 ( n22532,n22533,n22534,n22535 );
   nor U22049 ( n22535,n19999,n22449 );
   nor U22050 ( n22534,n22536,n21239 );
   not U22051 ( n21239,n22537 );
   and U22052 ( n22533,p2_u3088,p2_reg3_reg_11_ );
   nand U22053 ( n22531,n22499,n20000 );
   not U22054 ( n20000,n21238 );
   nand U22055 ( n22530,n22469,n22538 );
   nand U22056 ( n22538,n22539,n22540 );
   nand U22057 ( n22540,n22541,n22542,n22543 );
   nand U22058 ( n22541,n22544,n22545 );
   nand U22059 ( n22539,n22544,n22545,n22546 );
   nand U22060 ( n22546,n22543,n22542 );
   nand U22061 ( n22543,n22547,n22548 );
   nand U22062 ( n22529,n22451,n19602 );
   nand U22063 ( p2_u3207,n22549,n22550,n22551,n22552 );
   nor U22064 ( n22552,n22553,n22554,n22555 );
   nor U22065 ( n22555,n19857,n22488 );
   nor U22066 ( n22554,n19858,n22450 );
   nor U22067 ( n22553,p2_state_reg,n22556 );
   nand U22068 ( n22551,n22557,n19563 );
   or U22069 ( n22550,n22558,n22452 );
   xor U22070 ( n22558,n22559,n22560 );
   xor U22071 ( n22559,n22561,n22562 );
   nand U22072 ( n22549,n21577,n22480 );
   nand U22073 ( p2_u3206,n22563,n22564,n22565,n22566 );
   nor U22074 ( n22566,n22567,n22568,n22569 );
   nor U22075 ( n22569,n19945,n22449 );
   not U22076 ( n19945,n19590 );
   nor U22077 ( n22568,n19999,n22488 );
   not U22078 ( n19999,n19596 );
   nor U22079 ( n22567,p2_state_reg,n22570 );
   nand U22080 ( n22565,n22499,n19973 );
   not U22081 ( n19973,n21300 );
   nand U22082 ( n22564,n22571,n22572,n22469 );
   nand U22083 ( n22572,n22573,n22574,n22575 );
   nand U22084 ( n22575,n22576,n22577 );
   nand U22085 ( n22571,n22578,n22579,n22576,n22577 );
   nand U22086 ( n22578,n22580,n22574 );
   not U22087 ( n22580,n22581 );
   nand U22088 ( n22563,n21301,n22458 );
   nand U22089 ( p2_u3205,n22582,n22583,n22584,n22585 );
   nor U22090 ( n22585,n22586,n22587,n22588 );
   nor U22091 ( n22588,n19857,n22449 );
   not U22092 ( n19857,n19569 );
   nor U22093 ( n22587,n19906,n22488 );
   not U22094 ( n19906,n19575 );
   nor U22095 ( n22586,p2_state_reg,n22589 );
   nand U22096 ( n22584,n22499,n19883 );
   not U22097 ( n19883,n21490 );
   nand U22098 ( n22583,n22590,n22469 );
   xor U22099 ( n22590,n22591,n22592 );
   nand U22100 ( n22592,n22593,n22594 );
   nand U22101 ( n22582,n22595,n22480 );
   nand U22102 ( p2_u3204,n22596,n22597,n22598,n22599 );
   nand U22103 ( n22599,p2_reg3_reg_0_,n22528 );
   nand U22104 ( n22598,n22469,n22600 );
   xor U22105 ( n22600,n22601,n22602 );
   nand U22106 ( n22602,n22603,n22604 );
   nand U22107 ( n22601,n22605,n19632 );
   nand U22108 ( n22597,n22499,n20135 );
   nand U22109 ( n22596,n22557,n19629 );
   nand U22110 ( p2_u3203,n22606,n22607,n22608,n22609 );
   nor U22111 ( n22609,n22610,n22611,n22612 );
   nor U22112 ( n22612,n20022,n22488 );
   nor U22113 ( n22611,n20021,n22449 );
   not U22114 ( n20021,n19602 );
   nor U22115 ( n22610,p2_state_reg,n22613 );
   nand U22116 ( n22608,n22499,n20414 );
   not U22117 ( n20414,n20023 );
   or U22118 ( n22607,n22614,n22452 );
   xor U22119 ( n22614,n22615,n22616 );
   xor U22120 ( n22616,n22617,n22618 );
   nand U22121 ( n22606,n21176,n22458 );
   nand U22122 ( p2_u3202,n22619,n22620,n22621,n22622 );
   nor U22123 ( n22622,n22623,n22624,n22625 );
   nor U22124 ( n22625,n20083,n22488 );
   not U22125 ( n20083,n19623 );
   nor U22126 ( n22624,n20082,n22449 );
   not U22127 ( n20082,n19617 );
   nor U22128 ( n22623,p2_state_reg,n22626 );
   nand U22129 ( n22621,n22499,n20318 );
   not U22130 ( n20318,n20084 );
   or U22131 ( n22620,n22627,n22452 );
   xor U22132 ( n22627,n22628,n22629 );
   xor U22133 ( n22629,n22630,n22631 );
   nand U22134 ( n22619,n21021,n22458 );
   nand U22135 ( p2_u3201,n22632,n22633,n22634,n22635 );
   nor U22136 ( n22635,n22636,n22637,n22638 );
   nor U22137 ( n22638,n19831,n22449 );
   not U22138 ( n19831,n19557 );
   nor U22139 ( n22637,n19833,n22450 );
   nor U22140 ( n22636,p2_state_reg,n22639 );
   nand U22141 ( n22634,n22451,n19563 );
   nand U22142 ( n22633,n22469,n22640 );
   xor U22143 ( n22640,n22641,n22642 );
   nand U22144 ( n22641,n22643,n22644 );
   nand U22145 ( n22632,n21619,n22480 );
   nand U22146 ( p2_u3200,n22645,n22646,n22647,n22648 );
   nor U22147 ( n22648,n22649,n22650,n22651 );
   nor U22148 ( n22651,n21421,n22450 );
   nor U22149 ( n22650,n22536,n21422 );
   and U22150 ( n22649,p2_u3088,p2_reg3_reg_17_ );
   nand U22151 ( n22647,n22451,n19584 );
   nand U22152 ( n22646,n22652,n22653,n22469 );
   nand U22153 ( n22653,n22654,n22655 );
   nand U22154 ( n22655,n22656,n22657 );
   nand U22155 ( n22652,n22658,n22659,n22656,n22657 );
   nand U22156 ( n22658,n22660,n22661 );
   nand U22157 ( n22645,n22557,n19578 );
   nand U22158 ( p2_u3199,n22662,n22663,n22664,n22665 );
   nor U22159 ( n22665,n22666,n22667,n22668 );
   nor U22160 ( n22668,n20983,n22488 );
   not U22161 ( n20983,n19620 );
   nor U22162 ( n22667,n21113,n22449 );
   nor U22163 ( n22666,p2_state_reg,n22669 );
   nand U22164 ( n22664,n21031,n22458 );
   nand U22165 ( n22663,n22469,n22670 );
   nand U22166 ( n22670,n22671,n22672,n22673 );
   nand U22167 ( n22673,n22674,n22675 );
   nand U22168 ( n22672,n22676,n22677,n22678 );
   not U22169 ( n22678,n22679 );
   nand U22170 ( n22671,n22680,n22679 );
   xor U22171 ( n22680,n22677,n22676 );
   nand U22172 ( n22662,n22499,n20072 );
   nand U22173 ( p2_u3198,n22681,n22682,n22683,n22684 );
   nor U22174 ( n22684,n22685,n22686,n22687 );
   nor U22175 ( n22687,n19907,n22449 );
   not U22176 ( n19907,n19581 );
   nor U22177 ( n22686,n22536,n21379 );
   nor U22178 ( n22685,p2_state_reg,n22688 );
   nand U22179 ( n22683,n22499,n19934 );
   not U22180 ( n19934,n21378 );
   nand U22181 ( n22682,n22689,n22690,n22469 );
   or U22182 ( n22690,n22691,n22692 );
   xor U22183 ( n22691,n22693,n22694 );
   nand U22184 ( n22689,n22659,n22661,n22692 );
   nand U22185 ( n22681,n22451,n19587 );
   nand U22186 ( p2_u3197,n22695,n22696,n22697,n22698 );
   nor U22187 ( n22698,n22699,n22700,n22701 );
   nor U22188 ( n22701,n19814,n22449 );
   nor U22189 ( n22700,n19816,n22450 );
   and U22190 ( n22699,p2_u3088,p2_reg3_reg_25_ );
   nand U22191 ( n22697,n22451,n19560 );
   nand U22192 ( n22696,n22469,n22702 );
   nand U22193 ( n22702,n22703,n22704,n22705 );
   or U22194 ( n22705,n22476,n22477 );
   nand U22195 ( n22704,n22477,n22706,n22707 );
   nand U22196 ( n22703,n22708,n22709 );
   xor U22197 ( n22708,n22706,n22477 );
   and U22198 ( n22477,n22644,n22710 );
   nand U22199 ( n22695,n21638,n22480 );
   nand U22200 ( p2_u3196,n22711,n22712,n22713,n22714 );
   nor U22201 ( n22714,n22715,n22716,n22717 );
   nor U22202 ( n22717,n22536,n21281 );
   nor U22203 ( n22716,n19985,n22450 );
   nor U22204 ( n22715,p2_state_reg,n22718 );
   nand U22205 ( n22713,n22451,n19599 );
   nand U22206 ( n22712,n22719,n22720,n22469 );
   nand U22207 ( n22720,n22579,n22574,n22581 );
   or U22208 ( n22719,n22721,n22581 );
   xor U22209 ( n22721,n22722,n22723 );
   nand U22210 ( n22711,n22557,n19593 );
   nand U22211 ( p2_u3195,n22724,n22725,n22726,n22727 );
   nor U22212 ( n22727,n22728,n22729,n22730 );
   nor U22213 ( n22730,n21525,n22450 );
   nor U22214 ( n22729,n21533,n22488 );
   not U22215 ( n21533,n19572 );
   nor U22216 ( n22728,p2_state_reg,n22731 );
   nand U22217 ( n22726,n22557,n19566 );
   nand U22218 ( n22725,n22732,n22733,n22469 );
   nand U22219 ( n22733,n22734,n22735 );
   nand U22220 ( n22735,n22736,n22737 );
   nand U22221 ( n22732,n22738,n22593,n22736,n22737 );
   nand U22222 ( n22738,n22591,n22594 );
   nand U22223 ( n22724,n21526,n22480 );
   nand U22224 ( p2_u3194,n22739,n22740,n22741,n22742 );
   nand U22225 ( n22742,n22499,n20338 );
   nor U22226 ( n22741,n22743,n22744 );
   and U22227 ( n22744,n22528,p2_reg3_reg_1_ );
   nand U22228 ( n22528,n22536,p2_state_reg );
   nor U22229 ( n22743,n22452,n22745 );
   xor U22230 ( n22745,n22746,n22747 );
   nand U22231 ( n22746,n22748,n22749 );
   nand U22232 ( n22740,n22557,n19626 );
   nand U22233 ( n22739,n22451,n19632 );
   nand U22234 ( p2_u3193,n22750,n22751,n22752,n22753 );
   nor U22235 ( n22753,n22754,n22755,n22756 );
   nor U22236 ( n22756,n20060,n22488 );
   not U22237 ( n20060,n19611 );
   nor U22238 ( n22755,n22536,n21140 );
   nor U22239 ( n22754,p2_state_reg,n22757 );
   nand U22240 ( n22752,n22499,n20038 );
   nand U22241 ( n22751,n22758,n22469 );
   xor U22242 ( n22758,n22759,n22760 );
   and U22243 ( n22759,n22761,n22762 );
   nand U22244 ( n22750,n22557,n19605 );
   nand U22245 ( p2_u3192,n22763,n22764,n22765,n22766 );
   nor U22246 ( n22766,n22767,n22768,n22769 );
   nor U22247 ( n22769,n19775,n22488 );
   not U22248 ( n19775,n19551 );
   and U22249 ( n22768,n22480,n21745 );
   nor U22250 ( n22767,p2_state_reg,n22770 );
   nand U22251 ( n22765,n22499,n20575 );
   nand U22252 ( n22764,n22771,n22772,n22469 );
   nand U22253 ( n22772,n22773,n22774 );
   nand U22254 ( n22774,n22775,n22776 );
   nand U22255 ( n22775,n22777,n22778 );
   nand U22256 ( n22771,n22779,n22780 );
   nand U22257 ( n22780,n22781,n22778 );
   not U22258 ( n22781,n22782 );
   not U22259 ( n22779,n22773 );
   nand U22260 ( n22773,n22783,n22784 );
   nand U22261 ( n22784,n14937,n22786 );
   nand U22262 ( n22786,n21834,n21837 );
   nand U22263 ( n21837,n19792,n20575 );
   not U22264 ( n20575,n19778 );
   nand U22265 ( n21834,n19778,n19548 );
   nand U22266 ( n22783,n22787,n22788 );
   nand U22267 ( n22787,n22789,n22790 );
   nand U22268 ( n22790,n22791,n19778 );
   nand U22269 ( n22791,n22605,n19548 );
   nand U22270 ( n22789,n21750,n22605 );
   nor U22271 ( n21750,n19778,n19792 );
   not U22272 ( n19792,n19548 );
   nand U22273 ( n19778,n22792,n22793,n21921 );
   nand U22274 ( n22793,n16576,n17683 );
   or U22275 ( n22792,n20853,n16576 );
   nand U22276 ( n22763,n22557,n19545 );
   nand U22277 ( n19545,n22794,n22795,n22796,n22797 );
   nand U22278 ( n22797,n22798,n21758 );
   nor U22279 ( n21758,n22799,n22800,n22770 );
   not U22280 ( n22770,p2_reg3_reg_28_ );
   nand U22281 ( n22796,p2_reg0_reg_29_,n21826 );
   nand U22282 ( n22795,p2_reg1_reg_29_,n21827 );
   nand U22283 ( n22794,p2_reg2_reg_29_,n21825 );
   nand U22284 ( p2_u3191,n22801,n22802,n22803,n22804 );
   nor U22285 ( n22804,n22805,n22806,n22807 );
   nor U22286 ( n22807,n22536,n21473 );
   nor U22287 ( n22806,n19892,n22450 );
   and U22288 ( n22805,p2_u3088,p2_reg3_reg_19_ );
   nand U22289 ( n22803,n22557,n19572 );
   nand U22290 ( n22802,n22469,n22808 );
   nand U22291 ( n22808,n22809,n22810,n22811 );
   nand U22292 ( n22811,n22812,n22813 );
   nand U22293 ( n22810,n22814,n22815,n22816 );
   nand U22294 ( n22809,n22817,n22818 );
   xor U22295 ( n22817,n22814,n22815 );
   nand U22296 ( n22801,n22451,n19578 );
   nand U22297 ( p2_u3190,n22819,n22820,n22821,n22822 );
   nor U22298 ( n22822,n22823,n22824,n22825 );
   nor U22299 ( n22825,p2_reg3_reg_3_,n22536 );
   nor U22300 ( n22824,p2_state_reg,n21002 );
   nor U22301 ( n22823,n20099,n22488 );
   not U22302 ( n20099,n19626 );
   nand U22303 ( n22821,n22557,n19620 );
   nand U22304 ( n22820,n22826,n22827,n22469 );
   nand U22305 ( n22827,n22828,n22829 );
   nand U22306 ( n22829,n22830,n22831 );
   nand U22307 ( n22826,n22832,n22526,n22830,n22831 );
   nand U22308 ( n22832,n22833,n22527 );
   not U22309 ( n22833,n22523 );
   nand U22310 ( n22819,n22499,n20100 );
   nand U22311 ( p2_u3189,n22834,n22835,n22836,n22837 );
   nor U22312 ( n22837,n22838,n22839,n22840 );
   nor U22313 ( n22840,n19984,n22449 );
   not U22314 ( n19984,n19599 );
   nor U22315 ( n22839,n22536,n21198 );
   not U22316 ( n21198,n22841 );
   nor U22317 ( n22838,p2_state_reg,n22842 );
   nand U22318 ( n22836,n22499,n20011 );
   nand U22319 ( n22835,n22469,n22843 );
   xor U22320 ( n22843,n22844,n22845 );
   and U22321 ( n22845,n22542,n22548 );
   nand U22322 ( n22834,n22451,n19605 );
   nand U22323 ( p2_u3188,n22846,n22847,n22848,n22849 );
   nor U22324 ( n22849,n22850,n22851,n22852 );
   nor U22325 ( n22852,n19815,n22449 );
   not U22326 ( n19815,n19560 );
   nor U22327 ( n22851,n21586,n22450 );
   nor U22328 ( n22850,p2_state_reg,n22853 );
   nand U22329 ( n22848,n22451,n19566 );
   or U22330 ( n22847,n22854,n22452 );
   xor U22331 ( n22854,n22855,n22856 );
   xor U22332 ( n22855,n22857,n22858 );
   nand U22333 ( n22846,n21587,n22480 );
   nand U22334 ( p2_u3187,n22859,n22860,n22861,n22862 );
   nor U22335 ( n22862,n22863,n22864,n22865 );
   nor U22336 ( n22865,n19958,n22450 );
   nor U22337 ( n22864,n22536,n21340 );
   not U22338 ( n21340,n22866 );
   not U22339 ( n22536,n22458 );
   nor U22340 ( n22863,p2_state_reg,n22867 );
   nand U22341 ( n22861,n22451,n19593 );
   nand U22342 ( n22860,n22868,n22469 );
   xor U22343 ( n22868,n22869,n22870 );
   nand U22344 ( n22870,n22871,n22872 );
   nand U22345 ( n22859,n22557,n19587 );
   nand U22346 ( p2_u3186,n22873,n22874,n22875,n22876 );
   nor U22347 ( n22876,n22877,n22878,n22879 );
   nor U22348 ( n22879,n19814,n22488 );
   not U22349 ( n19814,n19554 );
   nor U22350 ( n22878,n21698,n22450 );
   nor U22351 ( n22877,p2_state_reg,n22799 );
   nand U22352 ( n22875,n22557,n19548 );
   nand U22353 ( n19548,n22880,n22881,n22882,n22883 );
   nand U22354 ( n22883,n22798,n21745 );
   xor U22355 ( n21745,n22884,p2_reg3_reg_28_ );
   nor U22356 ( n22884,n22800,n22799 );
   nand U22357 ( n22882,p2_reg0_reg_28_,n21826 );
   nand U22358 ( n22881,p2_reg1_reg_28_,n21827 );
   nand U22359 ( n22880,p2_reg2_reg_28_,n21825 );
   nand U22360 ( n22874,n22469,n22885 );
   nand U22361 ( n22885,n22886,n22887 );
   nand U22362 ( n22887,n22888,n22777 );
   nand U22363 ( n22888,n22778,n22776 );
   not U22364 ( n22776,n22889 );
   nand U22365 ( n22886,n22782,n22778 );
   nand U22366 ( n22778,n22890,n22891 );
   nor U22367 ( n22782,n22777,n22889 );
   nor U22368 ( n22889,n22891,n22890 );
   xor U22369 ( n22890,n22788,n21698 );
   nand U22370 ( n21698,n22892,n22893,n21921 );
   nand U22371 ( n22893,n16576,n18763 );
   or U22372 ( n22892,n20843,n16576 );
   nand U22373 ( n22891,n22605,n19551 );
   nand U22374 ( n19551,n22894,n22895,n22896,n22897 );
   nand U22375 ( n22897,n22798,n21699 );
   nand U22376 ( n22896,p2_reg0_reg_27_,n21826 );
   nand U22377 ( n22895,p2_reg1_reg_27_,n21827 );
   nand U22378 ( n22894,p2_reg2_reg_27_,n21825 );
   nand U22379 ( n22777,n22471,n22898 );
   nand U22380 ( n22898,n22472,n22899 );
   nand U22381 ( n22899,n22710,n22644,n22478 );
   nand U22382 ( n22478,n22706,n22709 );
   not U22383 ( n22706,n22900 );
   nand U22384 ( n22644,n22605,n19560,n22901 );
   xor U22385 ( n22901,n22785,n19833 );
   nand U22386 ( n22710,n22902,n22643 );
   nand U22387 ( n22643,n22903,n22904 );
   nand U22388 ( n22904,n22605,n19560 );
   nand U22389 ( n19560,n22905,n22906,n22907,n22908 );
   nand U22390 ( n22908,n21619,n22798 );
   nor U22391 ( n21619,n22909,n22910 );
   and U22392 ( n22909,n22639,n22911 );
   nand U22393 ( n22911,p2_reg3_reg_23_,n22912 );
   nand U22394 ( n22907,p2_reg0_reg_24_,n21826 );
   nand U22395 ( n22906,p2_reg1_reg_24_,n21827 );
   nand U22396 ( n22905,p2_reg2_reg_24_,n21825 );
   xor U22397 ( n22903,n19833,n22788 );
   nand U22398 ( n19833,n22913,n22914,n21921 );
   nand U22399 ( n22914,n16576,n19197 );
   or U22400 ( n22913,n20818,n16576 );
   not U22401 ( n22902,n22642 );
   nand U22402 ( n22642,n22915,n22916 );
   nand U22403 ( n22916,n22856,n22917 );
   or U22404 ( n22917,n22858,n22857 );
   xor U22405 ( n22856,n22788,n21586 );
   nand U22406 ( n21586,n22918,n22919,n21921 );
   nand U22407 ( n22919,n16576,n19201 );
   or U22408 ( n22918,n20811,n16576 );
   nand U22409 ( n22915,n22857,n22858 );
   nand U22410 ( n22858,n22920,n22921 );
   nand U22411 ( n22921,n22922,n22562 );
   nand U22412 ( n22562,n22923,n22737 );
   nand U22413 ( n22737,n22924,n22925 );
   nand U22414 ( n22925,n22605,n19569 );
   xor U22415 ( n22924,n21525,n22788 );
   nand U22416 ( n22923,n22734,n22736 );
   nand U22417 ( n22736,n22605,n19569,n22926 );
   xor U22418 ( n22926,n22785,n21525 );
   nand U22419 ( n21525,n22927,n22928,n21921 );
   nand U22420 ( n22928,n16576,n19209 );
   or U22421 ( n22927,n20794,n16576 );
   nand U22422 ( n19569,n22929,n22930,n22931,n22932 );
   nand U22423 ( n22932,n22798,n21526 );
   xor U22424 ( n21526,n22731,n22933 );
   nand U22425 ( n22931,p2_reg0_reg_21_,n21826 );
   nand U22426 ( n22930,p2_reg1_reg_21_,n21827 );
   nand U22427 ( n22929,p2_reg2_reg_21_,n21825 );
   and U22428 ( n22734,n22594,n22934 );
   nand U22429 ( n22934,n22935,n22593 );
   nand U22430 ( n22593,n22936,n22937 );
   nand U22431 ( n22937,n22605,n19572 );
   not U22432 ( n22936,n22938 );
   not U22433 ( n22935,n22591 );
   nor U22434 ( n22591,n22812,n22939 );
   and U22435 ( n22939,n22813,n22940 );
   nand U22436 ( n22940,n22818,n22815 );
   not U22437 ( n22813,n22814 );
   nand U22438 ( n22814,n22941,n22942 );
   nand U22439 ( n22942,n22943,n22512 );
   nand U22440 ( n22512,n22944,n22657 );
   nand U22441 ( n22657,n22945,n22946 );
   nand U22442 ( n22946,n22605,n19581 );
   xor U22443 ( n22945,n21421,n22788 );
   nand U22444 ( n22944,n22654,n22656 );
   nand U22445 ( n22656,n22605,n19581,n22947 );
   xor U22446 ( n22947,n14937,n21421 );
   nand U22447 ( n21421,n22948,n22949,n22950 );
   nand U22448 ( n22950,n21918,n21992 );
   nand U22449 ( n21992,n22951,n22952,n22953 );
   nand U22450 ( n22952,n20760,n20873 );
   nand U22451 ( n22951,p2_ir_reg_17_,n20759,p2_ir_reg_31_ );
   nand U22452 ( n22949,n22954,n22955 );
   nand U22453 ( n22948,n22956,n19225 );
   nand U22454 ( n19581,n22957,n22958,n22959,n22960 );
   nand U22455 ( n22960,n22798,n22961 );
   not U22456 ( n22961,n21422 );
   xor U22457 ( n21422,p2_reg3_reg_17_,n22962 );
   nand U22458 ( n22959,p2_reg0_reg_17_,n21826 );
   nand U22459 ( n22958,p2_reg1_reg_17_,n21827 );
   nand U22460 ( n22957,p2_reg2_reg_17_,n21825 );
   and U22461 ( n22654,n22661,n22963 );
   nand U22462 ( n22963,n22692,n22659 );
   nand U22463 ( n22659,n22693,n22694 );
   not U22464 ( n22692,n22660 );
   nand U22465 ( n22660,n22964,n22965 );
   nand U22466 ( n22965,n22454,n22966 );
   or U22467 ( n22966,n22456,n22457 );
   xor U22468 ( n22454,n14937,n20371 );
   nand U22469 ( n20371,n22967,n22968,n22969 );
   nand U22470 ( n22969,n22041,n21918 );
   not U22471 ( n22041,n22023 );
   nand U22472 ( n22023,n22970,n22971,n22972 );
   nand U22473 ( n22971,n20743,n20873 );
   nand U22474 ( n22970,p2_ir_reg_15_,n20742,p2_ir_reg_31_ );
   nand U22475 ( n22968,n22954,n20744 );
   nand U22476 ( n22967,n22956,p1_datao_reg_15_ );
   nand U22477 ( n22964,n22456,n22457 );
   nand U22478 ( n22457,n22973,n22871 );
   nand U22479 ( n22871,n22974,n22975 );
   nand U22480 ( n22973,n22869,n22872 );
   or U22481 ( n22872,n22975,n22974 );
   xor U22482 ( n22974,n22788,n19958 );
   not U22483 ( n19958,n20389 );
   nand U22484 ( n20389,n22976,n22977,n22978 );
   nand U22485 ( n22978,n22055,n21918 );
   not U22486 ( n22055,n22067 );
   nand U22487 ( n22067,n22979,n22980 );
   or U22488 ( n22980,p2_ir_reg_14_,p2_ir_reg_31_ );
   nand U22489 ( n22979,p2_ir_reg_31_,n20733 );
   nand U22490 ( n20733,n20742,n22981 );
   nand U22491 ( n22981,p2_ir_reg_14_,n22982 );
   not U22492 ( n20742,n20741 );
   nand U22493 ( n22977,n22954,n20734 );
   nand U22494 ( n22976,n22956,p1_datao_reg_14_ );
   nand U22495 ( n22975,n22605,n19590 );
   nand U22496 ( n19590,n22983,n22984,n22985,n22986 );
   nand U22497 ( n22986,n22866,n22798 );
   nor U22498 ( n22866,n22987,n22988 );
   and U22499 ( n22987,n22867,n22989 );
   or U22500 ( n22989,n22570,n22990 );
   nand U22501 ( n22985,p2_reg0_reg_14_,n21826 );
   nand U22502 ( n22984,p2_reg1_reg_14_,n21827 );
   nand U22503 ( n22983,p2_reg2_reg_14_,n21825 );
   and U22504 ( n22869,n22576,n22991 );
   nand U22505 ( n22991,n22992,n22577 );
   nand U22506 ( n22577,n22993,n22994 );
   nand U22507 ( n22994,n22605,n19593 );
   xor U22508 ( n22993,n21300,n22788 );
   nand U22509 ( n22992,n22574,n22573 );
   nand U22510 ( n22573,n22581,n22579 );
   nand U22511 ( n22579,n22722,n22723 );
   nand U22512 ( n22581,n22995,n22996 );
   nand U22513 ( n22996,n22997,n22544 );
   not U22514 ( n22997,n22548 );
   nand U22515 ( n22548,n22998,n22999,n22605 );
   nand U22516 ( n22999,n21212,n22788 );
   nand U22517 ( n21212,n21197,n19602 );
   not U22518 ( n21197,n20011 );
   nand U22519 ( n22998,n14937,n21228 );
   nand U22520 ( n21228,n20011,n19602 );
   and U22521 ( n22995,n22545,n23000 );
   nand U22522 ( n23000,n22542,n22544,n22844 );
   not U22523 ( n22844,n22547 );
   nand U22524 ( n22547,n23001,n23002 );
   nand U22525 ( n23002,n23003,n22617 );
   nand U22526 ( n22617,n23004,n22762 );
   nand U22527 ( n22762,n23005,n23006 );
   nand U22528 ( n23006,n22605,n19608 );
   xor U22529 ( n23005,n22785,n20038 );
   nand U22530 ( n23004,n23007,n22761 );
   nand U22531 ( n22761,n22605,n19608,n23008 );
   xor U22532 ( n23008,n20038,n22788 );
   not U22533 ( n20038,n21139 );
   nand U22534 ( n21139,n23009,n23010,n23011 );
   nand U22535 ( n23011,n21918,n22159 );
   nand U22536 ( n22159,n23012,n23013 );
   or U22537 ( n23013,p2_ir_reg_31_,p2_ir_reg_8_ );
   nand U22538 ( n23012,p2_ir_reg_31_,n23014 );
   nand U22539 ( n23014,n20683,n20682 );
   nand U22540 ( n20682,p2_ir_reg_8_,n23015 );
   nand U22541 ( n23010,n22954,n23016 );
   not U22542 ( n23016,n20684 );
   nand U22543 ( n23009,n22956,n19259 );
   not U22544 ( n23007,n22760 );
   nand U22545 ( n22760,n23017,n23018 );
   nand U22546 ( n23018,n22675,n23019,n22498,n23020 );
   not U22547 ( n22675,n22677 );
   nand U22548 ( n23017,n23019,n23021 );
   nand U22549 ( n23021,n23022,n22497,n23023 );
   nand U22550 ( n23023,n22679,n22498,n22676 );
   or U22551 ( n23003,n22618,n22615 );
   nand U22552 ( n23001,n22615,n22618 );
   nand U22553 ( n22618,n22605,n19605 );
   nand U22554 ( n19605,n23024,n23025,n23026,n23027 );
   nand U22555 ( n23027,n22798,n21176 );
   xor U22556 ( n21176,n22613,n23028 );
   nand U22557 ( n23026,p2_reg0_reg_9_,n21826 );
   nand U22558 ( n23025,p2_reg1_reg_9_,n21827 );
   nand U22559 ( n23024,p2_reg2_reg_9_,n21825 );
   xor U22560 ( n22615,n20023,n22788 );
   nand U22561 ( n20023,n23029,n23030,n23031 );
   nand U22562 ( n23031,n21918,n22223 );
   nand U22563 ( n22223,n23032,n23033,n23034 );
   nand U22564 ( n23033,n20873,n20692 );
   nand U22565 ( n23032,p2_ir_reg_31_,n20683,p2_ir_reg_9_ );
   not U22566 ( n20683,n20691 );
   nand U22567 ( n23030,n22954,n23035 );
   not U22568 ( n23035,n20693 );
   nand U22569 ( n23029,n22956,n19253 );
   nand U22570 ( n22544,n23036,n23037 );
   nand U22571 ( n23037,n22605,n19599 );
   not U22572 ( n23036,n23038 );
   nand U22573 ( n22542,n23039,n23040 );
   nand U22574 ( n23040,n22605,n19602 );
   nand U22575 ( n19602,n23041,n23042,n23043,n23044 );
   nand U22576 ( n23044,n22841,n22798 );
   nor U22577 ( n22841,n23045,n23046 );
   and U22578 ( n23045,n22842,n23047 );
   nand U22579 ( n23047,p2_reg3_reg_9_,n23048 );
   not U22580 ( n23048,n23028 );
   nand U22581 ( n23043,p2_reg0_reg_10_,n21826 );
   nand U22582 ( n23042,p2_reg1_reg_10_,n21827 );
   nand U22583 ( n23041,p2_reg2_reg_10_,n21825 );
   xor U22584 ( n23039,n22785,n20011 );
   nand U22585 ( n20011,n23049,n23050,n23051 );
   nand U22586 ( n23051,n22177,n21918 );
   not U22587 ( n22177,n22162 );
   nand U22588 ( n22162,n23052,n23053 );
   or U22589 ( n23053,p2_ir_reg_10_,p2_ir_reg_31_ );
   nand U22590 ( n23052,p2_ir_reg_31_,n20699 );
   nand U22591 ( n20699,n20708,n23054 );
   nand U22592 ( n23054,p2_ir_reg_10_,n23034 );
   nand U22593 ( n23050,n22954,n20700 );
   nand U22594 ( n23049,n22956,p1_datao_reg_10_ );
   nand U22595 ( n22545,n22605,n19599,n23038 );
   xor U22596 ( n23038,n14937,n21238 );
   nand U22597 ( n21238,n23055,n23056,n23057 );
   nand U22598 ( n23057,n21918,n22153 );
   nand U22599 ( n22153,n23058,n23059,n23060 );
   nand U22600 ( n23059,n20709,n20873 );
   nand U22601 ( n23058,p2_ir_reg_11_,n20708,p2_ir_reg_31_ );
   not U22602 ( n20708,n20707 );
   nand U22603 ( n23056,n22954,n23061 );
   not U22604 ( n23061,n20710 );
   nand U22605 ( n23055,n22956,n19045 );
   not U22606 ( n19045,p1_datao_reg_11_ );
   nand U22607 ( n19599,n23062,n23063,n23064,n23065 );
   nand U22608 ( n23065,n22798,n22537 );
   xor U22609 ( n22537,p2_reg3_reg_11_,n23046 );
   nand U22610 ( n23064,p2_reg0_reg_11_,n21826 );
   nand U22611 ( n23063,p2_reg1_reg_11_,n21827 );
   nand U22612 ( n23062,p2_reg2_reg_11_,n21825 );
   or U22613 ( n22574,n22723,n22722 );
   xor U22614 ( n22722,n22788,n19985 );
   nand U22615 ( n19985,n23066,n23067,n23068 );
   nand U22616 ( n23068,n21918,n22141 );
   nand U22617 ( n22141,n23069,n23070 );
   or U22618 ( n23070,p2_ir_reg_12_,p2_ir_reg_31_ );
   nand U22619 ( n23069,p2_ir_reg_31_,n20716 );
   nand U22620 ( n20716,n20725,n23071 );
   nand U22621 ( n23071,p2_ir_reg_12_,n23060 );
   nand U22622 ( n23067,n22954,n23072 );
   not U22623 ( n23072,n20717 );
   nand U22624 ( n23066,n22956,n19245 );
   nand U22625 ( n22723,n22605,n19596 );
   nand U22626 ( n19596,n23073,n23074,n23075,n23076 );
   nand U22627 ( n23076,n23077,n22798 );
   not U22628 ( n23077,n21281 );
   nand U22629 ( n21281,n23078,n22990 );
   nand U22630 ( n23078,n22718,n23079 );
   nand U22631 ( n23079,p2_reg3_reg_11_,n23046 );
   not U22632 ( n22718,p2_reg3_reg_12_ );
   nand U22633 ( n23075,p2_reg0_reg_12_,n21826 );
   nand U22634 ( n23074,p2_reg1_reg_12_,n21827 );
   nand U22635 ( n23073,p2_reg2_reg_12_,n21825 );
   nand U22636 ( n22576,n22605,n19593,n23080 );
   xor U22637 ( n23080,n22785,n21300 );
   nand U22638 ( n21300,n23081,n23082,n23083 );
   nand U22639 ( n23083,n21918,n22111 );
   nand U22640 ( n22111,n23084,n23085,n22982 );
   nand U22641 ( n23085,n20726,n20873 );
   nand U22642 ( n23084,p2_ir_reg_13_,n20725,p2_ir_reg_31_ );
   not U22643 ( n20725,n20724 );
   nand U22644 ( n23082,n22954,n23086 );
   not U22645 ( n23086,n20727 );
   nand U22646 ( n23081,n22956,n19070 );
   nand U22647 ( n19593,n23087,n23088,n23089,n23090 );
   nand U22648 ( n23090,n22798,n21301 );
   xor U22649 ( n21301,n22570,n22990 );
   nand U22650 ( n23089,p2_reg0_reg_13_,n21826 );
   nand U22651 ( n23088,p2_reg1_reg_13_,n21827 );
   nand U22652 ( n23087,p2_reg2_reg_13_,n21825 );
   nand U22653 ( n22456,n22605,n19587 );
   nand U22654 ( n19587,n23091,n23092,n23093,n23094 );
   nand U22655 ( n23094,n22798,n21369 );
   xor U22656 ( n21369,p2_reg3_reg_15_,n22988 );
   nand U22657 ( n23093,p2_reg0_reg_15_,n21826 );
   nand U22658 ( n23092,p2_reg1_reg_15_,n21827 );
   nand U22659 ( n23091,p2_reg2_reg_15_,n21825 );
   or U22660 ( n22661,n22694,n22693 );
   xor U22661 ( n22693,n22788,n21378 );
   nand U22662 ( n21378,n23095,n23096,n23097 );
   nand U22663 ( n23097,n21918,n22036 );
   nand U22664 ( n22036,n23098,n23099 );
   or U22665 ( n23099,p2_ir_reg_16_,p2_ir_reg_31_ );
   nand U22666 ( n23098,p2_ir_reg_31_,n20750 );
   nand U22667 ( n20750,n20759,n23100 );
   nand U22668 ( n23100,p2_ir_reg_16_,n22972 );
   not U22669 ( n20759,n20758 );
   nand U22670 ( n23096,n22954,n23101 );
   nand U22671 ( n23095,n22956,n19229 );
   not U22672 ( n19229,p1_datao_reg_16_ );
   nand U22673 ( n22694,n22605,n19584 );
   nand U22674 ( n19584,n23102,n23103,n23104,n23105 );
   nand U22675 ( n23105,n23106,n22798 );
   not U22676 ( n23106,n21379 );
   nand U22677 ( n21379,n23107,n22962 );
   nand U22678 ( n23107,n22688,n23108 );
   nand U22679 ( n23108,p2_reg3_reg_15_,n22988 );
   not U22680 ( n22688,p2_reg3_reg_16_ );
   nand U22681 ( n23104,p2_reg0_reg_16_,n21826 );
   nand U22682 ( n23103,p2_reg1_reg_16_,n21827 );
   nand U22683 ( n23102,p2_reg2_reg_16_,n21825 );
   or U22684 ( n22943,n22511,n22510 );
   nand U22685 ( n22941,n22510,n22511 );
   nand U22686 ( n22511,n22605,n19578 );
   nand U22687 ( n19578,n23109,n23110,n23111,n23112 );
   nand U22688 ( n23112,n22513,n22798 );
   not U22689 ( n22513,n21453 );
   nand U22690 ( n21453,n23113,n23114 );
   nand U22691 ( n23113,n22507,n23115 );
   nand U22692 ( n23115,p2_reg3_reg_17_,n23116 );
   not U22693 ( n22507,p2_reg3_reg_18_ );
   nand U22694 ( n23111,p2_reg0_reg_18_,n21826 );
   nand U22695 ( n23110,p2_reg1_reg_18_,n21827 );
   nand U22696 ( n23109,p2_reg2_reg_18_,n21825 );
   xor U22697 ( n22510,n22788,n19908 );
   nand U22698 ( n19908,n23117,n23118,n23119 );
   nand U22699 ( n23119,n21918,n21963 );
   nand U22700 ( n21963,n23120,n23121 );
   or U22701 ( n23121,p2_ir_reg_18_,p2_ir_reg_31_ );
   nand U22702 ( n23120,p2_ir_reg_31_,n20767 );
   nand U22703 ( n20767,n20776,n23122 );
   nand U22704 ( n23122,p2_ir_reg_18_,n22953 );
   nand U22705 ( n23118,n22954,n23123 );
   nand U22706 ( n23117,n22956,n19221 );
   nor U22707 ( n22812,n22815,n22818 );
   not U22708 ( n22818,n22816 );
   xor U22709 ( n22816,n22785,n19892 );
   nand U22710 ( n19892,n23124,n23125,n23126 );
   nand U22711 ( n23126,n21918,n21948 );
   nand U22712 ( n23125,n22954,n23127 );
   not U22713 ( n23127,n20778 );
   nand U22714 ( n23124,n22956,n19217 );
   nand U22715 ( n22815,n22605,n19575 );
   nand U22716 ( n19575,n23128,n23129,n23130,n23131 );
   nand U22717 ( n23131,n22798,n23132 );
   not U22718 ( n23132,n21473 );
   xor U22719 ( n21473,p2_reg3_reg_19_,n23114 );
   nand U22720 ( n23130,p2_reg0_reg_19_,n21826 );
   nand U22721 ( n23129,p2_reg1_reg_19_,n21827 );
   nand U22722 ( n23128,p2_reg2_reg_19_,n21825 );
   nand U22723 ( n22594,n22605,n19572,n22938 );
   xor U22724 ( n22938,n22785,n21490 );
   nand U22725 ( n21490,n23133,n23134,n21921 );
   nand U22726 ( n23134,n16576,n19213 );
   or U22727 ( n23133,n20785,n16576 );
   nand U22728 ( n19572,n23135,n23136,n23137,n23138 );
   nand U22729 ( n23138,n22595,n22798 );
   not U22730 ( n22595,n21491 );
   nand U22731 ( n21491,n23139,n22933 );
   nand U22732 ( n23139,n22589,n23140 );
   nand U22733 ( n23140,p2_reg3_reg_19_,n23141 );
   not U22734 ( n22589,p2_reg3_reg_20_ );
   nand U22735 ( n23137,p2_reg0_reg_20_,n21826 );
   nand U22736 ( n23136,p2_reg1_reg_20_,n21827 );
   nand U22737 ( n23135,p2_reg2_reg_20_,n21825 );
   or U22738 ( n22922,n22561,n22560 );
   nand U22739 ( n22920,n22560,n22561 );
   nand U22740 ( n22561,n22605,n19566 );
   nand U22741 ( n19566,n23142,n23143,n23144,n23145 );
   nand U22742 ( n23145,n21577,n22798 );
   and U22743 ( n21577,n23146,n23147 );
   nand U22744 ( n23146,n22556,n23148 );
   or U22745 ( n23148,n22731,n22933 );
   nand U22746 ( n23144,p2_reg0_reg_22_,n21826 );
   nand U22747 ( n23143,p2_reg1_reg_22_,n21827 );
   nand U22748 ( n23142,p2_reg2_reg_22_,n21825 );
   xor U22749 ( n22560,n22788,n19858 );
   nand U22750 ( n19858,n23149,n23150,n21921 );
   nand U22751 ( n23150,n16576,n19205 );
   or U22752 ( n23149,n20804,n16576 );
   nand U22753 ( n22857,n22605,n19563 );
   nand U22754 ( n19563,n23151,n23152,n23153,n23154 );
   nand U22755 ( n23154,n22798,n21587 );
   xor U22756 ( n21587,n22853,n23147 );
   nand U22757 ( n23153,p2_reg0_reg_23_,n21826 );
   nand U22758 ( n23152,p2_reg1_reg_23_,n21827 );
   nand U22759 ( n23151,p2_reg2_reg_23_,n21825 );
   and U22760 ( n22472,n22475,n22476 );
   nand U22761 ( n22476,n22707,n22900 );
   nand U22762 ( n22900,n22605,n19557 );
   nand U22763 ( n19557,n23155,n23156,n23157,n23158 );
   nand U22764 ( n23158,n22798,n21638 );
   xor U22765 ( n21638,p2_reg3_reg_25_,n22910 );
   nand U22766 ( n23157,p2_reg0_reg_25_,n21826 );
   nand U22767 ( n23156,p2_reg1_reg_25_,n21827 );
   nand U22768 ( n23155,p2_reg2_reg_25_,n21825 );
   not U22769 ( n22707,n22709 );
   xor U22770 ( n22709,n22785,n19816 );
   nand U22771 ( n19816,n23159,n23160,n21921 );
   nand U22772 ( n23160,n16576,n19193 );
   or U22773 ( n23159,n20827,n16576 );
   nand U22774 ( n22475,n23161,n23162 );
   nand U22775 ( n23162,n22605,n19554 );
   not U22776 ( n23161,n23163 );
   nand U22777 ( n22471,n22605,n19554,n23163 );
   xor U22778 ( n23163,n14937,n21656 );
   nand U22779 ( n21656,n23164,n23165,n21921 );
   nand U22780 ( n23165,n16576,n19189 );
   or U22781 ( n23164,n20834,n16576 );
   nand U22782 ( n19554,n23166,n23167,n23168,n23169 );
   nand U22783 ( n23169,n22479,n22798 );
   not U22784 ( n22479,n21657 );
   nand U22785 ( n21657,n22800,n23170 );
   nand U22786 ( n23170,n23171,n22466 );
   nand U22787 ( n23168,p2_reg0_reg_26_,n21826 );
   nand U22788 ( n23167,p2_reg1_reg_26_,n21827 );
   nand U22789 ( n23166,p2_reg2_reg_26_,n21825 );
   nand U22790 ( n22873,n21699,n22480 );
   nand U22791 ( n22480,n23172,n23173 );
   nand U22792 ( n23172,n23174,p2_state_reg );
   xor U22793 ( n21699,n22799,n22800 );
   or U22794 ( n22800,n22466,n23171 );
   nand U22795 ( n23171,p2_reg3_reg_25_,n22910 );
   nor U22796 ( n22910,n22853,n23147,n22639 );
   not U22797 ( n22639,p2_reg3_reg_24_ );
   not U22798 ( n23147,n22912 );
   nor U22799 ( n22912,n22731,n22933,n22556 );
   not U22800 ( n22556,p2_reg3_reg_22_ );
   nand U22801 ( n22933,p2_reg3_reg_19_,n23141,p2_reg3_reg_20_ );
   not U22802 ( n23141,n23114 );
   nand U22803 ( n23114,p2_reg3_reg_17_,n23116,p2_reg3_reg_18_ );
   not U22804 ( n23116,n22962 );
   nand U22805 ( n22962,p2_reg3_reg_15_,n22988,p2_reg3_reg_16_ );
   nor U22806 ( n22988,n22570,n22990,n22867 );
   not U22807 ( n22867,p2_reg3_reg_14_ );
   nand U22808 ( n22990,p2_reg3_reg_11_,n23046,p2_reg3_reg_12_ );
   nor U22809 ( n23046,n22842,n23028,n22613 );
   not U22810 ( n22613,p2_reg3_reg_9_ );
   not U22811 ( n22842,p2_reg3_reg_10_ );
   not U22812 ( n22570,p2_reg3_reg_13_ );
   not U22813 ( n22731,p2_reg3_reg_21_ );
   not U22814 ( n22853,p2_reg3_reg_23_ );
   not U22815 ( n22466,p2_reg3_reg_26_ );
   not U22816 ( n22799,p2_reg3_reg_27_ );
   nand U22817 ( p2_u3185,n23175,n23176,n23177,n23178 );
   nor U22818 ( n23178,n23179,n23180,n23181 );
   nor U22819 ( n23181,n21113,n22488 );
   nor U22820 ( n22451,n20215,n20216,n23182 );
   not U22821 ( n21113,n19614 );
   nor U22822 ( n23180,n20022,n22449 );
   nor U22823 ( n22557,n20215,n21828,n23182 );
   not U22824 ( n21828,n20216 );
   not U22825 ( n20022,n19608 );
   nand U22826 ( n19608,n23183,n23184,n23185,n23186 );
   nand U22827 ( n23186,n23187,n22798 );
   not U22828 ( n23187,n21140 );
   nand U22829 ( n21140,n23188,n23028 );
   nand U22830 ( n23028,p2_reg3_reg_7_,n23189,p2_reg3_reg_8_ );
   nand U22831 ( n23188,n22757,n23190 );
   nand U22832 ( n23190,p2_reg3_reg_7_,n23189 );
   not U22833 ( n23189,n23191 );
   not U22834 ( n22757,p2_reg3_reg_8_ );
   nand U22835 ( n23185,p2_reg0_reg_8_,n21826 );
   nand U22836 ( n23184,p2_reg1_reg_8_,n21827 );
   nand U22837 ( n23183,p2_reg2_reg_8_,n21825 );
   nor U22838 ( n23179,p2_state_reg,n23192 );
   nand U22839 ( n23177,n21103,n22458 );
   nand U22840 ( n22458,n23193,n23173 );
   nand U22841 ( n23173,n23194,p2_state_reg );
   nand U22842 ( n23194,n22436,n23195,n21932,n23196 );
   nand U22843 ( n21932,n20148,n20146 );
   not U22844 ( n20148,n22441 );
   nand U22845 ( n23195,n23197,n23182 );
   nand U22846 ( n23193,n23174,n20141 );
   and U22847 ( n23174,n23182,n23198 );
   nand U22848 ( n23198,n20215,n19777 );
   nand U22849 ( n20215,n20141,n20228,n20603 );
   nand U22850 ( n23176,n23199,n23200,n22469 );
   nand U22851 ( n22452,n20141,n23197,n23201 );
   nand U22852 ( n23197,n23202,n20314,n21924,n21043 );
   nand U22853 ( n21043,n20333,n20138 );
   nand U22854 ( n21924,n19741,n21948 );
   nand U22855 ( n20314,n21760,n20138 );
   nor U22856 ( n23202,n23203,n23204 );
   nor U22857 ( n23204,n20228,n20138 );
   nor U22858 ( n23203,n21820,n20145 );
   nand U22859 ( n23200,n23205,n22497,n23206 );
   nand U22860 ( n23206,n22494,n22498 );
   not U22861 ( n22494,n23207 );
   nand U22862 ( n23205,n23022,n23019 );
   nand U22863 ( n23199,n23208,n23022,n23019,n22498 );
   nand U22864 ( n22498,n22495,n22496 );
   nand U22865 ( n23019,n23209,n23210 );
   nand U22866 ( n23210,n22605,n19611 );
   xor U22867 ( n23209,n14937,n20049 );
   nand U22868 ( n23022,n22605,n19611,n23211 );
   xor U22869 ( n23211,n20049,n22788 );
   nand U22870 ( n19611,n23212,n23213,n23214,n23215 );
   nand U22871 ( n23215,n22798,n21103 );
   xor U22872 ( n21103,n23192,n23191 );
   not U22873 ( n23192,p2_reg3_reg_7_ );
   nand U22874 ( n23214,p2_reg0_reg_7_,n21826 );
   nand U22875 ( n23213,p2_reg1_reg_7_,n21827 );
   nand U22876 ( n23212,p2_reg2_reg_7_,n21825 );
   nand U22877 ( n23208,n23207,n22497 );
   or U22878 ( n22497,n22496,n22495 );
   xor U22879 ( n22495,n21066,n22788 );
   not U22880 ( n21066,n20061 );
   nand U22881 ( n20061,n23216,n23217,n23218 );
   nand U22882 ( n23218,n22290,n21918 );
   not U22883 ( n22290,n22300 );
   nand U22884 ( n22300,n23219,n23220 );
   or U22885 ( n23220,p2_ir_reg_31_,p2_ir_reg_6_ );
   nand U22886 ( n23219,p2_ir_reg_31_,n23221 );
   nand U22887 ( n23221,n20667,n20666 );
   nand U22888 ( n20666,p2_ir_reg_6_,n23222 );
   nand U22889 ( n23217,n22954,n20668 );
   nand U22890 ( n23216,n22956,p1_datao_reg_6_ );
   nand U22891 ( n22496,n19614,n22605 );
   nand U22892 ( n19614,n23223,n23224,n23225,n23226 );
   nand U22893 ( n23226,p2_reg0_reg_6_,n21826 );
   nand U22894 ( n23225,p2_reg1_reg_6_,n21827 );
   nand U22895 ( n23224,p2_reg2_reg_6_,n21825 );
   nand U22896 ( n23223,n22490,n22798 );
   not U22897 ( n22490,n21067 );
   nand U22898 ( n21067,n23227,n23191 );
   nand U22899 ( n23191,p2_reg3_reg_5_,n23228,p2_reg3_reg_6_ );
   nand U22900 ( n23227,n22489,n23229 );
   nand U22901 ( n23229,p2_reg3_reg_5_,n23228 );
   not U22902 ( n23228,n23230 );
   not U22903 ( n22489,p2_reg3_reg_6_ );
   nand U22904 ( n23207,n23020,n23231 );
   nand U22905 ( n23231,n23232,n22677 );
   nand U22906 ( n22677,n23233,n23234 );
   nand U22907 ( n23234,n23235,n22630 );
   nand U22908 ( n22630,n23236,n22831 );
   nand U22909 ( n22831,n23237,n23238 );
   nand U22910 ( n23238,n22605,n19623 );
   xor U22911 ( n23237,n22785,n20100 );
   nand U22912 ( n23236,n22828,n22830 );
   nand U22913 ( n22830,n22605,n19623,n23239 );
   xor U22914 ( n23239,n20100,n22788 );
   not U22915 ( n20100,n21015 );
   nand U22916 ( n21015,n23240,n23241,n23242 );
   nand U22917 ( n23242,n21918,n22362 );
   nand U22918 ( n22362,n23243,n23244,n23245 );
   nand U22919 ( n23244,n20873,n20644 );
   nand U22920 ( n23243,p2_ir_reg_31_,n20643,p2_ir_reg_3_ );
   nand U22921 ( n23241,n22954,n23246 );
   not U22922 ( n23246,n20645 );
   nand U22923 ( n23240,n22956,n19357 );
   nand U22924 ( n19623,n23247,n23248,n23249,n23250 );
   nand U22925 ( n23250,p2_reg0_reg_3_,n21826 );
   nand U22926 ( n23249,p2_reg1_reg_3_,n21827 );
   nand U22927 ( n23248,p2_reg2_reg_3_,n21825 );
   nand U22928 ( n23247,n22798,n21002 );
   and U22929 ( n22828,n22527,n23251 );
   nand U22930 ( n23251,n22526,n22523 );
   nand U22931 ( n22523,n22749,n23252 );
   nand U22932 ( n23252,n22747,n22748 );
   nand U22933 ( n22748,n23253,n23254 );
   nand U22934 ( n23254,n22605,n19629 );
   xor U22935 ( n23253,n20123,n22788 );
   nand U22936 ( n22747,n22604,n23255 );
   nand U22937 ( n23255,n22605,n19632,n22603 );
   or U22938 ( n22603,n23256,n22788 );
   nand U22939 ( n19632,n23257,n23258,n23259,n23260 );
   nand U22940 ( n23260,p2_reg0_reg_0_,n21826 );
   nand U22941 ( n23259,p2_reg1_reg_0_,n21827 );
   nand U22942 ( n23258,p2_reg2_reg_0_,n21825 );
   nand U22943 ( n23257,p2_reg3_reg_0_,n22798 );
   nand U22944 ( n22604,n23256,n22788 );
   xor U22945 ( n23256,n20135,n22788 );
   nand U22946 ( n20135,n23261,n23262,n23263 );
   nand U22947 ( n23263,p2_ir_reg_0_,n21918 );
   nand U22948 ( n23262,n20618,n22954 );
   nand U22949 ( n23261,n22956,p1_datao_reg_0_ );
   nand U22950 ( n22749,n22605,n19629,n23264 );
   xor U22951 ( n23264,n22785,n20123 );
   not U22952 ( n20123,n20338 );
   nand U22953 ( n20338,n23265,n23266,n23267 );
   or U22954 ( n23267,n22409,n21921 );
   nand U22955 ( n22409,n23268,n23269,n23270 );
   nand U22956 ( n23269,n20627,n20873 );
   nand U22957 ( n23268,p2_ir_reg_1_,p2_ir_reg_0_,p2_ir_reg_31_ );
   nand U22958 ( n23266,n22954,n20628 );
   nand U22959 ( n23265,n22956,p1_datao_reg_1_ );
   nand U22960 ( n19629,n23271,n23272,n23273,n23274 );
   nand U22961 ( n23274,p2_reg0_reg_1_,n21826 );
   nand U22962 ( n23273,p2_reg1_reg_1_,n21827 );
   nand U22963 ( n23272,p2_reg2_reg_1_,n21825 );
   nand U22964 ( n23271,p2_reg3_reg_1_,n22798 );
   nand U22965 ( n22526,n22524,n22525 );
   or U22966 ( n22527,n22525,n22524 );
   xor U22967 ( n22524,n20110,n22788 );
   not U22968 ( n20110,n20297 );
   nand U22969 ( n20297,n23275,n23276,n23277 );
   nand U22970 ( n23277,n22389,n21918 );
   not U22971 ( n22389,n22400 );
   nand U22972 ( n22400,n23278,n23279 );
   or U22973 ( n23279,p2_ir_reg_2_,p2_ir_reg_31_ );
   nand U22974 ( n23278,p2_ir_reg_31_,n20634 );
   nand U22975 ( n20634,n20643,n23280 );
   nand U22976 ( n23280,p2_ir_reg_2_,n23270 );
   not U22977 ( n20643,n20642 );
   nand U22978 ( n23276,n22954,n20635 );
   nand U22979 ( n23275,n22956,p1_datao_reg_2_ );
   nand U22980 ( n22525,n22605,n19626 );
   nand U22981 ( n19626,n23281,n23282,n23283,n23284 );
   nand U22982 ( n23284,p2_reg0_reg_2_,n21826 );
   nand U22983 ( n23283,p2_reg1_reg_2_,n21827 );
   nand U22984 ( n23282,p2_reg2_reg_2_,n21825 );
   nand U22985 ( n23281,p2_reg3_reg_2_,n22798 );
   or U22986 ( n23235,n22631,n22628 );
   nand U22987 ( n23233,n22628,n22631 );
   nand U22988 ( n22631,n22605,n19620 );
   nand U22989 ( n19620,n23285,n23286,n23287,n23288 );
   nand U22990 ( n23288,n21021,n22798 );
   and U22991 ( n21021,n23289,n23230 );
   nand U22992 ( n23289,n22626,n21002 );
   not U22993 ( n21002,p2_reg3_reg_3_ );
   not U22994 ( n22626,p2_reg3_reg_4_ );
   nand U22995 ( n23287,p2_reg0_reg_4_,n21826 );
   nand U22996 ( n23286,p2_reg1_reg_4_,n21827 );
   nand U22997 ( n23285,p2_reg2_reg_4_,n21825 );
   xor U22998 ( n22628,n20084,n22788 );
   nand U22999 ( n20084,n23290,n23291,n23292 );
   nand U23000 ( n23292,n21918,n22348 );
   nand U23001 ( n22348,n23293,n23294 );
   or U23002 ( n23294,p2_ir_reg_31_,p2_ir_reg_4_ );
   nand U23003 ( n23293,p2_ir_reg_31_,n23295 );
   nand U23004 ( n23295,n20651,n20650 );
   nand U23005 ( n20650,p2_ir_reg_4_,n23245 );
   nand U23006 ( n23291,n22954,n23296 );
   not U23007 ( n23296,n20652 );
   nand U23008 ( n23290,n22956,n19418 );
   not U23009 ( n19418,p1_datao_reg_4_ );
   nand U23010 ( n23232,n22676,n22679 );
   not U23011 ( n23020,n22674 );
   nor U23012 ( n22674,n22679,n22676 );
   and U23013 ( n22676,n22605,n19617 );
   nand U23014 ( n19617,n23297,n23298,n23299,n23300 );
   nand U23015 ( n23300,n22798,n21031 );
   xor U23016 ( n21031,n22669,n23230 );
   nand U23017 ( n23230,p2_reg3_reg_4_,p2_reg3_reg_3_ );
   not U23018 ( n22669,p2_reg3_reg_5_ );
   nand U23019 ( n23299,p2_reg0_reg_5_,n21826 );
   nand U23020 ( n23298,p2_reg1_reg_5_,n21827 );
   nand U23021 ( n23297,p2_reg2_reg_5_,n21825 );
   xor U23022 ( n23302,n20873,n20868 );
   not U23023 ( n20868,p2_ir_reg_30_ );
   not U23024 ( n23303,n23301 );
   nand U23025 ( n23301,n23304,n23305 );
   nand U23026 ( n23305,p2_ir_reg_29_,n20873 );
   nand U23027 ( n23304,p2_ir_reg_31_,n20858 );
   nand U23028 ( n20858,p2_ir_reg_29_,n20872 );
   nand U23029 ( n21042,n23307,n21948 );
   nor U23030 ( n23306,n20168,n23308 );
   not U23031 ( n23308,n20166 );
   nand U23032 ( n20166,n21948,n21820,n20167 );
   nor U23033 ( n22432,n21760,n20603,n20333 );
   nor U23034 ( n20333,n20146,n21820 );
   nor U23035 ( n20603,n20146,n20138 );
   nand U23036 ( n20146,n20137,n21948 );
   nor U23037 ( n21760,n20167,n21820,n21948 );
   xor U23038 ( n22679,n20072,n22788 );
   nor U23039 ( n23307,n20137,n21820 );
   nor U23040 ( n20168,n21948,n20228 );
   not U23041 ( n20072,n21030 );
   nand U23042 ( n21030,n23309,n23310,n23311 );
   nand U23043 ( n23311,n21918,n22310 );
   nand U23044 ( n22310,n23312,n23313,n23222 );
   nand U23045 ( n23313,n20873,n20660 );
   nand U23046 ( n23312,p2_ir_reg_31_,n20651,p2_ir_reg_5_ );
   not U23047 ( n20651,n20659 );
   nand U23048 ( n23310,n22954,n23314 );
   not U23049 ( n23314,n20661 );
   nand U23050 ( n23309,n22956,n19331 );
   nand U23051 ( n23175,n22499,n20049 );
   not U23052 ( n20049,n21102 );
   nand U23053 ( n21102,n23315,n23316,n23317 );
   nand U23054 ( n23317,n21918,n22258 );
   nand U23055 ( n22258,n23318,n23319,n23015 );
   nand U23056 ( n23319,n20873,n20676 );
   nand U23057 ( n23318,p2_ir_reg_31_,n20667,p2_ir_reg_7_ );
   not U23058 ( n20667,n20675 );
   nand U23059 ( n23316,n22954,n23320 );
   not U23060 ( n23320,n20677 );
   nand U23061 ( n23315,n22956,n19452 );
   not U23062 ( n19452,p1_datao_reg_7_ );
   not U23063 ( n22499,n22450 );
   nand U23064 ( n22450,n23321,n20141 );
   nor U23065 ( n20141,n22437,p2_u3088,n22435 );
   nand U23066 ( n23321,n21929,n23322 );
   nand U23067 ( n23322,n23201,n19739 );
   nand U23068 ( n20145,n20167,n20138 );
   not U23069 ( n20167,n20137 );
   not U23070 ( n23201,n23182 );
   nand U23071 ( n23182,n19731,n20144,n21931 );
   not U23072 ( n21931,n20143 );
   nand U23073 ( n20143,n20154,n23323 );
   or U23074 ( n23323,n20894,p2_d_reg_1_ );
   nand U23075 ( n20154,n23324,n23325 );
   nand U23076 ( n20144,n23326,n23327 );
   nand U23077 ( n23327,n23328,n23329,n23330,n23331 );
   nor U23078 ( n23331,n23332,n23333,n23334,n23335 );
   nand U23079 ( n23335,n20888,n20889,n20887 );
   not U23080 ( n20887,p2_d_reg_25_ );
   not U23081 ( n20889,p2_d_reg_27_ );
   not U23082 ( n20888,p2_d_reg_26_ );
   nand U23083 ( n23334,n20890,n20891,n20875,n20892 );
   not U23084 ( n20892,p2_d_reg_30_ );
   not U23085 ( n20875,p2_d_reg_2_ );
   not U23086 ( n20891,p2_d_reg_29_ );
   not U23087 ( n20890,p2_d_reg_28_ );
   nand U23088 ( n23333,n20893,n20876,n20877,n20878 );
   not U23089 ( n20878,p2_d_reg_5_ );
   not U23090 ( n20877,p2_d_reg_4_ );
   not U23091 ( n20876,p2_d_reg_3_ );
   not U23092 ( n20893,p2_d_reg_31_ );
   nand U23093 ( n23332,n20879,n20880,n20881,n20882 );
   not U23094 ( n20882,p2_d_reg_9_ );
   not U23095 ( n20881,p2_d_reg_8_ );
   not U23096 ( n20880,p2_d_reg_7_ );
   not U23097 ( n20879,p2_d_reg_6_ );
   nor U23098 ( n23330,n23336,p2_d_reg_10_,p2_d_reg_12_,p2_d_reg_11_ );
   nand U23099 ( n23336,n20883,n20884,n20885,n20886 );
   not U23100 ( n20886,p2_d_reg_16_ );
   not U23101 ( n20885,p2_d_reg_15_ );
   not U23102 ( n20884,p2_d_reg_14_ );
   not U23103 ( n20883,p2_d_reg_13_ );
   nor U23104 ( n23329,p2_d_reg_24_,p2_d_reg_23_,p2_d_reg_22_,p2_d_reg_21_ );
   nor U23105 ( n23328,p2_d_reg_20_,p2_d_reg_19_,p2_d_reg_18_,p2_d_reg_17_ );
   not U23106 ( n19731,n20140 );
   nand U23107 ( n20140,n20157,n23337 );
   or U23108 ( n23337,n20894,p2_d_reg_0_ );
   not U23109 ( n20894,n23326 );
   nor U23110 ( n23326,n23325,n23338 );
   and U23111 ( n23338,n23339,n23324 );
   xor U23112 ( n23339,n23340,p2_b_reg );
   nand U23113 ( n20157,n23341,n23325 );
   nand U23114 ( n21929,n20139,n19741 );
   not U23115 ( n19741,n19759 );
   nand U23116 ( n20137,n23342,n23343 );
   or U23117 ( n23343,p2_ir_reg_20_,p2_ir_reg_31_ );
   nand U23118 ( n23342,p2_ir_reg_31_,n23344 );
   nand U23119 ( n23344,n20784,n20783 );
   nand U23120 ( n20783,p2_ir_reg_20_,n23345 );
   nor U23121 ( n20149,n22434,n20228 );
   not U23122 ( n20139,n21948 );
   nand U23123 ( n21948,n23346,n23347,n23345 );
   nand U23124 ( n23347,n20777,n20873 );
   nand U23125 ( n23346,p2_ir_reg_19_,n20776,p2_ir_reg_31_ );
   not U23126 ( n20776,n20775 );
   nand U23127 ( p2_u3087,n22440,n23348 );
   nand U23128 ( n23348,n22441,n23196,n21921 );
   not U23129 ( n23196,n22437 );
   nor U23130 ( n22437,n23324,n23341,n23325 );
   nand U23131 ( n23325,n23349,n23350 );
   or U23132 ( n23350,p2_ir_reg_26_,p2_ir_reg_31_ );
   nand U23133 ( n23349,p2_ir_reg_31_,n23351 );
   nand U23134 ( n23351,n20833,n20832 );
   nand U23135 ( n20832,p2_ir_reg_26_,n23352 );
   nand U23136 ( n23352,n20825,n20826 );
   not U23137 ( n23341,n23340 );
   nand U23138 ( n23340,n23353,n23354 );
   nand U23139 ( n23354,n23355,n20816 );
   nand U23140 ( n20816,p2_ir_reg_24_,n20810 );
   nand U23141 ( n23353,p2_ir_reg_24_,n20873 );
   xor U23142 ( n23324,n20826,n23355 );
   nor U23143 ( n23355,n20873,n20825 );
   not U23144 ( n20826,p2_ir_reg_25_ );
   nand U23145 ( n22441,n22434,n20228 );
   not U23146 ( n20228,n21820 );
   nand U23147 ( n21820,n23356,n23357,n20802 );
   nand U23148 ( n23357,n20793,n20873 );
   nand U23149 ( n23356,p2_ir_reg_21_,n20784,p2_ir_reg_31_ );
   not U23150 ( n20784,n20792 );
   not U23151 ( n22434,n20138 );
   nand U23152 ( n20138,n23358,n23359,n23360 );
   nand U23153 ( n23359,n20803,n20873 );
   nand U23154 ( n23358,p2_ir_reg_22_,n20802,p2_ir_reg_31_ );
   and U23155 ( n22440,n23361,p2_state_reg );
   nand U23156 ( n23361,n22435,n21921 );
   nand U23157 ( n21921,n20216,n20217 );
   nand U23158 ( n20217,n23362,n23363,n20851 );
   nand U23159 ( n23363,n20842,n20873 );
   nand U23160 ( n23362,p2_ir_reg_27_,n20833,p2_ir_reg_31_ );
   not U23161 ( n20833,n20841 );
   nand U23162 ( n20216,n23364,n23365,n20872 );
   nand U23163 ( n20872,n20850,n20852 );
   not U23164 ( n20850,n20851 );
   nand U23165 ( n23365,n20852,n20873 );
   not U23166 ( n20873,p2_ir_reg_31_ );
   not U23167 ( n20852,p2_ir_reg_28_ );
   nand U23168 ( n23364,p2_ir_reg_28_,n20851,p2_ir_reg_31_ );
   nand U23169 ( n20851,n20841,n20842 );
   not U23170 ( n20842,p2_ir_reg_27_ );
   nor U23171 ( n20841,p2_ir_reg_25_,p2_ir_reg_26_,n20817 );
   not U23172 ( n20817,n20825 );
   nor U23173 ( n20825,n20810,p2_ir_reg_24_ );
   not U23174 ( n22435,n22436 );
   nand U23175 ( n22436,n23366,n23367 );
   or U23176 ( n23367,p2_ir_reg_23_,p2_ir_reg_31_ );
   nand U23177 ( n23366,p2_ir_reg_31_,n23368 );
   nand U23178 ( n23368,n20810,n20809 );
   nand U23179 ( n20809,p2_ir_reg_23_,n23360 );
   or U23180 ( n20810,n23360,p2_ir_reg_23_ );
   nand U23181 ( n23360,n20801,n20803 );
   not U23182 ( n20803,p2_ir_reg_22_ );
   not U23183 ( n20801,n20802 );
   nand U23184 ( n20802,n20792,n20793 );
   not U23185 ( n20793,p2_ir_reg_21_ );
   nor U23186 ( n20792,n23345,p2_ir_reg_20_ );
   nand U23187 ( n23345,n20775,n20777 );
   not U23188 ( n20777,p2_ir_reg_19_ );
   nor U23189 ( n20775,n22953,p2_ir_reg_18_ );
   nand U23190 ( n22953,n20758,n20760 );
   not U23191 ( n20760,p2_ir_reg_17_ );
   nor U23192 ( n20758,n22972,p2_ir_reg_16_ );
   nand U23193 ( n22972,n20741,n20743 );
   not U23194 ( n20743,p2_ir_reg_15_ );
   nor U23195 ( n20741,n22982,p2_ir_reg_14_ );
   nand U23196 ( n22982,n20724,n20726 );
   not U23197 ( n20726,p2_ir_reg_13_ );
   nor U23198 ( n20724,n23060,p2_ir_reg_12_ );
   nand U23199 ( n23060,n20707,n20709 );
   not U23200 ( n20709,p2_ir_reg_11_ );
   nor U23201 ( n20707,n23034,p2_ir_reg_10_ );
   nand U23202 ( n23034,n20691,n20692 );
   not U23203 ( n20692,p2_ir_reg_9_ );
   nor U23204 ( n20691,n23015,p2_ir_reg_8_ );
   nand U23205 ( n23015,n20675,n20676 );
   not U23206 ( n20676,p2_ir_reg_7_ );
   nor U23207 ( n20675,n23222,p2_ir_reg_6_ );
   nand U23208 ( n23222,n20659,n20660 );
   not U23209 ( n20660,p2_ir_reg_5_ );
   nor U23210 ( n20659,n23245,p2_ir_reg_4_ );
   nand U23211 ( n23245,n20642,n20644 );
   not U23212 ( n20644,p2_ir_reg_3_ );
   nor U23213 ( n20642,n23270,p2_ir_reg_2_ );
   nand U23214 ( n23270,n20626,n20627 );
   not U23215 ( n20627,p2_ir_reg_1_ );
   not U23216 ( n20626,p2_ir_reg_0_ );
   nand U23217 ( p1_u3591,n23369,n23370 );
   nand U23218 ( n23370,p1_datao_reg_31_,n23371 );
   nand U23219 ( n23369,p1_u4016,n23372 );
   nand U23220 ( p1_u3590,n23373,n23374 );
   nand U23221 ( n23374,p1_datao_reg_30_,n23371 );
   nand U23222 ( n23373,p1_u4016,n23375 );
   nand U23223 ( p1_u3589,n23376,n23377 );
   nand U23224 ( n23377,p1_datao_reg_29_,n23371 );
   nand U23225 ( n23376,p1_u4016,n23378 );
   nand U23226 ( p1_u3588,n23379,n23380 );
   nand U23227 ( n23380,p1_datao_reg_28_,n23371 );
   nand U23228 ( n23379,p1_u4016,n23381 );
   nand U23229 ( p1_u3587,n23382,n23383 );
   nand U23230 ( n23383,p1_datao_reg_27_,n23371 );
   nand U23231 ( n23382,p1_u4016,n23384 );
   nand U23232 ( p1_u3586,n23385,n23386 );
   nand U23233 ( n23386,p1_datao_reg_26_,n23371 );
   nand U23234 ( n23385,p1_u4016,n23387 );
   nand U23235 ( p1_u3585,n23388,n23389 );
   nand U23236 ( n23389,p1_datao_reg_25_,n23371 );
   nand U23237 ( n23388,p1_u4016,n23390 );
   nand U23238 ( p1_u3584,n23391,n23392 );
   nand U23239 ( n23392,p1_datao_reg_24_,n23371 );
   nand U23240 ( n23391,p1_u4016,n23393 );
   nand U23241 ( p1_u3583,n23394,n23395 );
   nand U23242 ( n23395,p1_datao_reg_23_,n23371 );
   nand U23243 ( n23394,p1_u4016,n23396 );
   nand U23244 ( p1_u3582,n23397,n23398 );
   nand U23245 ( n23398,p1_datao_reg_22_,n23371 );
   nand U23246 ( n23397,p1_u4016,n23399 );
   nand U23247 ( p1_u3581,n23400,n23401 );
   nand U23248 ( n23401,p1_datao_reg_21_,n23371 );
   nand U23249 ( n23400,p1_u4016,n23402 );
   nand U23250 ( p1_u3580,n23403,n23404 );
   nand U23251 ( n23404,p1_datao_reg_20_,n23371 );
   nand U23252 ( n23403,p1_u4016,n23405 );
   nand U23253 ( p1_u3579,n23406,n23407 );
   nand U23254 ( n23407,p1_datao_reg_19_,n23371 );
   nand U23255 ( n23406,p1_u4016,n23408 );
   nand U23256 ( p1_u3578,n23409,n23410 );
   nand U23257 ( n23410,p1_datao_reg_18_,n23371 );
   nand U23258 ( n23409,p1_u4016,n23411 );
   nand U23259 ( p1_u3577,n23412,n23413 );
   nand U23260 ( n23413,p1_datao_reg_17_,n23371 );
   nand U23261 ( n23412,p1_u4016,n23414 );
   nand U23262 ( p1_u3576,n23415,n23416 );
   nand U23263 ( n23416,p1_datao_reg_16_,n23371 );
   nand U23264 ( n23415,p1_u4016,n23417 );
   nand U23265 ( p1_u3575,n23418,n23419 );
   nand U23266 ( n23419,p1_datao_reg_15_,n23371 );
   nand U23267 ( n23418,p1_u4016,n23420 );
   nand U23268 ( p1_u3574,n23421,n23422 );
   nand U23269 ( n23422,p1_datao_reg_14_,n23371 );
   nand U23270 ( n23421,p1_u4016,n23423 );
   nand U23271 ( p1_u3573,n23424,n23425 );
   nand U23272 ( n23425,p1_datao_reg_13_,n23371 );
   nand U23273 ( n23424,p1_u4016,n23426 );
   nand U23274 ( p1_u3572,n23427,n23428 );
   nand U23275 ( n23428,p1_datao_reg_12_,n23371 );
   nand U23276 ( n23427,p1_u4016,n23429 );
   nand U23277 ( p1_u3571,n23430,n23431 );
   nand U23278 ( n23431,p1_datao_reg_11_,n23371 );
   nand U23279 ( n23430,p1_u4016,n23432 );
   nand U23280 ( p1_u3570,n23433,n23434 );
   nand U23281 ( n23434,p1_datao_reg_10_,n23371 );
   nand U23282 ( n23433,p1_u4016,n23435 );
   nand U23283 ( p1_u3569,n23436,n23437 );
   nand U23284 ( n23437,p1_datao_reg_9_,n23371 );
   nand U23285 ( n23436,p1_u4016,n23438 );
   nand U23286 ( p1_u3568,n23439,n23440 );
   nand U23287 ( n23440,p1_datao_reg_8_,n23371 );
   nand U23288 ( n23439,p1_u4016,n23441 );
   nand U23289 ( p1_u3567,n23442,n23443 );
   nand U23290 ( n23443,p1_datao_reg_7_,n23371 );
   nand U23291 ( n23442,p1_u4016,n23444 );
   nand U23292 ( p1_u3566,n23445,n23446 );
   nand U23293 ( n23446,p1_datao_reg_6_,n23371 );
   nand U23294 ( n23445,p1_u4016,n23447 );
   nand U23295 ( p1_u3565,n23448,n23449 );
   nand U23296 ( n23449,p1_datao_reg_5_,n23371 );
   nand U23297 ( n23448,p1_u4016,n23450 );
   nand U23298 ( p1_u3564,n23451,n23452 );
   nand U23299 ( n23452,p1_datao_reg_4_,n23371 );
   nand U23300 ( n23451,p1_u4016,n23453 );
   nand U23301 ( p1_u3563,n23454,n23455 );
   nand U23302 ( n23455,p1_datao_reg_3_,n23371 );
   nand U23303 ( n23454,p1_u4016,n23456 );
   nand U23304 ( p1_u3562,n23457,n23458 );
   nand U23305 ( n23458,p1_datao_reg_2_,n23371 );
   nand U23306 ( n23457,p1_u4016,n23459 );
   nand U23307 ( p1_u3561,n23460,n23461 );
   nand U23308 ( n23461,p1_datao_reg_1_,n23371 );
   nand U23309 ( n23460,p1_u4016,n23462 );
   nand U23310 ( p1_u3560,n23463,n23464 );
   nand U23311 ( n23464,p1_datao_reg_0_,n23371 );
   nand U23312 ( n23463,p1_u4016,n23465 );
   nand U23313 ( p1_u3559,n23466,n23467 );
   nand U23314 ( n23467,n23468,n23469 );
   nand U23315 ( n23466,p1_reg1_reg_31_,n23470 );
   nand U23316 ( p1_u3558,n23471,n23472 );
   nand U23317 ( n23472,p1_reg1_reg_30_,n23470 );
   nand U23318 ( n23471,n23468,n23473 );
   nand U23319 ( p1_u3557,n23474,n23475 );
   nand U23320 ( n23475,p1_reg1_reg_29_,n23470 );
   nand U23321 ( n23474,n23468,n23476 );
   nand U23322 ( p1_u3556,n23477,n23478 );
   nand U23323 ( n23478,p1_reg1_reg_28_,n23470 );
   nand U23324 ( n23477,n23468,n23479 );
   nand U23325 ( p1_u3555,n23480,n23481 );
   nand U23326 ( n23481,p1_reg1_reg_27_,n23470 );
   nand U23327 ( n23480,n23468,n23482 );
   nand U23328 ( p1_u3554,n23483,n23484 );
   nand U23329 ( n23484,p1_reg1_reg_26_,n23470 );
   nand U23330 ( n23483,n23468,n23485 );
   nand U23331 ( p1_u3553,n23486,n23487 );
   nand U23332 ( n23487,p1_reg1_reg_25_,n23470 );
   nand U23333 ( n23486,n23468,n23488 );
   nand U23334 ( p1_u3552,n23489,n23490 );
   nand U23335 ( n23490,p1_reg1_reg_24_,n23470 );
   nand U23336 ( n23489,n23468,n23491 );
   nand U23337 ( p1_u3551,n23492,n23493 );
   nand U23338 ( n23493,p1_reg1_reg_23_,n23470 );
   nand U23339 ( n23492,n23468,n23494 );
   nand U23340 ( p1_u3550,n23495,n23496 );
   nand U23341 ( n23496,p1_reg1_reg_22_,n23470 );
   nand U23342 ( n23495,n23468,n23497 );
   nand U23343 ( p1_u3549,n23498,n23499 );
   nand U23344 ( n23499,p1_reg1_reg_21_,n23470 );
   nand U23345 ( n23498,n23468,n23500 );
   nand U23346 ( p1_u3548,n23501,n23502 );
   nand U23347 ( n23502,p1_reg1_reg_20_,n23470 );
   nand U23348 ( n23501,n23468,n23503 );
   nand U23349 ( p1_u3547,n23504,n23505 );
   nand U23350 ( n23505,p1_reg1_reg_19_,n23470 );
   nand U23351 ( n23504,n23468,n23506 );
   nand U23352 ( p1_u3546,n23507,n23508 );
   nand U23353 ( n23508,p1_reg1_reg_18_,n23470 );
   nand U23354 ( n23507,n23468,n23509 );
   nand U23355 ( p1_u3545,n23510,n23511 );
   nand U23356 ( n23511,p1_reg1_reg_17_,n23470 );
   nand U23357 ( n23510,n23468,n23512 );
   nand U23358 ( p1_u3544,n23513,n23514 );
   nand U23359 ( n23514,p1_reg1_reg_16_,n23470 );
   nand U23360 ( n23513,n23468,n23515 );
   nand U23361 ( p1_u3543,n23516,n23517 );
   nand U23362 ( n23517,p1_reg1_reg_15_,n23470 );
   nand U23363 ( n23516,n23468,n23518 );
   nand U23364 ( p1_u3542,n23519,n23520 );
   nand U23365 ( n23520,p1_reg1_reg_14_,n23470 );
   nand U23366 ( n23519,n23468,n23521 );
   nand U23367 ( p1_u3541,n23522,n23523 );
   nand U23368 ( n23523,p1_reg1_reg_13_,n23470 );
   nand U23369 ( n23522,n23468,n23524 );
   nand U23370 ( p1_u3540,n23525,n23526 );
   nand U23371 ( n23526,p1_reg1_reg_12_,n23470 );
   nand U23372 ( n23525,n23468,n23527 );
   nand U23373 ( p1_u3539,n23528,n23529 );
   nand U23374 ( n23529,p1_reg1_reg_11_,n23470 );
   nand U23375 ( n23528,n23468,n23530 );
   nand U23376 ( p1_u3538,n23531,n23532 );
   nand U23377 ( n23532,p1_reg1_reg_10_,n23470 );
   nand U23378 ( n23531,n23468,n23533 );
   nand U23379 ( p1_u3537,n23534,n23535 );
   nand U23380 ( n23535,p1_reg1_reg_9_,n23470 );
   nand U23381 ( n23534,n23468,n23536 );
   nand U23382 ( p1_u3536,n23537,n23538 );
   nand U23383 ( n23538,p1_reg1_reg_8_,n23470 );
   nand U23384 ( n23537,n23468,n23539 );
   nand U23385 ( p1_u3535,n23540,n23541 );
   nand U23386 ( n23541,p1_reg1_reg_7_,n23470 );
   nand U23387 ( n23540,n23468,n23542 );
   nand U23388 ( p1_u3534,n23543,n23544 );
   nand U23389 ( n23544,p1_reg1_reg_6_,n23470 );
   nand U23390 ( n23543,n23468,n23545 );
   nand U23391 ( p1_u3533,n23546,n23547 );
   nand U23392 ( n23547,p1_reg1_reg_5_,n23470 );
   nand U23393 ( n23546,n23468,n23548 );
   nand U23394 ( p1_u3532,n23549,n23550 );
   nand U23395 ( n23550,p1_reg1_reg_4_,n23470 );
   nand U23396 ( n23549,n23468,n23551 );
   nand U23397 ( p1_u3531,n23552,n23553 );
   nand U23398 ( n23553,p1_reg1_reg_3_,n23470 );
   nand U23399 ( n23552,n23468,n23554 );
   nand U23400 ( p1_u3530,n23555,n23556 );
   nand U23401 ( n23556,p1_reg1_reg_2_,n23470 );
   nand U23402 ( n23555,n23468,n23557 );
   nand U23403 ( p1_u3529,n23558,n23559 );
   nand U23404 ( n23559,p1_reg1_reg_1_,n23470 );
   nand U23405 ( n23558,n23468,n23560 );
   nand U23406 ( p1_u3528,n23561,n23562 );
   nand U23407 ( n23562,p1_reg1_reg_0_,n23470 );
   nand U23408 ( n23561,n23468,n23563 );
   nand U23409 ( p1_u3527,n23567,n23568 );
   nand U23410 ( n23568,n23569,n23469 );
   nand U23411 ( n23469,n23570,n23571,n23572 );
   nand U23412 ( n23572,n23573,n23574 );
   nand U23413 ( n23570,n23575,n23576 );
   nand U23414 ( n23567,p1_reg0_reg_31_,n23577 );
   nand U23415 ( p1_u3526,n23578,n23579 );
   nand U23416 ( n23579,n23569,n23473 );
   nand U23417 ( n23473,n23580,n23571,n23581 );
   nand U23418 ( n23581,n23582,n23573 );
   nand U23419 ( n23580,n23583,n23584,n23575 );
   nand U23420 ( n23578,p1_reg0_reg_30_,n23577 );
   nand U23421 ( p1_u3525,n23585,n23586 );
   nand U23422 ( n23586,n23569,n23476 );
   nand U23423 ( n23476,n23587,n23588,n23589,n23590 );
   nand U23424 ( n23590,n23591,n23592 );
   nand U23425 ( n23589,n23575,n23593 );
   nand U23426 ( n23588,n23594,n23573 );
   not U23427 ( n23587,n23595 );
   nand U23428 ( n23585,p1_reg0_reg_29_,n23577 );
   nand U23429 ( p1_u3524,n23596,n23597 );
   nand U23430 ( n23597,n23569,n23479 );
   nand U23431 ( n23479,n23598,n23599,n23600,n23601 );
   nor U23432 ( n23601,n23602,n23603,n23604 );
   nor U23433 ( n23604,n23605,n23606 );
   nor U23434 ( n23603,n23607,n23608 );
   nand U23435 ( n23600,n23609,n23573 );
   nand U23436 ( n23599,n23610,n23611,n23575 );
   nand U23437 ( n23598,n23612,n23591 );
   nand U23438 ( n23596,p1_reg0_reg_28_,n23577 );
   nand U23439 ( p1_u3523,n23613,n23614 );
   nand U23440 ( n23614,n23569,n23482 );
   nand U23441 ( n23482,n23615,n23616,n23617 );
   nor U23442 ( n23617,n23618,n23619,n23620 );
   nor U23443 ( n23620,n23621,n23622 );
   and U23444 ( n23619,n23623,n23575 );
   nor U23445 ( n23618,n23624,n23625 );
   nand U23446 ( n23616,n23626,n23381 );
   nand U23447 ( n23613,p1_reg0_reg_27_,n23577 );
   nand U23448 ( p1_u3522,n23627,n23628 );
   nand U23449 ( n23628,n23569,n23485 );
   nand U23450 ( n23485,n23629,n23630,n23631 );
   nor U23451 ( n23631,n23632,n23633,n23634 );
   nor U23452 ( n23634,n23621,n23635 );
   and U23453 ( n23633,n23575,n23636,n23637 );
   nor U23454 ( n23632,n23624,n23638 );
   nand U23455 ( n23630,n23626,n23384 );
   nand U23456 ( n23627,p1_reg0_reg_26_,n23577 );
   nand U23457 ( p1_u3521,n23639,n23640 );
   nand U23458 ( n23640,n23569,n23488 );
   nand U23459 ( n23488,n23641,n23642,n23643,n23644 );
   nor U23460 ( n23644,n23645,n23646,n23647 );
   nor U23461 ( n23647,n23648,n23608 );
   nor U23462 ( n23646,n23624,n23649 );
   nor U23463 ( n23645,n23650,n23606 );
   nand U23464 ( n23643,n23651,n23652 );
   nand U23465 ( n23642,n23575,n23653 );
   nand U23466 ( n23641,n23654,n23655 );
   nand U23467 ( n23639,p1_reg0_reg_25_,n23577 );
   nand U23468 ( p1_u3520,n23656,n23657 );
   nand U23469 ( n23657,n23569,n23491 );
   nand U23470 ( n23491,n23658,n23659,n23660,n23661 );
   nor U23471 ( n23661,n23662,n23663,n23664 );
   nor U23472 ( n23664,n23665,n23608 );
   nor U23473 ( n23663,n23624,n23666 );
   nor U23474 ( n23662,n23667,n23606 );
   nand U23475 ( n23660,n23668,n23652 );
   nand U23476 ( n23659,n23669,n23670,n23575 );
   nand U23477 ( n23658,n23671,n23655 );
   nand U23478 ( n23656,p1_reg0_reg_24_,n23577 );
   nand U23479 ( p1_u3519,n23672,n23673 );
   nand U23480 ( n23673,n23569,n23494 );
   nand U23481 ( n23494,n23674,n23675,n23676 );
   nor U23482 ( n23676,n23677,n23678,n23679 );
   nor U23483 ( n23679,n23680,n23621 );
   and U23484 ( n23678,n23681,n23575 );
   nor U23485 ( n23677,n23624,n23682 );
   nand U23486 ( n23675,n23626,n23393 );
   nand U23487 ( n23672,p1_reg0_reg_23_,n23577 );
   nand U23488 ( p1_u3518,n23683,n23684 );
   nand U23489 ( n23684,n23569,n23497 );
   nand U23490 ( n23497,n23685,n23686,n23687,n23688 );
   nor U23491 ( n23688,n23689,n23690,n23691 );
   nor U23492 ( n23691,n23692,n23608 );
   nor U23493 ( n23690,n23624,n23693 );
   nor U23494 ( n23689,n23665,n23606 );
   nand U23495 ( n23687,n23694,n23655 );
   nand U23496 ( n23685,n23695,n23696,n23575 );
   nand U23497 ( n23683,p1_reg0_reg_22_,n23577 );
   nand U23498 ( p1_u3517,n23697,n23698 );
   nand U23499 ( n23698,n23569,n23500 );
   nand U23500 ( n23500,n23699,n23700,n23701 );
   nor U23501 ( n23701,n23702,n23703,n23704 );
   nor U23502 ( n23704,n23621,n23705 );
   and U23503 ( n23703,n23706,n23575 );
   nor U23504 ( n23702,n23624,n23707 );
   nand U23505 ( n23700,n23626,n23399 );
   nand U23506 ( n23697,p1_reg0_reg_21_,n23577 );
   nand U23507 ( p1_u3516,n23708,n23709 );
   nand U23508 ( n23709,n23569,n23503 );
   nand U23509 ( n23503,n23710,n23711,n23712 );
   nor U23510 ( n23712,n23713,n23714,n23715 );
   nor U23511 ( n23715,n23621,n23716 );
   and U23512 ( n23714,n23575,n23717,n23718 );
   nor U23513 ( n23713,n23624,n23719 );
   nand U23514 ( n23711,n23626,n23402 );
   nand U23515 ( n23708,p1_reg0_reg_20_,n23577 );
   nand U23516 ( p1_u3515,n23720,n23721 );
   nand U23517 ( n23721,n23569,n23506 );
   nand U23518 ( n23506,n23722,n23723,n23724,n23725 );
   nor U23519 ( n23725,n23726,n23727 );
   nor U23520 ( n23726,n23728,n23606 );
   nand U23521 ( n23724,n23729,n23573 );
   nand U23522 ( n23723,n23575,n23730 );
   nand U23523 ( n23722,n23731,n23591 );
   nand U23524 ( n23720,p1_reg0_reg_19_,n23577 );
   nand U23525 ( p1_u3513,n23732,n23733 );
   nand U23526 ( n23733,n23569,n23509 );
   nand U23527 ( n23509,n23734,n23735,n23736,n23737 );
   nor U23528 ( n23737,n23738,n23739,n23740 );
   nor U23529 ( n23740,n23741,n23608 );
   nor U23530 ( n23739,n23742,n23743 );
   nor U23531 ( n23738,n23744,n23606 );
   nand U23532 ( n23736,n23745,n23573 );
   nand U23533 ( n23735,n23746,n23655 );
   or U23534 ( n23734,n23747,n23748 );
   nand U23535 ( n23732,p1_reg0_reg_18_,n23577 );
   nand U23536 ( p1_u3510,n23749,n23750 );
   nand U23537 ( n23750,n23569,n23512 );
   nand U23538 ( n23512,n23751,n23752,n23753 );
   nor U23539 ( n23753,n23754,n23755,n23756 );
   nor U23540 ( n23756,n23621,n23757 );
   and U23541 ( n23755,n23758,n23575 );
   nor U23542 ( n23754,n23624,n23759 );
   nand U23543 ( n23752,n23626,n23411 );
   nand U23544 ( n23749,p1_reg0_reg_17_,n23577 );
   nand U23545 ( p1_u3507,n23760,n23761 );
   nand U23546 ( n23761,n23569,n23515 );
   nand U23547 ( n23515,n23762,n23763,n23764,n23765 );
   nand U23548 ( n23765,n23766,n23573 );
   nor U23549 ( n23764,n23767,n23768 );
   nor U23550 ( n23768,n23769,n23621 );
   and U23551 ( n23767,n23575,n23770,n23771 );
   nand U23552 ( n23763,n23626,n23414 );
   nand U23553 ( n23760,p1_reg0_reg_16_,n23577 );
   nand U23554 ( p1_u3504,n23772,n23773 );
   nand U23555 ( n23773,n23569,n23518 );
   nand U23556 ( n23518,n23774,n23775,n23776,n23777 );
   nor U23557 ( n23777,n23778,n23779,n23780 );
   nor U23558 ( n23780,n23781,n23608 );
   nor U23559 ( n23779,n23624,n23782 );
   nor U23560 ( n23778,n23783,n23606 );
   nand U23561 ( n23776,n23784,n23655 );
   nand U23562 ( n23774,n23575,n23785 );
   nand U23563 ( n23772,p1_reg0_reg_15_,n23577 );
   nand U23564 ( p1_u3501,n23786,n23787 );
   nand U23565 ( n23787,n23569,n23521 );
   nand U23566 ( n23521,n23788,n23789,n23790,n23791 );
   nor U23567 ( n23791,n23792,n23793,n23794 );
   nor U23568 ( n23794,n23795,n23606 );
   nor U23569 ( n23793,n23796,n23608 );
   or U23570 ( n23790,n23797,n23742 );
   nand U23571 ( n23789,n23798,n23655 );
   nand U23572 ( n23788,n23799,n23573 );
   nand U23573 ( n23786,p1_reg0_reg_14_,n23577 );
   nand U23574 ( p1_u3498,n23800,n23801 );
   nand U23575 ( n23801,n23569,n23524 );
   nand U23576 ( n23524,n23802,n23803,n23804 );
   nor U23577 ( n23804,n23805,n23806,n23807 );
   nor U23578 ( n23807,n23621,n23808 );
   and U23579 ( n23806,n23809,n23575 );
   nor U23580 ( n23805,n23624,n23810 );
   nand U23581 ( n23803,n23626,n23423 );
   nand U23582 ( n23800,p1_reg0_reg_13_,n23577 );
   nand U23583 ( p1_u3495,n23811,n23812 );
   nand U23584 ( n23812,n23569,n23527 );
   nand U23585 ( n23527,n23813,n23814,n23815,n23816 );
   nor U23586 ( n23816,n23817,n23818,n23819 );
   nor U23587 ( n23819,n23820,n23608 );
   nor U23588 ( n23818,n23742,n23821 );
   nor U23589 ( n23817,n23796,n23606 );
   nand U23590 ( n23815,n23822,n23573 );
   nand U23591 ( n23814,n23823,n23655 );
   nand U23592 ( n23813,n23824,n23652 );
   nand U23593 ( n23811,p1_reg0_reg_12_,n23577 );
   nand U23594 ( p1_u3492,n23825,n23826 );
   nand U23595 ( n23826,n23569,n23530 );
   nand U23596 ( n23530,n23827,n23828,n23829 );
   nor U23597 ( n23829,n23830,n23831,n23832 );
   nor U23598 ( n23832,n23621,n23833 );
   and U23599 ( n23831,n23834,n23575 );
   nor U23600 ( n23830,n23624,n23835 );
   nand U23601 ( n23828,n23626,n23429 );
   nand U23602 ( n23825,p1_reg0_reg_11_,n23577 );
   nand U23603 ( p1_u3489,n23836,n23837 );
   nand U23604 ( n23837,n23569,n23533 );
   nand U23605 ( n23533,n23838,n23839,n23840 );
   nor U23606 ( n23840,n23841,n23842,n23843 );
   nor U23607 ( n23843,n23621,n23844 );
   and U23608 ( n23842,n23575,n23845,n23846 );
   nor U23609 ( n23841,n23624,n23847 );
   nand U23610 ( n23839,n23626,n23432 );
   nand U23611 ( n23836,p1_reg0_reg_10_,n23577 );
   nand U23612 ( p1_u3486,n23848,n23849 );
   nand U23613 ( n23849,n23569,n23536 );
   nand U23614 ( n23536,n23850,n23851,n23852,n23853 );
   nor U23615 ( n23853,n23854,n23855,n23856 );
   nor U23616 ( n23856,n23857,n23608 );
   nor U23617 ( n23855,n23624,n23858 );
   nor U23618 ( n23854,n23859,n23606 );
   nand U23619 ( n23852,n23860,n23652 );
   nand U23620 ( n23851,n23575,n23861 );
   nand U23621 ( n23850,n23862,n23655 );
   nand U23622 ( n23848,p1_reg0_reg_9_,n23577 );
   nand U23623 ( p1_u3483,n23863,n23864 );
   nand U23624 ( n23864,n23569,n23539 );
   nand U23625 ( n23539,n23865,n23866,n23867 );
   nor U23626 ( n23867,n23868,n23869,n23870 );
   nor U23627 ( n23870,n23621,n23871 );
   and U23628 ( n23869,n23575,n23872,n23873 );
   nor U23629 ( n23868,n23624,n23874 );
   nand U23630 ( n23866,n23626,n23438 );
   nand U23631 ( n23863,p1_reg0_reg_8_,n23577 );
   nand U23632 ( p1_u3480,n23875,n23876 );
   nand U23633 ( n23876,n23569,n23542 );
   nand U23634 ( n23542,n23877,n23878,n23879 );
   nor U23635 ( n23879,n23880,n23881,n23882 );
   nor U23636 ( n23882,n23621,n23883 );
   and U23637 ( n23881,n23884,n23575 );
   nor U23638 ( n23880,n23624,n23885 );
   nand U23639 ( n23878,n23626,n23441 );
   nand U23640 ( n23875,p1_reg0_reg_7_,n23577 );
   nand U23641 ( p1_u3477,n23886,n23887 );
   nand U23642 ( n23887,n23569,n23545 );
   nand U23643 ( n23545,n23888,n23889,n23890 );
   nor U23644 ( n23890,n23891,n23892,n23893 );
   nor U23645 ( n23893,n23621,n23894 );
   and U23646 ( n23892,n23575,n23895,n23896 );
   nor U23647 ( n23891,n23624,n23897 );
   nand U23648 ( n23889,n23626,n23444 );
   nand U23649 ( n23886,p1_reg0_reg_6_,n23577 );
   nand U23650 ( p1_u3474,n23898,n23899 );
   nand U23651 ( n23899,n23569,n23548 );
   nand U23652 ( n23548,n23900,n23901,n23902 );
   nor U23653 ( n23902,n23903,n23904,n23905 );
   nor U23654 ( n23905,n23906,n23621 );
   and U23655 ( n23904,n23907,n23575 );
   nor U23656 ( n23903,n23624,n23908 );
   nand U23657 ( n23901,n23626,n23447 );
   nand U23658 ( n23898,p1_reg0_reg_5_,n23577 );
   nand U23659 ( p1_u3471,n23909,n23910 );
   nand U23660 ( n23910,n23569,n23551 );
   nand U23661 ( n23551,n23911,n23912,n23913,n23914 );
   nor U23662 ( n23914,n23915,n23916,n23917 );
   nor U23663 ( n23917,n23918,n23608 );
   nor U23664 ( n23916,n23624,n23919 );
   nor U23665 ( n23915,n23920,n23606 );
   or U23666 ( n23913,n23921,n23748 );
   nand U23667 ( n23912,n23922,n23923,n23575 );
   nand U23668 ( n23911,n23924,n23655 );
   nand U23669 ( n23909,p1_reg0_reg_4_,n23577 );
   nand U23670 ( p1_u3468,n23925,n23926 );
   nand U23671 ( n23926,n23569,n23554 );
   nand U23672 ( n23554,n23927,n23928,n23929,n23930 );
   nor U23673 ( n23930,n23931,n23932 );
   nor U23674 ( n23931,n23933,n23606 );
   nand U23675 ( n23929,n23934,n23573 );
   nand U23676 ( n23928,n23575,n23935 );
   nand U23677 ( n23927,n23936,n23655 );
   nand U23678 ( n23925,p1_reg0_reg_3_,n23577 );
   nand U23679 ( p1_u3465,n23937,n23938 );
   nand U23680 ( n23938,n23569,n23557 );
   nand U23681 ( n23557,n23939,n23940,n23941,n23942 );
   nor U23682 ( n23942,n23943,n23944,n23945 );
   nor U23683 ( n23945,n23946,n23608 );
   nor U23684 ( n23944,n23624,n23947 );
   nor U23685 ( n23943,n23918,n23606 );
   nand U23686 ( n23941,n23948,n23655 );
   nand U23687 ( n23939,n23949,n23950,n23575 );
   nand U23688 ( n23937,p1_reg0_reg_2_,n23577 );
   nand U23689 ( p1_u3462,n23951,n23952 );
   nand U23690 ( n23952,n23569,n23560 );
   nand U23691 ( n23560,n23953,n23954,n23955,n23956 );
   nor U23692 ( n23956,n23957,n23958,n23959 );
   nor U23693 ( n23959,n23960,n23608 );
   nor U23694 ( n23958,n23624,n23961 );
   nor U23695 ( n23957,n23962,n23606 );
   nand U23696 ( n23955,n23963,n23652 );
   nand U23697 ( n23954,n23575,n23964 );
   nand U23698 ( n23953,n23965,n23655 );
   or U23699 ( n23655,n23966,n23591 );
   nand U23700 ( n23951,p1_reg0_reg_1_,n23577 );
   nand U23701 ( p1_u3459,n23967,n23968 );
   nand U23702 ( n23968,n23569,n23563 );
   nand U23703 ( n23563,n23969,n23970,n23971,n23972 );
   nand U23704 ( n23972,n23973,n23974 );
   nand U23705 ( n23973,n23624,n23742 );
   nand U23706 ( n23573,n23975,n23976 );
   nand U23707 ( n23971,n23977,n23591 );
   not U23708 ( n23591,n23621 );
   nand U23709 ( n23970,n23626,n23462 );
   nand U23710 ( n23967,p1_reg0_reg_0_,n23577 );
   and U23711 ( n23564,n23981,n23982,n23983 );
   nand U23712 ( n23981,n23984,n23985,n23986 );
   nand U23713 ( n23986,n23987,n23988 );
   nand U23714 ( n23988,n23989,n23990 );
   nand U23715 ( p1_u3446,n23991,n23992 );
   nand U23716 ( n23992,p1_d_reg_1_,n23993 );
   nand U23717 ( n23991,n23994,n23995 );
   nand U23718 ( p1_u3445,n23996,n23997 );
   nand U23719 ( n23997,p1_d_reg_0_,n23993 );
   nand U23720 ( n23996,n23994,n23998 );
   nand U23721 ( p1_u3356,n23999,n24000,n24001,n24002 );
   nor U23722 ( n24002,n24003,n24004,n24005 );
   and U23723 ( n24005,n23592,n24006 );
   and U23724 ( n24004,n24007,n24008 );
   and U23725 ( n24003,n23593,n24009 );
   xor U23726 ( n23593,n23611,n23594 );
   nand U23727 ( n24001,n24010,n23594 );
   nand U23728 ( n24000,p1_reg2_reg_29_,n24011 );
   nand U23729 ( n23999,n24012,n23595 );
   nand U23730 ( n23595,n24013,n24014,n24015,n24016 );
   nand U23731 ( n24016,n23592,n23966 );
   xor U23732 ( n23592,n24017,n24018 );
   nand U23733 ( n24018,n24019,n24020 );
   or U23734 ( n24020,n24021,n24022,n24023 );
   nand U23735 ( n24015,n23652,n24024 );
   nand U23736 ( n24024,n24025,n24026,n24027 );
   nand U23737 ( n24027,n24017,n24028,n24029 );
   nand U23738 ( n24026,n24030,n24031 );
   nand U23739 ( n24031,n24028,n24032 );
   or U23740 ( n24032,n24033,n24029 );
   not U23741 ( n24029,n24034 );
   nand U23742 ( n24028,n24035,n23381 );
   nand U23743 ( n24025,n24033,n24017 );
   nor U23744 ( n24033,n23381,n24035 );
   nand U23745 ( n24014,n24036,n23381 );
   nand U23746 ( n24013,n24037,n23375 );
   nand U23747 ( p1_u3355,n24038,n24039,n24040 );
   nand U23748 ( n24040,n24041,n20618 );
   nand U23749 ( n24039,p1_ir_reg_0_,n24042 );
   or U23750 ( n24042,n24043,n24044 );
   nand U23751 ( n24038,n24045,p2_datao_reg_0_ );
   nand U23752 ( p1_u3354,n24046,n24047,n24048,n24049 );
   nand U23753 ( n24049,n24044,n24050 );
   nand U23754 ( n24048,n24045,p2_datao_reg_1_ );
   nand U23755 ( n24047,n24043,p1_ir_reg_1_ );
   nand U23756 ( n24046,n24041,n20628 );
   nand U23757 ( p1_u3353,n24051,n24052,n24053,n24054 );
   nand U23758 ( n24054,n24055,n24056,n24044 );
   nand U23759 ( n24053,n24045,p2_datao_reg_2_ );
   nand U23760 ( n24052,n24043,p1_ir_reg_2_ );
   nand U23761 ( n24051,n24041,n20635 );
   nand U23762 ( p1_u3352,n24057,n24058,n24059,n24060 );
   nand U23763 ( n24060,n24061,n24044 );
   nand U23764 ( n24059,n24045,p2_datao_reg_3_ );
   nand U23765 ( n24058,n24043,p1_ir_reg_3_ );
   nand U23766 ( n24057,n24041,n20645 );
   nand U23767 ( p1_u3351,n24062,n24063,n24064,n24065 );
   nand U23768 ( n24065,n24066,n24067,n24044 );
   nand U23769 ( n24064,n24045,p2_datao_reg_4_ );
   nand U23770 ( n24063,n24043,p1_ir_reg_4_ );
   nand U23771 ( n24062,n24041,n20652 );
   nand U23772 ( p1_u3350,n24068,n24069,n24070,n24071 );
   nand U23773 ( n24071,p1_ir_reg_5_,n24072 );
   nand U23774 ( n24072,n24073,n24074 );
   nand U23775 ( n24074,n24044,n24075 );
   nand U23776 ( n24070,n24044,n24067,n24076 );
   nand U23777 ( n24069,n24045,p2_datao_reg_5_ );
   nand U23778 ( n24068,n24041,n20661 );
   nand U23779 ( p1_u3349,n24077,n24078,n24079,n24080 );
   nand U23780 ( n24080,n24081,n24082,n24044 );
   nand U23781 ( n24079,n24045,p2_datao_reg_6_ );
   nand U23782 ( n24078,n24043,p1_ir_reg_6_ );
   nand U23783 ( n24077,n24041,n20668 );
   nand U23784 ( p1_u3348,n24083,n24084,n24085,n24086 );
   nand U23785 ( n24086,p1_ir_reg_7_,n24087 );
   nand U23786 ( n24087,n24073,n24088 );
   nand U23787 ( n24088,n24044,n24089 );
   nand U23788 ( n24085,n24044,n24082,n24090 );
   nand U23789 ( n24084,n24045,p2_datao_reg_7_ );
   nand U23790 ( n24083,n24041,n20677 );
   nand U23791 ( p1_u3347,n24091,n24092,n24093,n24094 );
   nand U23792 ( n24094,n24095,n24096,n24044 );
   nand U23793 ( n24093,n24045,p2_datao_reg_8_ );
   nand U23794 ( n24092,n24043,p1_ir_reg_8_ );
   nand U23795 ( n24091,n24041,n20684 );
   nand U23796 ( p1_u3346,n24097,n24098,n24099,n24100 );
   nand U23797 ( n24100,n24101,n24044 );
   nand U23798 ( n24099,n24045,p2_datao_reg_9_ );
   nand U23799 ( n24098,n24043,p1_ir_reg_9_ );
   nand U23800 ( n24097,n24041,n20693 );
   nand U23801 ( p1_u3345,n24102,n24103,n24104,n24105 );
   nand U23802 ( n24105,n24106,n24044 );
   not U23803 ( n24106,n24107 );
   nand U23804 ( n24104,n24045,p2_datao_reg_10_ );
   nand U23805 ( n24103,n24043,p1_ir_reg_10_ );
   nand U23806 ( n24102,n24041,n20700 );
   nand U23807 ( p1_u3344,n24108,n24109,n24110,n24111 );
   nand U23808 ( n24111,n24112,n24044 );
   nand U23809 ( n24110,n24045,p2_datao_reg_11_ );
   nand U23810 ( n24109,n24043,p1_ir_reg_11_ );
   nand U23811 ( n24108,n24041,n20710 );
   nand U23812 ( p1_u3343,n24113,n24114,n24115,n24116 );
   nand U23813 ( n24116,n24117,n24118,n24044 );
   nand U23814 ( n24115,n24045,p2_datao_reg_12_ );
   nand U23815 ( n24114,n24043,p1_ir_reg_12_ );
   nand U23816 ( n24113,n24041,n20717 );
   nand U23817 ( p1_u3342,n24119,n24120,n24121,n24122 );
   nand U23818 ( n24122,p1_ir_reg_13_,n24123 );
   nand U23819 ( n24123,n24073,n24124 );
   nand U23820 ( n24124,n24044,n24125 );
   nand U23821 ( n24121,n24044,n24118,n24126 );
   nand U23822 ( n24120,n24045,p2_datao_reg_13_ );
   nand U23823 ( n24119,n24041,n20727 );
   nand U23824 ( p1_u3341,n24127,n24128,n24129,n24130 );
   nand U23825 ( n24130,n24131,n24044 );
   not U23826 ( n24131,n24132 );
   nand U23827 ( n24129,n24045,p2_datao_reg_14_ );
   nand U23828 ( n24128,n24043,p1_ir_reg_14_ );
   nand U23829 ( n24127,n24041,n20734 );
   nand U23830 ( p1_u3340,n24133,n24134,n24135,n24136 );
   nand U23831 ( n24136,p1_ir_reg_15_,n24137 );
   nand U23832 ( n24137,n24073,n24138 );
   nand U23833 ( n24138,n24044,n24139 );
   nand U23834 ( n24135,n24044,n24140,n24141 );
   nand U23835 ( n24134,n24045,p2_datao_reg_15_ );
   nand U23836 ( n24133,n24041,n20744 );
   nand U23837 ( p1_u3339,n24142,n24143,n24144,n24145 );
   nand U23838 ( n24145,n24146,n24147,n24044 );
   nand U23839 ( n24144,n24045,p2_datao_reg_16_ );
   nand U23840 ( n24143,n24043,p1_ir_reg_16_ );
   nand U23841 ( n24142,n24041,n20751 );
   nand U23842 ( p1_u3338,n24148,n24149,n24150,n24151 );
   nand U23843 ( n24151,p1_ir_reg_17_,n24152 );
   nand U23844 ( n24152,n24073,n24153 );
   nand U23845 ( n24153,n24044,n24154 );
   nand U23846 ( n24150,n24044,n24147,n24155 );
   nand U23847 ( n24149,n24045,p2_datao_reg_17_ );
   nand U23848 ( n24148,n24041,n20761 );
   nand U23849 ( p1_u3337,n24156,n24157,n24158,n24159 );
   nand U23850 ( n24159,p1_ir_reg_18_,n24160 );
   nand U23851 ( n24160,n24073,n24161 );
   nand U23852 ( n24161,n24044,n24162 );
   nand U23853 ( n24158,n24044,n24163,n24164 );
   nand U23854 ( n24157,n24045,p2_datao_reg_18_ );
   nand U23855 ( n24156,n24041,n20768 );
   nand U23856 ( p1_u3336,n24165,n24166,n24167,n24168 );
   nand U23857 ( n24168,n24169,n24170,n24044 );
   nand U23858 ( n24167,n24045,p2_datao_reg_19_ );
   nand U23859 ( n24166,n24043,p1_ir_reg_19_ );
   nand U23860 ( n24165,n24041,n20778 );
   nand U23861 ( p1_u3335,n24171,n24172,n24173,n24174 );
   nand U23862 ( n24174,n24175,n24176,n24044 );
   nand U23863 ( n24173,n24045,p2_datao_reg_20_ );
   nand U23864 ( n24172,n24043,p1_ir_reg_20_ );
   nand U23865 ( n24171,n24041,n20785 );
   nand U23866 ( p1_u3334,n24177,n24178,n24179,n24180 );
   nand U23867 ( n24180,p1_ir_reg_21_,n24181 );
   nand U23868 ( n24181,n24073,n24182 );
   nand U23869 ( n24182,n24044,n24183 );
   nand U23870 ( n24179,n24044,n24176,n24184 );
   nand U23871 ( n24178,n24045,p2_datao_reg_21_ );
   nand U23872 ( n24177,n24041,n20794 );
   nand U23873 ( p1_u3333,n24185,n24186,n24187,n24188 );
   nand U23874 ( n24188,n24189,n24190,n24044 );
   nand U23875 ( n24187,n24045,p2_datao_reg_22_ );
   nand U23876 ( n24186,n24043,p1_ir_reg_22_ );
   nand U23877 ( n24185,n24041,n20804 );
   nand U23878 ( p1_u3332,n24191,n24192,n24193,n24194 );
   nand U23879 ( n24194,p1_ir_reg_23_,n24195 );
   nand U23880 ( n24195,n24073,n24196 );
   nand U23881 ( n24196,n24044,n24197 );
   nand U23882 ( n24193,n24044,n24190,n24198 );
   nand U23883 ( n24192,n24045,p2_datao_reg_23_ );
   nand U23884 ( n24191,n24041,n20811 );
   nand U23885 ( p1_u3331,n24199,n24200,n24201,n24202 );
   nand U23886 ( n24202,n24203,n24204,n24044 );
   nand U23887 ( n24201,n24045,p2_datao_reg_24_ );
   nand U23888 ( n24200,n24043,p1_ir_reg_24_ );
   nand U23889 ( n24199,n24041,n20818 );
   nand U23890 ( p1_u3330,n24205,n24206,n24207,n24208 );
   nand U23891 ( n24208,p1_ir_reg_25_,n24209 );
   nand U23892 ( n24209,n24073,n24210 );
   nand U23893 ( n24210,n24044,n24211 );
   nand U23894 ( n24207,n24044,n24204,n24212 );
   nand U23895 ( n24206,n24045,p2_datao_reg_25_ );
   nand U23896 ( n24205,n24041,n20827 );
   nand U23897 ( p1_u3329,n24213,n24214,n24215,n24216 );
   nand U23898 ( n24216,n24217,n24218,n24044 );
   nand U23899 ( n24215,n24045,p2_datao_reg_26_ );
   nand U23900 ( n24214,n24043,p1_ir_reg_26_ );
   nand U23901 ( n24213,n24041,n20834 );
   nand U23902 ( p1_u3328,n24219,n24220,n24221,n24222 );
   nand U23903 ( n24222,p1_ir_reg_27_,n24223 );
   nand U23904 ( n24223,n24073,n24224 );
   nand U23905 ( n24224,n24044,n24225 );
   nand U23906 ( n24221,n24044,n24218,n24226 );
   nand U23907 ( n24220,n24045,p2_datao_reg_27_ );
   nand U23908 ( n24219,n24041,n20843 );
   nand U23909 ( p1_u3327,n24227,n24228,n24229,n24230 );
   nand U23910 ( n24230,n24231,n24232,n24044 );
   nand U23911 ( n24229,n24045,p2_datao_reg_28_ );
   nand U23912 ( n24228,n24043,p1_ir_reg_28_ );
   nand U23913 ( n24227,n24041,n20853 );
   nand U23914 ( p1_u3326,n24233,n24234,n24235,n24236 );
   nand U23915 ( n24236,p1_ir_reg_29_,n24237 );
   nand U23916 ( n24237,n24073,n24238 );
   nand U23917 ( n24238,n24239,n24044 );
   nand U23918 ( n24235,n24044,n24232,n24240 );
   nand U23919 ( n24234,n24045,p2_datao_reg_29_ );
   nand U23920 ( n24233,n24041,n20860 );
   nand U23921 ( p1_u3325,n24241,n24242,n24243,n24244 );
   nand U23922 ( n24244,p1_ir_reg_30_,n24245 );
   nand U23923 ( n24245,n24073,n24246 );
   nand U23924 ( n24246,n24247,n24044 );
   nand U23925 ( n24243,n24044,n24248,n24249 );
   nand U23926 ( n24242,n24045,p2_datao_reg_30_ );
   nand U23927 ( n24241,n24041,n20869 );
   nand U23928 ( p1_u3324,n24250,n24251,n24252 );
   nand U23929 ( n24252,n24041,n24253 );
   nand U23930 ( n24251,n24044,n24249,n24247 );
   not U23931 ( n24247,n24248 );
   nand U23932 ( n24248,n24239,n24240 );
   nand U23933 ( n24073,p1_state_reg,n24254 );
   nand U23934 ( n24250,n24045,p2_datao_reg_31_ );
   nor U23935 ( p1_u3323,n23994,n24255 );
   and U23936 ( p1_u3322,n23993,p1_d_reg_3_ );
   and U23937 ( p1_u3321,n23993,p1_d_reg_4_ );
   and U23938 ( p1_u3320,n23993,p1_d_reg_5_ );
   nor U23939 ( p1_u3319,n23994,n24256 );
   and U23940 ( p1_u3318,n23993,p1_d_reg_7_ );
   and U23941 ( p1_u3317,n23993,p1_d_reg_8_ );
   and U23942 ( p1_u3316,n23993,p1_d_reg_9_ );
   nor U23943 ( p1_u3315,n23994,n24257 );
   and U23944 ( p1_u3314,n23993,p1_d_reg_11_ );
   and U23945 ( p1_u3313,n23993,p1_d_reg_12_ );
   nor U23946 ( p1_u3312,n23994,n24258 );
   and U23947 ( p1_u3311,n23993,p1_d_reg_14_ );
   and U23948 ( p1_u3310,n23993,p1_d_reg_15_ );
   nor U23949 ( p1_u3309,n23994,n24259 );
   nor U23950 ( p1_u3308,n23994,n24260 );
   nor U23951 ( p1_u3307,n23994,n24261 );
   nor U23952 ( p1_u3306,n23994,n24262 );
   and U23953 ( p1_u3305,n23993,p1_d_reg_20_ );
   and U23954 ( p1_u3304,n23993,p1_d_reg_21_ );
   and U23955 ( p1_u3303,n23993,p1_d_reg_22_ );
   and U23956 ( p1_u3302,n23993,p1_d_reg_23_ );
   and U23957 ( p1_u3301,n23993,p1_d_reg_24_ );
   and U23958 ( p1_u3300,n23993,p1_d_reg_25_ );
   and U23959 ( p1_u3299,n23993,p1_d_reg_26_ );
   nor U23960 ( p1_u3298,n23994,n24263 );
   and U23961 ( p1_u3297,n23993,p1_d_reg_28_ );
   nor U23962 ( p1_u3296,n23994,n24264 );
   and U23963 ( p1_u3295,n23993,p1_d_reg_30_ );
   and U23964 ( p1_u3294,n23993,p1_d_reg_31_ );
   nand U23965 ( p1_u3293,n24266,n24267,n24268,n24269 );
   nor U23966 ( n24269,n24270,n24271,n24272 );
   nor U23967 ( n24272,n23969,n24011 );
   and U23968 ( n23969,n24273,n24274 );
   nand U23969 ( n24274,n24275,n23652 );
   nand U23970 ( n24275,n24276,n24277 );
   nand U23971 ( n24277,n24278,n23465 );
   nand U23972 ( n24273,n23977,n23966 );
   nor U23973 ( n24271,n24012,n24279 );
   and U23974 ( n24270,p1_reg3_reg_0_,n24008 );
   nand U23975 ( n24268,n24006,n23977 );
   nand U23976 ( n24267,n24280,n23974 );
   nand U23977 ( n24280,n24281,n24282 );
   nand U23978 ( n24266,n24283,n23462 );
   nand U23979 ( p1_u3292,n24284,n24285,n24286,n24287 );
   nor U23980 ( n24287,n24288,n24289,n24290,n24291 );
   and U23981 ( n24291,n24292,n23965 );
   xor U23982 ( n23965,n24293,n24294 );
   nor U23983 ( n24290,n23960,n24295 );
   and U23984 ( n24289,n23964,n24009 );
   xor U23985 ( n23964,n23974,n24296 );
   and U23986 ( n24288,n23963,n24297 );
   xor U23987 ( n23963,n24298,n24294 );
   nor U23988 ( n24286,n24299,n24300 );
   nor U23989 ( n24300,n24301,n24302 );
   nor U23990 ( n24299,n23962,n24303 );
   nand U23991 ( n24285,n24010,n24296 );
   nand U23992 ( n24284,p1_reg2_reg_1_,n24011 );
   nand U23993 ( p1_u3291,n24304,n24305,n24306,n24307 );
   nor U23994 ( n24307,n24308,n24309,n24310,n24311 );
   nor U23995 ( n24311,n23918,n24303 );
   and U23996 ( n24310,n24292,n23948 );
   and U23997 ( n23948,n24312,n24313 );
   nand U23998 ( n24313,n24314,n24315 );
   not U23999 ( n24315,n24316 );
   nand U24000 ( n24312,n24317,n24318,n24316 );
   nor U24001 ( n24316,n24319,n24320 );
   nor U24002 ( n24309,n23946,n24295 );
   and U24003 ( n24308,n24009,n23950,n23949 );
   nand U24004 ( n23949,n24321,n24322 );
   nand U24005 ( n24322,n23961,n24278 );
   nor U24006 ( n24306,n24323,n24324 );
   nor U24007 ( n24324,n24011,n23940 );
   nand U24008 ( n23940,n24325,n24326,n24327 );
   nand U24009 ( n24326,n24328,n24317 );
   not U24010 ( n24328,n24329 );
   nand U24011 ( n24325,n24314,n24330 );
   nor U24012 ( n24323,n24012,n24331 );
   nand U24013 ( n24305,n24008,p1_reg3_reg_2_ );
   nand U24014 ( n24304,n24010,n24321 );
   nand U24015 ( p1_u3290,n24332,n24333,n24334,n24335 );
   nor U24016 ( n24335,n24336,n24337,n24338,n24339 );
   nor U24017 ( n24339,n24340,n24281 );
   nor U24018 ( n24338,p1_reg3_reg_3_,n24302 );
   and U24019 ( n24337,n23932,n24012 );
   nand U24020 ( n23932,n24341,n24342,n24343 );
   nand U24021 ( n24343,n24036,n23459 );
   nand U24022 ( n24342,n24344,n24345 );
   nand U24023 ( n24344,n24346,n24347 );
   nand U24024 ( n24341,n24348,n24345 );
   nand U24025 ( n24345,n24349,n24350 );
   nand U24026 ( n24350,n24317,n24329,n24351 );
   nand U24027 ( n24349,n24352,n24353 );
   nor U24028 ( n24336,n24012,n24354 );
   nand U24029 ( n24334,n24283,n23453 );
   nand U24030 ( n24333,n24009,n23935 );
   xor U24031 ( n23935,n24355,n24340 );
   nand U24032 ( n24332,n23936,n24292 );
   xor U24033 ( n23936,n24352,n24356 );
   nand U24034 ( n24356,n24357,n24358 );
   nand U24035 ( n24358,n24319,n24359 );
   nand U24036 ( p1_u3289,n24360,n24361,n24362,n24363 );
   nor U24037 ( n24363,n24364,n24365,n24366,n24367 );
   nor U24038 ( n24367,n23918,n24295 );
   nor U24039 ( n24366,n24368,n24302 );
   nor U24040 ( n24365,n23921,n24369 );
   xor U24041 ( n23921,n24370,n24371 );
   and U24042 ( n24364,n24009,n23923,n23922 );
   nand U24043 ( n23922,n24372,n24373 );
   nand U24044 ( n24373,n24355,n24340 );
   nor U24045 ( n24362,n24374,n24375 );
   nor U24046 ( n24375,n23920,n24303 );
   and U24047 ( n24374,n24292,n23924 );
   xor U24048 ( n23924,n24370,n24376 );
   nand U24049 ( n24361,n24010,n24372 );
   nand U24050 ( n24360,p1_reg2_reg_4_,n24011 );
   nand U24051 ( p1_u3288,n24377,n24378,n24379,n24380 );
   nor U24052 ( n24380,n24381,n24382,n24383,n24384 );
   nor U24053 ( n24384,n23908,n24281 );
   and U24054 ( n24383,n24385,n24008 );
   nor U24055 ( n24382,n23900,n24011 );
   and U24056 ( n23900,n24386,n24387,n24388,n24389 );
   nor U24057 ( n24389,n24390,n24391,n24392,n24393 );
   nor U24058 ( n24393,n23906,n24394 );
   nor U24059 ( n24392,n23906,n24395 );
   nor U24060 ( n24391,n24347,n24396 );
   nor U24061 ( n24390,n24397,n24396 );
   nor U24062 ( n24388,n24398,n24399 );
   nor U24063 ( n24399,n24400,n24396 );
   nor U24064 ( n24398,n23906,n24401 );
   not U24065 ( n23906,n24402 );
   or U24066 ( n24387,n24396,n24403 );
   nand U24067 ( n24396,n24404,n24405 );
   nand U24068 ( n24405,n24406,n24407,n24408 );
   nand U24069 ( n24404,n24409,n24410 );
   nand U24070 ( n24386,n24036,n23453 );
   nor U24071 ( n24381,n24012,n24411 );
   nand U24072 ( n24379,n24283,n23447 );
   nand U24073 ( n24378,n24009,n23907 );
   xor U24074 ( n23907,n24412,n23923 );
   nand U24075 ( n24377,n24006,n24402 );
   xor U24076 ( n24402,n24413,n24409 );
   nor U24077 ( n24413,n24414,n24415 );
   nor U24078 ( n24414,n24416,n24376 );
   nand U24079 ( p1_u3287,n24417,n24418,n24419,n24420 );
   nor U24080 ( n24420,n24421,n24422,n24423,n24424 );
   nor U24081 ( n24424,n23897,n24281 );
   nor U24082 ( n24423,n24425,n24302 );
   nor U24083 ( n24422,n23888,n24011 );
   and U24084 ( n23888,n24426,n24427 );
   nor U24085 ( n24427,n24428,n24429,n24430,n24431 );
   nor U24086 ( n24431,n24432,n24400 );
   nor U24087 ( n24430,n24401,n23894 );
   nor U24088 ( n24429,n24432,n24403 );
   nor U24089 ( n24428,n24432,n24347 );
   nor U24090 ( n24426,n24433,n24434,n24435,n24436 );
   nor U24091 ( n24436,n23920,n23608 );
   nor U24092 ( n24435,n24394,n23894 );
   nor U24093 ( n24434,n24432,n24397 );
   nor U24094 ( n24432,n24437,n24438 );
   nor U24095 ( n24438,n24439,n24440 );
   nand U24096 ( n24440,n24441,n24442 );
   nand U24097 ( n24442,n24410,n24407 );
   not U24098 ( n24410,n24408 );
   not U24099 ( n24439,n24406 );
   nor U24100 ( n24437,n24443,n24444 );
   nor U24101 ( n24433,n24395,n23894 );
   nor U24102 ( n24421,n24012,n24445 );
   nand U24103 ( n24419,n24283,n23444 );
   nand U24104 ( n24418,n23896,n23895,n24009 );
   nand U24105 ( n23896,n24446,n24447 );
   nand U24106 ( n24447,n24448,n23908 );
   or U24107 ( n24417,n24449,n23894 );
   xor U24108 ( n23894,n24441,n24450 );
   nand U24109 ( p1_u3286,n24451,n24452,n24453,n24454 );
   nor U24110 ( n24454,n24455,n24456,n24457,n24458 );
   nor U24111 ( n24458,n23885,n24281 );
   and U24112 ( n24457,n24459,n24008 );
   nor U24113 ( n24456,n23877,n24011 );
   and U24114 ( n23877,n24460,n24461,n24462,n24463 );
   nor U24115 ( n24463,n24464,n24465,n24466,n24467 );
   nor U24116 ( n24467,n24394,n23883 );
   nor U24117 ( n24466,n24401,n23883 );
   nor U24118 ( n24465,n24395,n23883 );
   nor U24119 ( n24464,n24400,n24468 );
   nor U24120 ( n24462,n24469,n24470 );
   nor U24121 ( n24470,n24471,n23608 );
   nor U24122 ( n24469,n24397,n24468 );
   nand U24123 ( n24461,n24472,n24473 );
   nand U24124 ( n24460,n24472,n24474 );
   not U24125 ( n24472,n24468 );
   nand U24126 ( n24468,n24475,n24476 );
   nand U24127 ( n24476,n24477,n24478 );
   nand U24128 ( n24475,n24479,n24480 );
   nor U24129 ( n24455,n24012,n24481 );
   nand U24130 ( n24453,n24283,n23441 );
   nand U24131 ( n24452,n24009,n23884 );
   xor U24132 ( n23884,n23895,n24482 );
   or U24133 ( n24451,n24449,n23883 );
   nand U24134 ( n23883,n24483,n24484 );
   nand U24135 ( n24484,n24485,n24486,n24487 );
   nand U24136 ( n24483,n24488,n24489,n24479 );
   nand U24137 ( n24488,n24450,n24486 );
   not U24138 ( n24450,n24490 );
   nand U24139 ( p1_u3285,n24491,n24492,n24493,n24494 );
   nor U24140 ( n24494,n24495,n24496,n24497,n24498 );
   nor U24141 ( n24498,n23874,n24281 );
   nor U24142 ( n24497,n24499,n24302 );
   nor U24143 ( n24496,n23865,n24011 );
   and U24144 ( n23865,n24500,n24501,n24502,n24503 );
   nor U24145 ( n24503,n24504,n24505,n24506,n24507 );
   nor U24146 ( n24507,n24508,n24403 );
   xor U24147 ( n24508,n24509,n24510 );
   nor U24148 ( n24506,n24511,n24400 );
   nor U24149 ( n24511,n24512,n24513 );
   not U24150 ( n24513,n24514 );
   nor U24151 ( n24512,n24509,n24510 );
   nor U24152 ( n24505,n24395,n23871 );
   not U24153 ( n23871,n24515 );
   nor U24154 ( n24504,n24516,n23608 );
   nand U24155 ( n24502,n24515,n24517 );
   nand U24156 ( n24501,n24518,n24519 );
   nand U24157 ( n24519,n24520,n24514 );
   nand U24158 ( n24514,n24509,n24510 );
   nand U24159 ( n24520,n24521,n24522 );
   nand U24160 ( n24518,n24347,n24397 );
   nand U24161 ( n24500,n24515,n24523 );
   nor U24162 ( n24495,n24012,n24524 );
   nand U24163 ( n24493,n24283,n23438 );
   nand U24164 ( n24492,n23873,n23872,n24009 );
   nand U24165 ( n23873,n24525,n24526 );
   nand U24166 ( n24526,n24527,n23885 );
   nand U24167 ( n24491,n24006,n24515 );
   xor U24168 ( n24515,n24521,n24528 );
   nand U24169 ( p1_u3284,n24529,n24530,n24531,n24532 );
   nor U24170 ( n24532,n24533,n24534,n24535,n24536 );
   and U24171 ( n24536,n24011,p1_reg2_reg_9_ );
   nor U24172 ( n24535,n23858,n24281 );
   and U24173 ( n24534,n24537,n24008 );
   nor U24174 ( n24533,n23859,n24303 );
   nor U24175 ( n24531,n24538,n24539 );
   and U24176 ( n24539,n24292,n23862 );
   xor U24177 ( n23862,n24540,n24541 );
   nor U24178 ( n24538,n23857,n24295 );
   nand U24179 ( n24530,n24297,n23860 );
   nand U24180 ( n23860,n24542,n24543 );
   nand U24181 ( n24543,n24544,n24540 );
   not U24182 ( n24544,n24545 );
   nand U24183 ( n24542,n24546,n24545 );
   nand U24184 ( n24546,n24547,n24548 );
   nand U24185 ( n24529,n24009,n23861 );
   xor U24186 ( n23861,n23858,n24549 );
   nand U24187 ( p1_u3283,n24550,n24551,n24552,n24553 );
   nor U24188 ( n24553,n24554,n24555,n24556,n24557 );
   nor U24189 ( n24557,n23847,n24281 );
   nor U24190 ( n24556,n24558,n24302 );
   nor U24191 ( n24555,n23838,n24011 );
   and U24192 ( n23838,n24559,n24560,n24561,n24562 );
   nor U24193 ( n24562,n24563,n24564,n24565,n24566 );
   nor U24194 ( n24566,n24397,n24567 );
   nor U24195 ( n24565,n24394,n23844 );
   nor U24196 ( n24564,n24401,n23844 );
   nor U24197 ( n24563,n24395,n23844 );
   nand U24198 ( n24561,n24568,n24473 );
   nand U24199 ( n24560,n24568,n24569 );
   nand U24200 ( n24569,n24403,n24400 );
   not U24201 ( n24568,n24567 );
   nand U24202 ( n24567,n24570,n24571 );
   nand U24203 ( n24571,n24572,n24573,n24574 );
   nand U24204 ( n24570,n24575,n24576 );
   nand U24205 ( n24559,n24036,n23438 );
   nor U24206 ( n24554,n24012,n24577 );
   nand U24207 ( n24552,n24283,n23432 );
   nand U24208 ( n24551,n23846,n23845,n24009 );
   nand U24209 ( n23846,n24578,n24579 );
   nand U24210 ( n24579,n24549,n23858 );
   or U24211 ( n24550,n24449,n23844 );
   nand U24212 ( n23844,n24580,n24581 );
   nand U24213 ( n24581,n24582,n24583,n24584 );
   nand U24214 ( n24580,n24585,n24586,n24575 );
   nand U24215 ( n24585,n24541,n24583 );
   not U24216 ( n24541,n24587 );
   nand U24217 ( p1_u3282,n24588,n24589,n24590,n24591 );
   nor U24218 ( n24591,n24592,n24593,n24594,n24595 );
   nor U24219 ( n24595,n23835,n24281 );
   nor U24220 ( n24594,n24596,n24302 );
   nor U24221 ( n24593,n23827,n24011 );
   and U24222 ( n23827,n24597,n24598 );
   nor U24223 ( n24598,n24599,n24600,n24601,n24602 );
   nor U24224 ( n24602,n24603,n24400 );
   nor U24225 ( n24601,n24395,n23833 );
   nor U24226 ( n24600,n23859,n23608 );
   nor U24227 ( n24599,n24603,n24347 );
   nor U24228 ( n24597,n24604,n24605,n24606,n24607 );
   nor U24229 ( n24607,n24603,n24397 );
   and U24230 ( n24603,n24608,n24609,n24610 );
   not U24231 ( n24610,n24611 );
   nand U24232 ( n24609,n24612,n24574 );
   nand U24233 ( n24608,n24576,n24613 );
   nor U24234 ( n24606,n24394,n23833 );
   nor U24235 ( n24605,n24401,n23833 );
   nor U24236 ( n24604,n24614,n24403 );
   nor U24237 ( n24614,n24611,n24615,n24616 );
   nor U24238 ( n24616,n24617,n24574 );
   and U24239 ( n24615,n24574,n24612 );
   not U24240 ( n24574,n24576 );
   nor U24241 ( n24576,n24618,n24619 );
   nand U24242 ( n24611,n24620,n24621 );
   nand U24243 ( n24621,n24622,n24612 );
   nor U24244 ( n24612,n24623,n24624 );
   not U24245 ( n24622,n24572 );
   nand U24246 ( n24620,n24624,n24613 );
   not U24247 ( n24613,n24617 );
   nand U24248 ( n24617,n24625,n24626 );
   not U24249 ( n24624,n24573 );
   nor U24250 ( n24592,n24012,n24627 );
   nand U24251 ( n24590,n24283,n23429 );
   nand U24252 ( n24589,n24009,n23834 );
   xor U24253 ( n23834,n23845,n24628 );
   or U24254 ( n24588,n24449,n23833 );
   xor U24255 ( n23833,n24623,n24629 );
   nand U24256 ( p1_u3281,n24630,n24631,n24632,n24633 );
   nor U24257 ( n24633,n24634,n24635,n24636,n24637 );
   nor U24258 ( n24637,n24012,n24638 );
   nor U24259 ( n24636,n24639,n24281 );
   nor U24260 ( n24635,n24640,n24302 );
   nor U24261 ( n24634,n23796,n24303 );
   nor U24262 ( n24632,n24641,n24642 );
   nor U24263 ( n24642,n23821,n24282 );
   nand U24264 ( n23821,n24643,n24644 );
   nand U24265 ( n24644,n24645,n23822 );
   nand U24266 ( n24645,n24646,n23835 );
   and U24267 ( n24641,n24292,n23823 );
   xor U24268 ( n23823,n24647,n24648 );
   nand U24269 ( n24631,n24297,n23824 );
   xor U24270 ( n23824,n24649,n24647 );
   or U24271 ( n24630,n24295,n23820 );
   nand U24272 ( p1_u3280,n24650,n24651,n24652,n24653 );
   nor U24273 ( n24653,n24654,n24655,n24656,n24657 );
   nor U24274 ( n24657,n23810,n24281 );
   nor U24275 ( n24656,n24658,n24302 );
   nor U24276 ( n24655,n23802,n24011 );
   and U24277 ( n23802,n24659,n24660,n24661,n24662 );
   nor U24278 ( n24662,n24663,n24664,n24665,n24666 );
   nor U24279 ( n24666,n24394,n23808 );
   nor U24280 ( n24665,n24401,n23808 );
   nor U24281 ( n24664,n24395,n23808 );
   nor U24282 ( n24663,n24347,n24667 );
   nor U24283 ( n24661,n24668,n24669 );
   nor U24284 ( n24669,n24670,n23608 );
   nor U24285 ( n24668,n24403,n24667 );
   not U24286 ( n24667,n24671 );
   nand U24287 ( n24660,n24671,n24348 );
   nand U24288 ( n24659,n24671,n24672 );
   xor U24289 ( n24671,n24673,n24674 );
   nor U24290 ( n24654,n24012,n24675 );
   nand U24291 ( n24652,n24283,n23423 );
   nand U24292 ( n24651,n24009,n23809 );
   xor U24293 ( n23809,n24676,n24643 );
   or U24294 ( n24650,n24449,n23808 );
   nand U24295 ( n23808,n24677,n24678 );
   nand U24296 ( n24678,n24679,n24680,n24674 );
   nand U24297 ( n24679,n24681,n24682 );
   not U24298 ( n24682,n24648 );
   nand U24299 ( n24677,n24683,n24681,n24684 );
   not U24300 ( n24684,n24674 );
   nand U24301 ( n24683,n24648,n24680 );
   nor U24302 ( n24648,n24685,n24686 );
   nand U24303 ( p1_u3279,n24687,n24688,n24689,n24690 );
   nor U24304 ( n24690,n24691,n24692,n24693,n24694 );
   nor U24305 ( n24694,n23795,n24303 );
   nor U24306 ( n24693,n23797,n24282 );
   nand U24307 ( n23797,n24695,n24696 );
   nand U24308 ( n24696,n24697,n23799 );
   nand U24309 ( n24697,n24698,n23810 );
   and U24310 ( n24692,n24292,n23798 );
   xor U24311 ( n23798,n24699,n24700 );
   nor U24312 ( n24691,n23796,n24295 );
   nor U24313 ( n24689,n24701,n24702 );
   nor U24314 ( n24702,n24703,n24281 );
   nor U24315 ( n24701,n24704,n24302 );
   nand U24316 ( n24688,p1_reg2_reg_14_,n24011 );
   nand U24317 ( n24687,n24012,n23792 );
   nand U24318 ( n23792,n24705,n24706 );
   nand U24319 ( n24706,n24707,n24708,n24473 );
   nand U24320 ( n24707,n24709,n24710 );
   nand U24321 ( n24705,n24711,n24708,n24712 );
   nand U24322 ( n24708,n24700,n24713 );
   nand U24323 ( n24711,n24714,n24710,n24715 );
   nand U24324 ( p1_u3278,n24716,n24717,n24718,n24719 );
   nor U24325 ( n24719,n24720,n24721,n24722,n24723 );
   nor U24326 ( n24723,n23783,n24303 );
   and U24327 ( n24722,n24292,n23784 );
   xor U24328 ( n23784,n24724,n24725 );
   nor U24329 ( n24721,n23781,n24295 );
   and U24330 ( n24720,n23785,n24009 );
   xor U24331 ( n23785,n24695,n24726 );
   nor U24332 ( n24718,n24727,n24728 );
   nor U24333 ( n24728,n24011,n23775 );
   nand U24334 ( n23775,n24729,n24730,n23652 );
   nand U24335 ( n24730,n24731,n24732,n24733 );
   nand U24336 ( n24729,n24725,n24734 );
   nor U24337 ( n24727,n24012,n24735 );
   nand U24338 ( n24717,n24008,n24736 );
   nand U24339 ( n24716,n24010,n24726 );
   nand U24340 ( p1_u3277,n24737,n24738,n24739,n24740 );
   nor U24341 ( n24740,n24741,n24742,n24743,n24744 );
   nor U24342 ( n24744,n24745,n24281 );
   nor U24343 ( n24743,n24746,n24302 );
   nor U24344 ( n24742,n23762,n24011 );
   and U24345 ( n23762,n24747,n24748 );
   nor U24346 ( n24748,n24749,n24750,n24751,n24752 );
   nor U24347 ( n24752,n24753,n24400 );
   nor U24348 ( n24751,n23769,n24395 );
   nor U24349 ( n24750,n23795,n23608 );
   nor U24350 ( n24749,n24753,n24347 );
   nor U24351 ( n24747,n24754,n24755,n24756,n24757 );
   nor U24352 ( n24757,n24753,n24397 );
   and U24353 ( n24753,n24758,n24759,n24760 );
   not U24354 ( n24760,n24761 );
   nand U24355 ( n24759,n24762,n24733 );
   nand U24356 ( n24758,n24734,n24763 );
   nor U24357 ( n24756,n23769,n24394 );
   nor U24358 ( n24755,n23769,n24401 );
   nor U24359 ( n24754,n24764,n24403 );
   nor U24360 ( n24764,n24761,n24765,n24766 );
   nor U24361 ( n24766,n24767,n24733 );
   and U24362 ( n24765,n24733,n24762 );
   not U24363 ( n24733,n24734 );
   nor U24364 ( n24734,n24709,n24768 );
   nand U24365 ( n24761,n24769,n24770 );
   nand U24366 ( n24770,n24771,n24762 );
   nor U24367 ( n24762,n24772,n24773 );
   not U24368 ( n24771,n24731 );
   nand U24369 ( n24769,n24773,n24763 );
   not U24370 ( n24763,n24767 );
   nand U24371 ( n24767,n24774,n24775 );
   not U24372 ( n24773,n24732 );
   nor U24373 ( n24741,n24012,n24776 );
   nand U24374 ( n24739,n24283,n23414 );
   nand U24375 ( n24738,n23771,n23770,n24009 );
   nand U24376 ( n23771,n23766,n24777 );
   nand U24377 ( n24777,n24778,n23782 );
   or U24378 ( n24737,n24449,n23769 );
   xor U24379 ( n23769,n24772,n24779 );
   nand U24380 ( p1_u3276,n24780,n24781,n24782,n24783 );
   nor U24381 ( n24783,n24784,n24785,n24786,n24787 );
   nor U24382 ( n24787,n23759,n24281 );
   nor U24383 ( n24786,n24788,n24302 );
   nor U24384 ( n24785,n23751,n24011 );
   and U24385 ( n23751,n24789,n24790,n24791,n24792 );
   nor U24386 ( n24792,n24793,n24794,n24795,n24796 );
   nor U24387 ( n24796,n24797,n24397 );
   nor U24388 ( n24795,n24797,n24400 );
   nor U24389 ( n24794,n23783,n23608 );
   nor U24390 ( n24793,n24797,n24403 );
   nor U24391 ( n24791,n24798,n24799 );
   nor U24392 ( n24799,n24395,n23757 );
   nor U24393 ( n24798,n24797,n24347 );
   xor U24394 ( n24797,n24800,n24801 );
   nand U24395 ( n24790,n24802,n24523 );
   nand U24396 ( n24789,n24802,n24517 );
   nor U24397 ( n24784,n24012,n24803 );
   nand U24398 ( n24782,n24283,n23411 );
   nand U24399 ( n24781,n24009,n23758 );
   xor U24400 ( n23758,n24804,n23770 );
   nand U24401 ( n24780,n24006,n24802 );
   not U24402 ( n24802,n23757 );
   nand U24403 ( n23757,n24805,n24806 );
   nand U24404 ( n24806,n24807,n24808,n24809 );
   nand U24405 ( n24805,n24810,n24811,n24800 );
   not U24406 ( n24800,n24809 );
   nand U24407 ( n24810,n24808,n24812 );
   nand U24408 ( p1_u3275,n24813,n24814,n24815,n24816 );
   nor U24409 ( n24816,n24817,n24818,n24819,n24820 );
   nor U24410 ( n24820,n24012,n24821 );
   nor U24411 ( n24819,n24822,n24281 );
   nor U24412 ( n24818,n24823,n24302 );
   nor U24413 ( n24817,n23744,n24303 );
   nor U24414 ( n24815,n24824,n24825 );
   nor U24415 ( n24825,n23741,n24295 );
   nor U24416 ( n24824,n23747,n24369 );
   xor U24417 ( n23747,n24826,n24827 );
   nand U24418 ( n24814,n23746,n24292 );
   xor U24419 ( n23746,n24828,n24829 );
   or U24420 ( n24813,n24282,n23743 );
   nand U24421 ( n23743,n24830,n24831 );
   nand U24422 ( n24831,n24832,n23745 );
   nand U24423 ( n24832,n24833,n23759 );
   nand U24424 ( p1_u3274,n24834,n24835,n24836,n24837 );
   nor U24425 ( n24837,n24838,n24839,n24840,n24841 );
   nor U24426 ( n24841,n24842,n24281 );
   nor U24427 ( n24840,n24843,n24302 );
   and U24428 ( n24839,n23727,n24012 );
   nand U24429 ( n23727,n24844,n24845,n24846 );
   nand U24430 ( n24846,n24036,n23411 );
   or U24431 ( n24845,n24847,n23748 );
   xor U24432 ( n24847,n24848,n24849 );
   nand U24433 ( n24844,n23731,n23966 );
   nor U24434 ( n24838,n24012,n24850 );
   nand U24435 ( n24836,n24283,n23405 );
   nand U24436 ( n24835,n24009,n23730 );
   xor U24437 ( n23730,n24851,n24842 );
   nand U24438 ( n24834,n24006,n23731 );
   xor U24439 ( n23731,n24848,n24852 );
   nand U24440 ( p1_u3273,n24853,n24854,n24855,n24856 );
   nor U24441 ( n24856,n24857,n24858,n24859,n24860 );
   nor U24442 ( n24860,n23719,n24281 );
   nor U24443 ( n24859,n24861,n24302 );
   nor U24444 ( n24858,n23710,n24011 );
   and U24445 ( n23710,n24862,n24863,n24864,n24865 );
   nor U24446 ( n24865,n24866,n24867,n24868,n24869 );
   nor U24447 ( n24869,n24394,n23716 );
   nor U24448 ( n24868,n24401,n23716 );
   nor U24449 ( n24867,n24395,n23716 );
   nor U24450 ( n24866,n24400,n24870 );
   nor U24451 ( n24864,n24871,n24872 );
   nor U24452 ( n24872,n23744,n23608 );
   nor U24453 ( n24871,n24397,n24870 );
   nand U24454 ( n24863,n24873,n24473 );
   not U24455 ( n24473,n24347 );
   nand U24456 ( n24862,n24873,n24474 );
   not U24457 ( n24873,n24870 );
   xor U24458 ( n24870,n24874,n24875 );
   and U24459 ( n24857,n24011,p1_reg2_reg_20_ );
   nand U24460 ( n24855,n24283,n23402 );
   nand U24461 ( n24854,n23718,n23717,n24009 );
   nand U24462 ( n23718,n24876,n24877 );
   nand U24463 ( n24877,n24851,n24842 );
   or U24464 ( n24853,n24449,n23716 );
   nand U24465 ( n23716,n24878,n24879 );
   nand U24466 ( n24879,n24880,n24881,n24882 );
   nand U24467 ( n24880,n24852,n24883 );
   nand U24468 ( n24878,n24874,n24883,n24884 );
   nand U24469 ( n24884,n24885,n24886 );
   nand U24470 ( p1_u3272,n24887,n24888,n24889,n24890 );
   nor U24471 ( n24890,n24891,n24892,n24893,n24894 );
   nor U24472 ( n24894,n23707,n24281 );
   nor U24473 ( n24893,n24895,n24302 );
   nor U24474 ( n24892,n23699,n24011 );
   and U24475 ( n23699,n24896,n24897,n24898,n24899 );
   nor U24476 ( n24899,n24900,n24901 );
   nor U24477 ( n24901,n23728,n23608 );
   nor U24478 ( n24900,n24346,n24902,n24903 );
   nor U24479 ( n24903,n24904,n24905,n24906 );
   and U24480 ( n24902,n24904,n24907 );
   or U24481 ( n24898,n23705,n24908 );
   nand U24482 ( n24897,n24517,n24909,n24910,n24911 );
   nand U24483 ( n24896,n24912,n24913,n24914 );
   nand U24484 ( n24914,n24400,n24347 );
   nand U24485 ( n24913,n24915,n24916 );
   nand U24486 ( n24912,n24907,n24904 );
   and U24487 ( n24891,n24011,p1_reg2_reg_21_ );
   nand U24488 ( n24889,n24283,n23399 );
   nand U24489 ( n24888,n24009,n23706 );
   xor U24490 ( n23706,n24917,n23717 );
   or U24491 ( n24887,n24449,n23705 );
   nand U24492 ( n23705,n24910,n24911,n24909 );
   nand U24493 ( n24909,n24882,n24885,n24907 );
   nand U24494 ( n24911,n24907,n24918 );
   not U24495 ( n24907,n24919 );
   nand U24496 ( n24910,n24920,n24919,n24921 );
   nand U24497 ( n24920,n24882,n24885 );
   not U24498 ( n24885,n24852 );
   nor U24499 ( n24852,n24922,n24923 );
   nand U24500 ( p1_u3271,n24924,n24925,n24926,n24927 );
   nor U24501 ( n24927,n24928,n24929,n24930,n24931 );
   nor U24502 ( n24931,n23665,n24303 );
   and U24503 ( n24930,n24292,n23694 );
   xor U24504 ( n23694,n24932,n24933 );
   nor U24505 ( n24929,n23692,n24295 );
   and U24506 ( n24928,n24009,n23696,n23695 );
   nand U24507 ( n23695,n24934,n24935 );
   nand U24508 ( n24935,n24936,n23707 );
   nor U24509 ( n24926,n24937,n24938 );
   nor U24510 ( n24938,n24011,n23686 );
   nand U24511 ( n23686,n24939,n24940,n23652 );
   nand U24512 ( n24940,n24941,n24942,n24943 );
   nand U24513 ( n24939,n24932,n24944 );
   and U24514 ( n24937,n24011,p1_reg2_reg_22_ );
   nand U24515 ( n24925,n24008,n24945 );
   not U24516 ( n24008,n24302 );
   nand U24517 ( n24924,n24010,n24934 );
   nand U24518 ( p1_u3270,n24946,n24947,n24948,n24949 );
   nor U24519 ( n24949,n24950,n24951,n24952,n24953 );
   nor U24520 ( n24953,n23682,n24281 );
   nor U24521 ( n24952,n24954,n24302 );
   nor U24522 ( n24951,n23674,n24011 );
   and U24523 ( n23674,n24955,n24956,n24957,n24958 );
   nor U24524 ( n24958,n24959,n24960,n24961,n24962 );
   nor U24525 ( n24962,n23680,n24395 );
   nor U24526 ( n24961,n23680,n24394 );
   nor U24527 ( n24960,n24963,n23608 );
   nor U24528 ( n24959,n24964,n24347 );
   nor U24529 ( n24957,n24965,n24966 );
   nor U24530 ( n24966,n24964,n24403 );
   nor U24531 ( n24965,n24964,n24397 );
   and U24532 ( n24964,n24967,n24968 );
   nand U24533 ( n24967,n24969,n24970 );
   nand U24534 ( n24970,n24942,n24943 );
   not U24535 ( n24969,n24971 );
   nand U24536 ( n24956,n24523,n24972 );
   nand U24537 ( n24955,n24973,n24974,n24348 );
   nand U24538 ( n24974,n24943,n24942,n24975 );
   not U24539 ( n24943,n24944 );
   nand U24540 ( n24973,n24968,n24971 );
   nand U24541 ( n24971,n24975,n24941 );
   nand U24542 ( n24968,n24976,n24977 );
   nand U24543 ( n24977,n24944,n24941 );
   nor U24544 ( n24944,n24915,n24905 );
   and U24545 ( n24976,n24978,n24942 );
   and U24546 ( n24950,n24011,p1_reg2_reg_23_ );
   nand U24547 ( n24948,n24283,n23393 );
   nand U24548 ( n24947,n24009,n23681 );
   xor U24549 ( n23681,n23696,n24979 );
   nand U24550 ( n24946,n24006,n24972 );
   not U24551 ( n24972,n23680 );
   xor U24552 ( n23680,n24978,n24980 );
   nand U24553 ( p1_u3269,n24981,n24982,n24983,n24984 );
   nor U24554 ( n24984,n24985,n24986,n24987,n24988 );
   and U24555 ( n24988,n24011,p1_reg2_reg_24_ );
   nor U24556 ( n24987,n23666,n24281 );
   nor U24557 ( n24986,n24989,n24302 );
   nor U24558 ( n24985,n23667,n24303 );
   nor U24559 ( n24983,n24990,n24991 );
   and U24560 ( n24991,n24292,n23671 );
   xor U24561 ( n23671,n24992,n24993 );
   nor U24562 ( n24990,n23665,n24295 );
   nand U24563 ( n24982,n23669,n23670,n24009 );
   nand U24564 ( n23669,n24994,n24995 );
   nand U24565 ( n24995,n24996,n23682 );
   nand U24566 ( n24981,n24297,n23668 );
   xor U24567 ( n23668,n24993,n24997 );
   nand U24568 ( p1_u3268,n24998,n24999,n25000,n25001 );
   nor U24569 ( n25001,n25002,n25003,n25004,n25005 );
   and U24570 ( n25005,n24011,p1_reg2_reg_25_ );
   nor U24571 ( n25004,n23649,n24281 );
   nor U24572 ( n25003,n25006,n24302 );
   nor U24573 ( n25002,n23650,n24303 );
   nor U24574 ( n25000,n25007,n25008 );
   and U24575 ( n25008,n24292,n23654 );
   xor U24576 ( n23654,n25009,n25010 );
   nand U24577 ( n24292,n24449,n25011 );
   nand U24578 ( n25011,n24012,n23966 );
   nand U24579 ( n23966,n24908,n24394 );
   nor U24580 ( n24908,n25012,n24523 );
   nor U24581 ( n25007,n23648,n24295 );
   nand U24582 ( n24999,n24297,n23651 );
   xor U24583 ( n23651,n25013,n25014 );
   not U24584 ( n25013,n25010 );
   not U24585 ( n24297,n24369 );
   nand U24586 ( n24369,n24012,n23652 );
   nand U24587 ( n24998,n24009,n23653 );
   xor U24588 ( n23653,n25015,n23649 );
   nand U24589 ( p1_u3267,n25016,n25017,n25018,n25019 );
   nor U24590 ( n25019,n25020,n25021,n25022,n25023 );
   nor U24591 ( n25023,n23638,n24281 );
   nor U24592 ( n25022,n25024,n24302 );
   nor U24593 ( n25021,n23629,n24011 );
   and U24594 ( n23629,n25025,n25026,n25027,n25028 );
   nor U24595 ( n25028,n25029,n25030,n25031,n25032 );
   nor U24596 ( n25032,n24394,n23635 );
   nor U24597 ( n25031,n24401,n23635 );
   nor U24598 ( n25030,n24395,n23635 );
   nor U24599 ( n25029,n24400,n25033,n25034 );
   nor U24600 ( n25027,n25035,n25036 );
   nor U24601 ( n25036,n24347,n25033,n25034 );
   nor U24602 ( n25035,n24397,n25033,n25034 );
   nor U24603 ( n25034,n25037,n25038 );
   not U24604 ( n25037,n25039 );
   nor U24605 ( n25033,n25040,n25041 );
   nand U24606 ( n25026,n24036,n23390 );
   nand U24607 ( n25025,n25042,n25043,n24474 );
   nand U24608 ( n25043,n25044,n25045 );
   or U24609 ( n25042,n25046,n25038,n25045 );
   and U24610 ( n25020,n24011,p1_reg2_reg_26_ );
   nand U24611 ( n25018,n24283,n23384 );
   nand U24612 ( n25017,n23637,n23636,n24009 );
   nand U24613 ( n23637,n25047,n25048 );
   nand U24614 ( n25048,n25015,n23649 );
   or U24615 ( n25016,n24449,n23635 );
   nand U24616 ( n23635,n25049,n25050 );
   nand U24617 ( n25050,n25051,n25052,n25040 );
   nand U24618 ( n25051,n25053,n25054 );
   not U24619 ( n25053,n25009 );
   nand U24620 ( n25049,n25055,n25054,n25044 );
   not U24621 ( n25044,n25040 );
   nand U24622 ( n25055,n25052,n25009 );
   nand U24623 ( n25009,n25056,n25057 );
   nand U24624 ( n25057,n25058,n24992 );
   nand U24625 ( p1_u3266,n25059,n25060,n25061,n25062 );
   nor U24626 ( n25062,n25063,n25064,n25065,n25066 );
   nor U24627 ( n25066,n23625,n24281 );
   nor U24628 ( n25065,n25067,n24302 );
   nor U24629 ( n25064,n23615,n24011 );
   and U24630 ( n23615,n25068,n25069,n25070,n25071 );
   nor U24631 ( n25071,n25072,n25073,n25074,n25075 );
   nor U24632 ( n25075,n25076,n24400 );
   nor U24633 ( n25076,n25077,n25078 );
   nor U24634 ( n25078,n25079,n25046,n25080 );
   nor U24635 ( n25080,n25038,n25041 );
   not U24636 ( n25041,n25045 );
   not U24637 ( n25077,n25081 );
   nor U24638 ( n25074,n23622,n24401 );
   and U24639 ( n25073,n25082,n24474 );
   nor U24640 ( n25072,n23622,n24394 );
   nor U24641 ( n25070,n25083,n25084 );
   nor U24642 ( n25084,n23650,n23608 );
   nor U24643 ( n25083,n25085,n24347 );
   xor U24644 ( n25085,n25086,n25079 );
   nand U24645 ( n25069,n24672,n25082 );
   nand U24646 ( n25082,n25087,n25081 );
   nand U24647 ( n25081,n25086,n25079 );
   or U24648 ( n25087,n25079,n25086 );
   nor U24649 ( n25086,n25039,n25038 );
   nand U24650 ( n25068,n25012,n25088 );
   and U24651 ( n25063,n24011,p1_reg2_reg_27_ );
   nand U24652 ( n25061,n24283,n23381 );
   not U24653 ( n24283,n24303 );
   nand U24654 ( n25060,n24009,n23623 );
   xor U24655 ( n23623,n23636,n25089 );
   nand U24656 ( n25059,n24006,n25088 );
   not U24657 ( n25088,n23622 );
   xor U24658 ( n23622,n25079,n25090 );
   nand U24659 ( n25090,n25091,n25092,n25093 );
   nand U24660 ( n25091,n25094,n25054,n25095 );
   nand U24661 ( p1_u3265,n25096,n25097,n25098,n25099 );
   nor U24662 ( n25099,n25100,n25101,n25102,n25103 );
   and U24663 ( n25103,n23612,n24006 );
   not U24664 ( n24006,n24449 );
   nor U24665 ( n25102,n23605,n24303 );
   nand U24666 ( n24303,n24012,n23626 );
   nor U24667 ( n25101,n23607,n24295 );
   nand U24668 ( n24295,n24012,n24036 );
   not U24669 ( n24036,n23608 );
   and U24670 ( n25100,n24009,n23611,n23610 );
   nand U24671 ( n23610,n23609,n25107 );
   nand U24672 ( n25107,n25108,n23625 );
   nor U24673 ( n25098,n25109,n25110 );
   nor U24674 ( n25110,n24035,n24281 );
   nor U24675 ( n25109,n25111,n24302 );
   nand U24676 ( n25097,p1_reg2_reg_28_,n24011 );
   nand U24677 ( n25096,n24012,n23602 );
   nand U24678 ( n23602,n25113,n25114 );
   nand U24679 ( n25114,n23612,n25115 );
   nand U24680 ( n25115,n25116,n24395 );
   xor U24681 ( n23612,n25117,n25118 );
   nor U24682 ( n25117,n24022,n24023 );
   nand U24683 ( n24023,n25119,n25120,n25121 );
   nand U24684 ( n25121,n23387,n25122,n25047 );
   nand U24685 ( n25119,n25095,n25122,n25094,n25054 );
   nand U24686 ( n25095,n25052,n25058 );
   nor U24687 ( n24022,n25092,n25123 );
   nand U24688 ( n25092,n25124,n25056,n25094,n25054 );
   not U24689 ( n25124,n24992 );
   nand U24690 ( n24992,n25125,n25126 );
   nand U24691 ( n25126,n23665,n25127 );
   or U24692 ( n25127,n24980,n23682 );
   nand U24693 ( n25125,n23682,n24980 );
   nand U24694 ( n24980,n25128,n25129 );
   nand U24695 ( n25129,n24963,n25130 );
   nand U24696 ( n25130,n24934,n24933 );
   or U24697 ( n25128,n24933,n24934 );
   nand U24698 ( n24933,n25131,n25132,n25133 );
   nand U24699 ( n25133,n25134,n25135 );
   nand U24700 ( n25135,n24921,n25136 );
   nand U24701 ( n25136,n24922,n24882 );
   not U24702 ( n24921,n24918 );
   nand U24703 ( n24918,n24881,n25137 );
   nand U24704 ( n25137,n25138,n25139 );
   not U24705 ( n25138,n24883 );
   nand U24706 ( n25131,n24882,n25134,n24923 );
   and U24707 ( n24923,n25140,n24829 );
   nand U24708 ( n24829,n25141,n25142 );
   nand U24709 ( n25142,n25143,n25144 );
   nand U24710 ( n25143,n24808,n24807 );
   nand U24711 ( n24807,n24779,n24811 );
   not U24712 ( n24779,n24812 );
   nand U24713 ( n24812,n25145,n25146 );
   nand U24714 ( n25146,n23795,n25147 );
   nand U24715 ( n25147,n24724,n24726 );
   not U24716 ( n24724,n25148 );
   nand U24717 ( n25145,n23782,n25148 );
   nand U24718 ( n25148,n25149,n25150 );
   nand U24719 ( n25150,n23781,n25151 );
   nand U24720 ( n25151,n23799,n24699 );
   or U24721 ( n25149,n24699,n23799 );
   nand U24722 ( n24699,n25152,n25153 );
   nand U24723 ( n25153,n25154,n24681,n24685 );
   and U24724 ( n24685,n24629,n25155 );
   nand U24725 ( n25155,n23820,n23835 );
   nand U24726 ( n24629,n25156,n25157 );
   nand U24727 ( n25157,n25158,n25159 );
   nand U24728 ( n25158,n24583,n24582 );
   nand U24729 ( n24582,n24586,n24587 );
   nand U24730 ( n24587,n25160,n25161 );
   nand U24731 ( n25160,n24528,n25162 );
   nand U24732 ( n24528,n25163,n25164 );
   nand U24733 ( n25164,n25165,n25166 );
   nand U24734 ( n25166,n24516,n23885 );
   nand U24735 ( n25165,n24486,n24485 );
   nand U24736 ( n24485,n24490,n24489 );
   nand U24737 ( n24490,n25167,n25168,n25169 );
   nand U24738 ( n25169,n24416,n24412 );
   nand U24739 ( n25168,n24376,n25170,n25171 );
   nand U24740 ( n25171,n23920,n23908 );
   nand U24741 ( n24376,n25172,n25173,n25174 );
   nand U24742 ( n25174,n25175,n23934 );
   nand U24743 ( n25173,n25176,n24359,n24319 );
   and U24744 ( n24319,n24293,n25177 );
   nand U24745 ( n25177,n23946,n23961 );
   nand U24746 ( n25176,n23918,n24340 );
   nand U24747 ( n25172,n25178,n23456 );
   nand U24748 ( n25178,n24357,n24340 );
   not U24749 ( n24357,n25175 );
   nand U24750 ( n25175,n25179,n25180 );
   nand U24751 ( n25180,n24320,n24359 );
   nand U24752 ( n25167,n25181,n23450 );
   or U24753 ( n25181,n24412,n24416 );
   nand U24754 ( n25163,n24482,n23444 );
   nand U24755 ( n25152,n25154,n25182 );
   nand U24756 ( n25182,n25183,n24680,n25184 );
   nand U24757 ( n25183,n24686,n24681 );
   nand U24758 ( n25140,n25185,n24822 );
   and U24759 ( n24882,n24886,n25139 );
   nand U24760 ( n25113,n25186,n24327 );
   nand U24761 ( n24327,n24403,n24347,n24397,n24400 );
   xor U24762 ( n25186,n25118,n24034 );
   nand U24763 ( n24034,n25187,n25188 );
   nand U24764 ( n25188,n25189,n25190 );
   nand U24765 ( n25190,n23607,n25089 );
   or U24766 ( n25189,n25038,n25039 );
   nor U24767 ( n25039,n25045,n25046 );
   nor U24768 ( n25046,n23387,n23638 );
   nand U24769 ( n25045,n25191,n25192 );
   nand U24770 ( n25192,n23667,n25193 );
   or U24771 ( n25193,n25014,n25194 );
   nand U24772 ( n25191,n25014,n25194 );
   nand U24773 ( n25014,n25195,n25196 );
   nand U24774 ( n25196,n23648,n25197 );
   nand U24775 ( n25197,n23666,n24997 );
   or U24776 ( n25195,n24997,n23666 );
   nand U24777 ( n24997,n25198,n25199 );
   nand U24778 ( n25199,n25200,n24942,n24915 );
   nor U24779 ( n24915,n24904,n24906 );
   nor U24780 ( n24906,n23402,n23707 );
   nand U24781 ( n24904,n25201,n25202 );
   nand U24782 ( n25202,n23728,n25203 );
   or U24783 ( n25203,n24875,n24876 );
   nand U24784 ( n25201,n24875,n24876 );
   nand U24785 ( n24875,n25204,n25205 );
   nand U24786 ( n25205,n23744,n25206 );
   or U24787 ( n25206,n24849,n23729 );
   nand U24788 ( n25204,n24849,n23729 );
   nand U24789 ( n24849,n25207,n25208 );
   nand U24790 ( n25208,n25185,n25209 );
   or U24791 ( n25209,n24827,n23745 );
   nand U24792 ( n25207,n24827,n23745 );
   nand U24793 ( n24827,n25210,n25211 );
   nand U24794 ( n25211,n23741,n25212 );
   nand U24795 ( n25212,n23759,n24801 );
   or U24796 ( n25210,n24801,n23759 );
   nand U24797 ( n24801,n25213,n25214 );
   nand U24798 ( n25214,n24775,n25215 );
   nand U24799 ( n25215,n24774,n25216 );
   nand U24800 ( n25216,n24768,n24732 );
   not U24801 ( n24768,n24710 );
   nand U24802 ( n24710,n24703,n23423 );
   and U24803 ( n24774,n24731,n25217 );
   nand U24804 ( n25217,n24745,n23417 );
   nand U24805 ( n24731,n23782,n23420 );
   nand U24806 ( n25213,n24775,n24732,n24709 );
   and U24807 ( n24709,n24715,n24714 );
   nand U24808 ( n24714,n23781,n23799 );
   not U24809 ( n23781,n23423 );
   not U24810 ( n24715,n24713 );
   nand U24811 ( n24713,n25218,n25219 );
   nand U24812 ( n25219,n23796,n25220 );
   nand U24813 ( n25220,n24673,n23810 );
   not U24814 ( n24673,n25221 );
   nand U24815 ( n25218,n25221,n24676 );
   nand U24816 ( n25221,n25222,n25223 );
   nand U24817 ( n25223,n24670,n25224 );
   nand U24818 ( n25224,n24639,n24649 );
   or U24819 ( n25222,n24649,n24639 );
   nand U24820 ( n24649,n25225,n25226 );
   nand U24821 ( n25226,n24626,n25227 );
   nand U24822 ( n25227,n24625,n25228 );
   nand U24823 ( n25228,n24619,n24573 );
   not U24824 ( n24619,n24548 );
   nand U24825 ( n24548,n23858,n23438 );
   and U24826 ( n24625,n24572,n25229 );
   nand U24827 ( n25229,n23835,n23432 );
   nand U24828 ( n24572,n23847,n23435 );
   nand U24829 ( n25225,n24626,n24573,n24618 );
   and U24830 ( n24618,n24545,n24547 );
   nand U24831 ( n24547,n25230,n25231 );
   nand U24832 ( n24545,n25232,n25233 );
   nand U24833 ( n25233,n25234,n23441 );
   nand U24834 ( n25234,n24509,n24525 );
   nand U24835 ( n25232,n23874,n24522 );
   not U24836 ( n24522,n24509 );
   nor U24837 ( n24509,n25235,n24477 );
   nor U24838 ( n24477,n24480,n25236 );
   nor U24839 ( n25236,n23444,n23885 );
   nand U24840 ( n24480,n25237,n24443 );
   nand U24841 ( n24443,n25238,n24407,n25239 );
   nand U24842 ( n25239,n23897,n23447 );
   nand U24843 ( n24407,n23908,n23450 );
   nand U24844 ( n25238,n24406,n24408 );
   nand U24845 ( n24408,n25240,n25241 );
   nand U24846 ( n25241,n25242,n24371 );
   nand U24847 ( n24371,n25243,n25244 );
   nand U24848 ( n25244,n24353,n25245 );
   nand U24849 ( n25245,n23918,n23934 );
   nand U24850 ( n24353,n24317,n24329 );
   nand U24851 ( n24329,n25246,n24318 );
   nand U24852 ( n24318,n23962,n24321 );
   not U24853 ( n25246,n24330 );
   nand U24854 ( n24330,n25247,n25248 );
   nand U24855 ( n25248,n23946,n25249 );
   nand U24856 ( n25249,n23961,n24276 );
   nand U24857 ( n25247,n24298,n24296 );
   not U24858 ( n24298,n24276 );
   nand U24859 ( n24276,n23960,n23974 );
   nand U24860 ( n24317,n23947,n23459 );
   nand U24861 ( n25243,n24340,n23456 );
   nand U24862 ( n25242,n23933,n24372 );
   nand U24863 ( n25240,n23919,n23453 );
   nand U24864 ( n24406,n23920,n24412 );
   not U24865 ( n25237,n24444 );
   nor U24866 ( n24444,n23447,n23897 );
   not U24867 ( n25235,n24478 );
   nand U24868 ( n24478,n23885,n23444 );
   nand U24869 ( n24573,n23859,n24578 );
   nand U24870 ( n24626,n23820,n24628 );
   nand U24871 ( n24732,n23795,n24726 );
   nand U24872 ( n24775,n23783,n23766 );
   nand U24873 ( n25198,n25250,n25200 );
   nand U24874 ( n25200,n23665,n24979 );
   nand U24875 ( n25250,n25251,n24941,n25252 );
   nand U24876 ( n25252,n23682,n23396 );
   nand U24877 ( n24941,n23693,n23399 );
   nand U24878 ( n25251,n24905,n24942 );
   nand U24879 ( n24942,n24963,n24934 );
   not U24880 ( n24905,n24916 );
   nand U24881 ( n24916,n23707,n23402 );
   nor U24882 ( n25038,n25047,n23650 );
   nand U24883 ( n25187,n23625,n23384 );
   nand U24884 ( p1_u3264,n25253,n25254,n25255,n25256 );
   nand U24885 ( n25255,n23583,n23584,n24009 );
   nand U24886 ( n23583,n23582,n25257 );
   or U24887 ( n25257,n23611,n23594 );
   nand U24888 ( n25254,n24010,n23582 );
   nand U24889 ( n25253,p1_reg2_reg_30_,n24011 );
   nand U24890 ( p1_u3263,n25258,n25259,n25260,n25256 );
   or U24891 ( n25256,n23571,n24011 );
   nand U24892 ( n23571,n24037,n23372 );
   nand U24893 ( n24037,n25261,n25262 );
   nand U24894 ( n25262,n23626,n25263 );
   not U24895 ( n23626,n23606 );
   nand U24896 ( n25261,n25265,n25105 );
   nand U24897 ( n25260,n24009,n23576 );
   xor U24898 ( n23576,n23584,n23574 );
   or U24899 ( n23584,n23582,n23594,n23611 );
   nand U24900 ( n23611,n23625,n24035,n25108 );
   not U24901 ( n25108,n23636 );
   nand U24902 ( n23636,n23649,n23638,n25015 );
   not U24903 ( n25015,n23670 );
   nand U24904 ( n23670,n23666,n23682,n24996 );
   not U24905 ( n24996,n23696 );
   nand U24906 ( n23696,n23707,n23693,n24936 );
   not U24907 ( n24936,n23717 );
   nand U24908 ( n23717,n23719,n24842,n24851 );
   not U24909 ( n24851,n24830 );
   nand U24910 ( n24830,n23759,n24822,n24833 );
   not U24911 ( n24833,n23770 );
   nand U24912 ( n23770,n24745,n23782,n24778 );
   not U24913 ( n24778,n24695 );
   nand U24914 ( n24695,n23810,n24703,n24698 );
   not U24915 ( n24698,n24643 );
   nand U24916 ( n24643,n23835,n24639,n24646 );
   not U24917 ( n24646,n23845 );
   nand U24918 ( n23845,n23847,n23858,n24549 );
   not U24919 ( n24549,n23872 );
   nand U24920 ( n23872,n23885,n23874,n24527 );
   not U24921 ( n24527,n23895 );
   nand U24922 ( n23895,n23908,n23897,n24448 );
   not U24923 ( n24448,n23923 );
   nand U24924 ( n23923,n24340,n23919,n24355 );
   not U24925 ( n24355,n23950 );
   nand U24926 ( n23950,n23961,n24278,n23947 );
   not U24927 ( n24340,n23934 );
   not U24928 ( n23908,n24412 );
   not U24929 ( n23885,n24482 );
   not U24930 ( n24703,n23799 );
   not U24931 ( n23782,n24726 );
   not U24932 ( n23682,n24979 );
   not U24933 ( n23625,n25089 );
   nand U24934 ( n24282,n25266,n24012 );
   nand U24935 ( n25259,n24010,n23574 );
   not U24936 ( n24010,n24281 );
   nand U24937 ( n25258,p1_reg2_reg_31_,n24011 );
   nand U24938 ( n25268,n25269,n25270 );
   nand U24939 ( n25270,n25271,n23983,n25272,n23980 );
   nand U24940 ( p1_u3262,n25273,n25274,n25275,n25276 );
   nor U24941 ( n25276,n25277,n25278 );
   nor U24942 ( n25277,n15117,n25279 );
   not U24943 ( n15117,p1_addr_reg_19_ );
   nand U24944 ( n25275,n25280,n23979 );
   nand U24945 ( n25274,n25281,n25282,n25283 );
   nand U24946 ( n25282,n25284,n25285,n25286 );
   xor U24947 ( n25286,p1_reg1_reg_19_,n23979 );
   nand U24948 ( n25285,n25287,n25288 );
   nand U24949 ( n25281,n25287,n25289,n25290 );
   xor U24950 ( n25290,n25291,p1_reg1_reg_19_ );
   nand U24951 ( n25289,p1_reg1_reg_18_,n25284 );
   nand U24952 ( n25284,n25292,n25293 );
   nand U24953 ( n25287,n25294,n25295 );
   nand U24954 ( n25273,n25296,n25297,n25298 );
   nand U24955 ( n25297,n25299,n25300,n25301 );
   xor U24956 ( n25301,p1_reg2_reg_19_,n23979 );
   nand U24957 ( n25300,n25302,n24821 );
   nand U24958 ( n25296,n25302,n25303,n25304 );
   xor U24959 ( n25304,n23979,n24850 );
   not U24960 ( n24850,p1_reg2_reg_19_ );
   nand U24961 ( n25303,p1_reg2_reg_18_,n25299 );
   nand U24962 ( n25299,n25305,n25293 );
   not U24963 ( n25305,n25306 );
   nand U24964 ( n25302,n25294,n25306 );
   nand U24965 ( p1_u3261,n25307,n25308,n25309,n25310 );
   nand U24966 ( n25310,n25294,n25311 );
   nand U24967 ( n25311,n25312,n25313,n25314 );
   nand U24968 ( n25314,n25298,n25315 );
   xor U24969 ( n25315,n25306,n24821 );
   not U24970 ( n24821,p1_reg2_reg_18_ );
   nand U24971 ( n25312,n25283,n25316 );
   xor U24972 ( n25316,p1_reg1_reg_18_,n25292 );
   nand U24973 ( n25309,n25317,n25293 );
   nand U24974 ( n25317,n25318,n25319 );
   nand U24975 ( n25319,n25320,n25283 );
   xor U24976 ( n25320,n25292,n25288 );
   not U24977 ( n25288,p1_reg1_reg_18_ );
   not U24978 ( n25292,n25295 );
   nand U24979 ( n25295,n25321,n25322,n25323 );
   nand U24980 ( n25323,n25324,n25325 );
   nand U24981 ( n25322,p1_reg1_reg_17_,n25326 );
   nand U24982 ( n25326,n25327,n25328 );
   or U24983 ( n25321,n25328,n25327 );
   nand U24984 ( n25318,n25329,n25298 );
   xor U24985 ( n25329,p1_reg2_reg_18_,n25306 );
   nand U24986 ( n25306,n25330,n25331,n25332 );
   nand U24987 ( n25332,n25333,n25334 );
   nand U24988 ( n25331,p1_reg2_reg_17_,n25335 );
   nand U24989 ( n25335,n25327,n25336 );
   or U24990 ( n25330,n25336,n25327 );
   nand U24991 ( n25308,n25337,p1_addr_reg_18_ );
   nand U24992 ( n25307,p1_reg3_reg_18_,p1_u3086 );
   nand U24993 ( p1_u3260,n25338,n25339,n25340,n25341 );
   nor U24994 ( n25341,n25342,n25343 );
   nor U24995 ( n25342,n15128,n25279 );
   not U24996 ( n15128,p1_addr_reg_17_ );
   nand U24997 ( n25340,n25280,n25344 );
   nand U24998 ( n25339,n25345,n25346,n25283 );
   nand U24999 ( n25346,n25347,n25348,n25325 );
   and U25000 ( n25325,n25349,n25350 );
   or U25001 ( n25349,n25344,p1_reg1_reg_17_ );
   nand U25002 ( n25348,n25351,n25328 );
   nand U25003 ( n25347,n25344,p1_reg1_reg_17_ );
   nand U25004 ( n25345,n25352,n25328,n25353 );
   xor U25005 ( n25353,p1_reg1_reg_17_,n25327 );
   nand U25006 ( n25328,n25354,p1_reg1_reg_16_ );
   nand U25007 ( n25352,n25324,n25350 );
   nand U25008 ( n25350,n25355,n25356 );
   not U25009 ( n25324,n25351 );
   nand U25010 ( n25338,n25357,n25358,n25298 );
   nand U25011 ( n25358,n25359,n25360,n25334 );
   and U25012 ( n25334,n25361,n25362 );
   nand U25013 ( n25361,n25327,n24803 );
   not U25014 ( n24803,p1_reg2_reg_17_ );
   nand U25015 ( n25360,n25363,n25336 );
   nand U25016 ( n25359,n25344,p1_reg2_reg_17_ );
   nand U25017 ( n25357,n25364,n25336,n25365 );
   xor U25018 ( n25365,p1_reg2_reg_17_,n25327 );
   nand U25019 ( n25336,n25354,p1_reg2_reg_16_ );
   nand U25020 ( n25364,n25333,n25362 );
   nand U25021 ( n25362,n25355,n24776 );
   not U25022 ( n25333,n25363 );
   nand U25023 ( p1_u3259,n25366,n25367,n25368,n25369 );
   nand U25024 ( n25369,n25355,n25370 );
   nand U25025 ( n25370,n25371,n25372 );
   nand U25026 ( n25372,n25283,n25373 );
   xor U25027 ( n25373,n25351,n25356 );
   not U25028 ( n25356,p1_reg1_reg_16_ );
   nand U25029 ( n25371,n25298,n25374 );
   xor U25030 ( n25374,n25363,n24776 );
   not U25031 ( n24776,p1_reg2_reg_16_ );
   nand U25032 ( n25368,n25354,n25375 );
   nand U25033 ( n25375,n25376,n25313,n25377 );
   nand U25034 ( n25377,n25378,n25298 );
   xor U25035 ( n25378,p1_reg2_reg_16_,n25363 );
   nand U25036 ( n25363,n25379,n25380 );
   nand U25037 ( n25380,n25381,n24735 );
   or U25038 ( n25381,n25382,n25383 );
   nand U25039 ( n25379,n25383,n25382 );
   nand U25040 ( n25376,n25384,n25283 );
   xor U25041 ( n25384,p1_reg1_reg_16_,n25351 );
   nand U25042 ( n25351,n25385,n25386 );
   nand U25043 ( n25386,n25387,n25388 );
   or U25044 ( n25387,n25389,n25383 );
   nand U25045 ( n25385,n25383,n25389 );
   nand U25046 ( n25367,n25337,p1_addr_reg_16_ );
   nand U25047 ( n25366,p1_reg3_reg_16_,p1_u3086 );
   nand U25048 ( p1_u3258,n25390,n25391,n25392,n25393 );
   nand U25049 ( n25393,n25394,n25395 );
   nand U25050 ( n25395,n25396,n25313,n25397 );
   nand U25051 ( n25397,n25398,n25298 );
   xor U25052 ( n25398,p1_reg2_reg_15_,n25382 );
   nand U25053 ( n25396,n25399,n25283 );
   xor U25054 ( n25399,p1_reg1_reg_15_,n25389 );
   nand U25055 ( n25392,n25383,n25400 );
   nand U25056 ( n25400,n25401,n25402 );
   nand U25057 ( n25402,n25283,n25403 );
   xor U25058 ( n25403,n25389,n25388 );
   not U25059 ( n25388,p1_reg1_reg_15_ );
   nand U25060 ( n25389,n25404,n25405 );
   nand U25061 ( n25405,n25406,n25407 );
   or U25062 ( n25406,n25408,n25409 );
   nand U25063 ( n25404,n25409,n25408 );
   nand U25064 ( n25401,n25298,n25410 );
   xor U25065 ( n25410,n25382,n24735 );
   not U25066 ( n24735,p1_reg2_reg_15_ );
   nand U25067 ( n25382,n25411,n25412 );
   nand U25068 ( n25412,n25413,n25414 );
   or U25069 ( n25413,n25415,n25409 );
   nand U25070 ( n25411,n25409,n25415 );
   nand U25071 ( n25391,n25337,p1_addr_reg_15_ );
   nand U25072 ( n25390,p1_reg3_reg_15_,p1_u3086 );
   nand U25073 ( p1_u3257,n25416,n25417,n25418,n25419 );
   nand U25074 ( n25419,n25409,n25420 );
   nand U25075 ( n25420,n25421,n25422 );
   nand U25076 ( n25422,n25283,n25423 );
   xor U25077 ( n25423,n25408,n25407 );
   not U25078 ( n25407,p1_reg1_reg_14_ );
   nand U25079 ( n25421,n25298,n25424 );
   xor U25080 ( n25424,n25414,n25415 );
   not U25081 ( n25414,p1_reg2_reg_14_ );
   nand U25082 ( n25418,n25425,n25426 );
   nand U25083 ( n25426,n25427,n25313,n25428 );
   nand U25084 ( n25428,n25429,n25298 );
   xor U25085 ( n25429,n25415,p1_reg2_reg_14_ );
   nand U25086 ( n25415,n25430,n25431 );
   nand U25087 ( n25430,n25432,n25433,n25434 );
   nand U25088 ( n25427,n25435,n25283 );
   xor U25089 ( n25435,p1_reg1_reg_14_,n25408 );
   nand U25090 ( n25408,n25436,n25437 );
   nand U25091 ( n25436,n25438,n25439,n25440 );
   nand U25092 ( n25417,n25337,p1_addr_reg_14_ );
   nand U25093 ( n25416,p1_reg3_reg_14_,p1_u3086 );
   nand U25094 ( p1_u3256,n25441,n25442,n25443,n25444 );
   nor U25095 ( n25444,n25445,n25446 );
   nor U25096 ( n25445,n15142,n25279 );
   not U25097 ( n15142,p1_addr_reg_13_ );
   nand U25098 ( n25443,n25280,n25447 );
   nand U25099 ( n25442,n25448,n25449,n25283 );
   nand U25100 ( n25449,n25440,n25450,n25451,n25437 );
   or U25101 ( n25437,p1_reg1_reg_13_,n25447 );
   nand U25102 ( n25450,n25452,n25439 );
   nand U25103 ( n25440,n25447,p1_reg1_reg_13_ );
   nand U25104 ( n25448,n25438,n25439,n25453 );
   xor U25105 ( n25453,p1_reg1_reg_13_,n25454 );
   nand U25106 ( n25441,n25455,n25456,n25298 );
   nand U25107 ( n25456,n25434,n25457,n25458,n25431 );
   nand U25108 ( n25431,n24675,n25454 );
   not U25109 ( n24675,p1_reg2_reg_13_ );
   nand U25110 ( n25457,n25459,n25433 );
   nand U25111 ( n25434,n25447,p1_reg2_reg_13_ );
   nand U25112 ( n25455,n25432,n25433,n25460 );
   xor U25113 ( n25460,p1_reg2_reg_13_,n25454 );
   nand U25114 ( p1_u3255,n25461,n25462,n25463,n25464 );
   nor U25115 ( n25464,n25465,n25466 );
   nor U25116 ( n25465,n15147,n25279 );
   not U25117 ( n15147,p1_addr_reg_12_ );
   nand U25118 ( n25463,n25467,n25468 );
   nand U25119 ( n25468,n25469,n25313,n25470 );
   nand U25120 ( n25470,p1_reg2_reg_12_,n25471,n25298 );
   nand U25121 ( n25469,p1_reg1_reg_12_,n25472,n25283 );
   nand U25122 ( n25462,n25473,n25438,n25283 );
   nand U25123 ( n25438,n25451,n25472 );
   nand U25124 ( n25473,n25452,n25474 );
   nand U25125 ( n25474,n25439,n25451 );
   or U25126 ( n25451,n25467,p1_reg1_reg_12_ );
   nand U25127 ( n25439,n25467,p1_reg1_reg_12_ );
   not U25128 ( n25452,n25472 );
   nand U25129 ( n25472,n25475,n25476 );
   nand U25130 ( n25476,n25477,n25478 );
   nand U25131 ( n25478,n25479,n25480 );
   nand U25132 ( n25475,n25481,p1_reg1_reg_11_ );
   nand U25133 ( n25461,n25482,n25432,n25298 );
   nand U25134 ( n25432,n25458,n25471 );
   nand U25135 ( n25482,n25459,n25483 );
   nand U25136 ( n25483,n25433,n25458 );
   nand U25137 ( n25458,n25484,n24638 );
   not U25138 ( n24638,p1_reg2_reg_12_ );
   nand U25139 ( n25433,n25467,p1_reg2_reg_12_ );
   not U25140 ( n25459,n25471 );
   nand U25141 ( n25471,n25485,n25486 );
   nand U25142 ( n25486,n25487,n25488 );
   nand U25143 ( n25488,n25479,n24627 );
   nand U25144 ( n25485,n25481,p1_reg2_reg_11_ );
   nand U25145 ( p1_u3254,n25489,n25490,n25491,n25492 );
   nand U25146 ( n25492,n25479,n25493 );
   nand U25147 ( n25493,n25494,n25495 );
   nand U25148 ( n25495,n25283,n25496 );
   xor U25149 ( n25496,n25477,p1_reg1_reg_11_ );
   nand U25150 ( n25494,n25298,n25497 );
   xor U25151 ( n25497,n25487,p1_reg2_reg_11_ );
   nand U25152 ( n25491,n25481,n25498 );
   nand U25153 ( n25498,n25499,n25313,n25500 );
   nand U25154 ( n25500,n25501,n25298 );
   xor U25155 ( n25501,n24627,n25487 );
   and U25156 ( n25487,n25502,n25503 );
   nand U25157 ( n25502,n25504,n25505,n25506 );
   not U25158 ( n24627,p1_reg2_reg_11_ );
   nand U25159 ( n25499,n25507,n25283 );
   xor U25160 ( n25507,n25480,n25477 );
   and U25161 ( n25477,n25508,n25509 );
   nand U25162 ( n25508,n25510,n25511,n25512 );
   not U25163 ( n25480,p1_reg1_reg_11_ );
   nand U25164 ( n25490,n25337,p1_addr_reg_11_ );
   nand U25165 ( n25489,p1_reg3_reg_11_,p1_u3086 );
   nand U25166 ( p1_u3253,n25513,n25514,n25515,n25516 );
   nor U25167 ( n25516,n25517,n25518 );
   nor U25168 ( n25517,n15155,n25279 );
   not U25169 ( n15155,p1_addr_reg_10_ );
   nand U25170 ( n25515,n25280,n25519 );
   nand U25171 ( n25514,n25520,n25521,n25283 );
   nand U25172 ( n25521,n25512,n25522,n25523,n25509 );
   or U25173 ( n25509,n25519,p1_reg1_reg_10_ );
   nand U25174 ( n25512,n25519,p1_reg1_reg_10_ );
   nand U25175 ( n25520,n25510,n25511,n25524 );
   xor U25176 ( n25524,p1_reg1_reg_10_,n25525 );
   nand U25177 ( n25510,n25523,n25526 );
   nand U25178 ( n25513,n25527,n25528,n25298 );
   nand U25179 ( n25528,n25506,n25529,n25530,n25503 );
   nand U25180 ( n25503,n25525,n24577 );
   not U25181 ( n24577,p1_reg2_reg_10_ );
   nand U25182 ( n25506,n25519,p1_reg2_reg_10_ );
   nand U25183 ( n25527,n25504,n25505,n25531 );
   xor U25184 ( n25531,p1_reg2_reg_10_,n25525 );
   nand U25185 ( n25504,n25530,n25532 );
   nand U25186 ( p1_u3252,n25533,n25534,n25535,n25536 );
   nor U25187 ( n25536,n25537,n25538 );
   nor U25188 ( n25537,n15092,n25279 );
   not U25189 ( n15092,p1_addr_reg_9_ );
   nand U25190 ( n25535,n25539,n25540 );
   nand U25191 ( n25540,n25541,n25313,n25542 );
   nand U25192 ( n25542,p1_reg2_reg_9_,n25532,n25298 );
   nand U25193 ( n25541,p1_reg1_reg_9_,n25526,n25283 );
   nand U25194 ( n25534,n25543,n25544,n25283 );
   nand U25195 ( n25544,n25545,n25546 );
   nand U25196 ( n25543,n25522,n25523 );
   not U25197 ( n25523,n25545 );
   nor U25198 ( n25545,n25539,p1_reg1_reg_9_ );
   nand U25199 ( n25522,n25546,n25511 );
   nand U25200 ( n25511,n25539,p1_reg1_reg_9_ );
   not U25201 ( n25546,n25526 );
   nand U25202 ( n25526,n25547,n25548 );
   nand U25203 ( n25547,n25549,n25550 );
   nand U25204 ( n25533,n25551,n25552,n25298 );
   nand U25205 ( n25552,n25553,n25554 );
   nand U25206 ( n25551,n25529,n25530 );
   not U25207 ( n25530,n25553 );
   nor U25208 ( n25553,n25539,p1_reg2_reg_9_ );
   nand U25209 ( n25529,n25554,n25505 );
   nand U25210 ( n25505,n25539,p1_reg2_reg_9_ );
   not U25211 ( n25554,n25532 );
   nand U25212 ( n25532,n25555,n25556 );
   nand U25213 ( n25555,n25557,n25558 );
   nand U25214 ( p1_u3251,n25559,n25560,n25561,n25562 );
   nor U25215 ( n25562,n25563,n25564 );
   nor U25216 ( n25563,n15089,n25279 );
   not U25217 ( n15089,p1_addr_reg_8_ );
   nand U25218 ( n25561,n25280,n25565 );
   or U25219 ( n25560,n25566,n25567 );
   xor U25220 ( n25566,n25550,n25568 );
   nand U25221 ( n25568,n25549,n25548 );
   nand U25222 ( n25548,n25565,p1_reg1_reg_8_ );
   or U25223 ( n25549,n25565,p1_reg1_reg_8_ );
   nand U25224 ( n25550,n25569,n25570 );
   nand U25225 ( n25570,p1_reg1_reg_7_,n25571 );
   nand U25226 ( n25571,n25572,n25573 );
   nand U25227 ( n25569,n25574,n25575 );
   nand U25228 ( n25559,n25576,n25298 );
   xor U25229 ( n25576,n25577,n25558 );
   nand U25230 ( n25558,n25578,n25579 );
   nand U25231 ( n25579,p1_reg2_reg_7_,n25580 );
   nand U25232 ( n25580,n25581,n25573 );
   nand U25233 ( n25578,n25574,n25582 );
   and U25234 ( n25577,n25556,n25557 );
   nand U25235 ( n25557,n25583,n24524 );
   not U25236 ( n24524,p1_reg2_reg_8_ );
   nand U25237 ( n25556,n25565,p1_reg2_reg_8_ );
   nand U25238 ( p1_u3250,n25584,n25585,n25586,n25587 );
   nor U25239 ( n25587,n25588,n25589 );
   nor U25240 ( n25588,n15086,n25279 );
   not U25241 ( n15086,p1_addr_reg_7_ );
   nand U25242 ( n25586,n25574,n25590 );
   nand U25243 ( n25590,n25591,n25313,n25592 );
   nand U25244 ( n25592,n25593,n24481,n25298 );
   not U25245 ( n24481,p1_reg2_reg_7_ );
   nand U25246 ( n25591,n25594,n25595,n25283 );
   not U25247 ( n25595,p1_reg1_reg_7_ );
   nand U25248 ( n25585,n25596,n25594,n25283 );
   nand U25249 ( n25594,n25597,n25598,n25599 );
   xor U25250 ( n25599,p1_reg1_reg_7_,n25574 );
   nand U25251 ( n25597,n25600,n25601 );
   nand U25252 ( n25596,n25572,n25602 );
   nand U25253 ( n25602,n25573,p1_reg1_reg_7_ );
   not U25254 ( n25572,n25575 );
   nand U25255 ( n25575,n25601,n25603 );
   nand U25256 ( n25584,n25604,n25593,n25298 );
   nand U25257 ( n25593,n25605,n25606,n25607 );
   xor U25258 ( n25607,p1_reg2_reg_7_,n25574 );
   nand U25259 ( n25605,n25608,n25609 );
   nand U25260 ( n25604,n25581,n25610 );
   nand U25261 ( n25610,n25573,p1_reg2_reg_7_ );
   not U25262 ( n25581,n25582 );
   nand U25263 ( n25582,n25609,n25611 );
   nand U25264 ( p1_u3249,n25612,n25613,n25614,n25615 );
   nor U25265 ( n25615,n25616,n25617 );
   nor U25266 ( n25616,n15168,n25279 );
   not U25267 ( n15168,p1_addr_reg_6_ );
   nand U25268 ( n25614,n25618,n25619 );
   nand U25269 ( n25619,n25620,n25313,n25621 );
   nand U25270 ( n25621,p1_reg2_reg_6_,n25622,n25298 );
   nand U25271 ( n25620,p1_reg1_reg_6_,n25623,n25283 );
   nand U25272 ( n25613,n25624,n25603,n25283 );
   nand U25273 ( n25603,n25623,n25598 );
   nand U25274 ( n25624,n25600,n25625 );
   nand U25275 ( n25625,n25601,n25598 );
   or U25276 ( n25598,n25618,p1_reg1_reg_6_ );
   nand U25277 ( n25601,n25618,p1_reg1_reg_6_ );
   not U25278 ( n25600,n25623 );
   nand U25279 ( n25623,n25626,n25627 );
   nand U25280 ( n25627,p1_reg1_reg_5_,n25628 );
   nand U25281 ( n25628,n25629,n25630 );
   nand U25282 ( n25626,n25631,n25632 );
   nand U25283 ( n25612,n25633,n25611,n25298 );
   nand U25284 ( n25611,n25622,n25606 );
   nand U25285 ( n25633,n25608,n25634 );
   nand U25286 ( n25634,n25609,n25606 );
   nand U25287 ( n25606,n25635,n24445 );
   not U25288 ( n24445,p1_reg2_reg_6_ );
   nand U25289 ( n25609,n25618,p1_reg2_reg_6_ );
   not U25290 ( n25608,n25622 );
   nand U25291 ( n25622,n25636,n25637 );
   nand U25292 ( n25637,p1_reg2_reg_5_,n25638 );
   nand U25293 ( n25638,n25639,n25630 );
   nand U25294 ( n25636,n25631,n25640 );
   nand U25295 ( p1_u3248,n25641,n25642,n25643,n25644 );
   nor U25296 ( n25644,n25645,n25646 );
   nor U25297 ( n25645,n15172,n25279 );
   not U25298 ( n15172,p1_addr_reg_5_ );
   nand U25299 ( n25643,n25631,n25647 );
   nand U25300 ( n25647,n25648,n25313,n25649 );
   nand U25301 ( n25649,n25650,n24411,n25298 );
   not U25302 ( n24411,p1_reg2_reg_5_ );
   nand U25303 ( n25648,n25651,n25652,n25283 );
   not U25304 ( n25652,p1_reg1_reg_5_ );
   nand U25305 ( n25642,n25653,n25651,n25283 );
   nand U25306 ( n25651,n25654,n25655,n25656 );
   xor U25307 ( n25656,p1_reg1_reg_5_,n25631 );
   nand U25308 ( n25654,n25657,n25658 );
   nand U25309 ( n25653,n25629,n25659 );
   nand U25310 ( n25659,n25630,p1_reg1_reg_5_ );
   not U25311 ( n25629,n25632 );
   nand U25312 ( n25632,n25658,n25660 );
   nand U25313 ( n25660,n25661,n25655 );
   nand U25314 ( n25641,n25662,n25650,n25298 );
   nand U25315 ( n25650,n25663,n25664,n25665 );
   xor U25316 ( n25665,p1_reg2_reg_5_,n25631 );
   nand U25317 ( n25663,n25666,n25667 );
   nand U25318 ( n25662,n25639,n25668 );
   nand U25319 ( n25668,n25630,p1_reg2_reg_5_ );
   not U25320 ( n25639,n25640 );
   nand U25321 ( n25640,n25667,n25669 );
   nand U25322 ( n25669,n25670,n25664 );
   nand U25323 ( p1_u3247,n25671,n25672,n25673,n25674 );
   nor U25324 ( n25674,n25675,n25676,n25677 );
   nor U25325 ( n25677,n25567,n25678,n25679 );
   nor U25326 ( n25679,n25680,n25661 );
   and U25327 ( n25680,n25655,n25658 );
   nand U25328 ( n25658,n25681,p1_reg1_reg_4_ );
   not U25329 ( n25655,n25682 );
   nor U25330 ( n25678,n25682,n25657 );
   not U25331 ( n25657,n25661 );
   nor U25332 ( n25682,n25681,p1_reg1_reg_4_ );
   not U25333 ( n25676,n25683 );
   nor U25334 ( n25675,n25684,n25685,n25686 );
   nor U25335 ( n25686,n25687,n25670 );
   and U25336 ( n25687,n25664,n25667 );
   nand U25337 ( n25667,n25681,p1_reg2_reg_4_ );
   not U25338 ( n25664,n25688 );
   nor U25339 ( n25685,n25688,n25666 );
   not U25340 ( n25666,n25670 );
   nor U25341 ( n25688,n25681,p1_reg2_reg_4_ );
   nand U25342 ( n25673,p1_reg3_reg_4_,p1_u3086 );
   nand U25343 ( n25672,n25681,n25689 );
   nand U25344 ( n25689,n25690,n25313,n25691 );
   nand U25345 ( n25691,p1_reg1_reg_4_,n25661,n25283 );
   nand U25346 ( n25661,n25692,n25693 );
   nand U25347 ( n25693,p1_reg1_reg_3_,n25694 );
   or U25348 ( n25694,n25695,n25696 );
   nand U25349 ( n25692,n25696,n25695 );
   nand U25350 ( n25690,p1_reg2_reg_4_,n25670,n25298 );
   nand U25351 ( n25670,n25697,n25698 );
   nand U25352 ( n25698,p1_reg2_reg_3_,n25699 );
   or U25353 ( n25699,n25700,n25696 );
   nand U25354 ( n25697,n25696,n25700 );
   nand U25355 ( n25671,n25337,p1_addr_reg_4_ );
   nand U25356 ( p1_u3246,n25701,n25702,n25703,n25704 );
   nor U25357 ( n25704,n25705,n25706 );
   nor U25358 ( n25705,n15179,n25279 );
   not U25359 ( n15179,p1_addr_reg_3_ );
   nand U25360 ( n25703,n25280,n25696 );
   nand U25361 ( n25702,n25283,n25707 );
   xor U25362 ( n25707,n25708,n25696 );
   xor U25363 ( n25708,n25695,p1_reg1_reg_3_ );
   nand U25364 ( n25695,n25709,n25710 );
   nand U25365 ( n25710,n25711,n25712 );
   nand U25366 ( n25701,n25298,n25713 );
   xor U25367 ( n25713,n25714,n25715 );
   xor U25368 ( n25714,n25700,n24354 );
   not U25369 ( n24354,p1_reg2_reg_3_ );
   nand U25370 ( n25700,n25716,n25717 );
   nand U25371 ( n25717,n25718,n25719 );
   nand U25372 ( p1_u3245,n25720,n25683,n25721,n25722 );
   nor U25373 ( n25722,n25723,n25724,n25725 );
   and U25374 ( n25725,p1_addr_reg_2_,n25337 );
   nor U25375 ( n25724,n25726,n25313 );
   nor U25376 ( n25723,p1_state_reg,n25727 );
   nand U25377 ( n25721,n25728,n25729,n25298 );
   nand U25378 ( n25729,n25716,n25719,n25718 );
   nand U25379 ( n25719,n25726,n24331 );
   not U25380 ( n24331,p1_reg2_reg_2_ );
   nand U25381 ( n25716,n25730,p1_reg2_reg_2_ );
   nand U25382 ( n25728,n25731,n25732 );
   not U25383 ( n25732,n25718 );
   nand U25384 ( n25718,n25733,n25734 );
   nand U25385 ( n25734,n25735,n25736 );
   not U25386 ( n25735,n25737 );
   xor U25387 ( n25731,p1_reg2_reg_2_,n25726 );
   nand U25388 ( n25683,n25738,n25739,p1_u4016 );
   nand U25389 ( n25739,n25740,n25741,n25106 );
   nand U25390 ( n25741,n25742,n25737 );
   nand U25391 ( n25740,n25743,n25744 );
   nand U25392 ( n25738,n25745,n25746 );
   nand U25393 ( n25745,n25106,n25747 );
   nand U25394 ( n25747,n25742,n24279 );
   nand U25395 ( n25720,n25748,n25749,n25283 );
   nand U25396 ( n25749,n25709,n25712,n25711 );
   or U25397 ( n25712,n25730,p1_reg1_reg_2_ );
   nand U25398 ( n25709,n25730,p1_reg1_reg_2_ );
   nand U25399 ( n25748,n25750,n25751 );
   not U25400 ( n25751,n25711 );
   nand U25401 ( n25711,n25752,n25753 );
   nand U25402 ( n25753,p1_reg1_reg_0_,n25754,p1_ir_reg_0_ );
   xor U25403 ( n25750,p1_reg1_reg_2_,n25726 );
   nand U25404 ( p1_u3244,n25755,n25756,n25757,n25758 );
   nor U25405 ( n25758,n25759,n25760 );
   nor U25406 ( n25760,p1_state_reg,n24301 );
   nor U25407 ( n25759,n15188,n25279 );
   not U25408 ( n15188,p1_addr_reg_1_ );
   nand U25409 ( n25757,n25280,n25761 );
   not U25410 ( n25280,n25313 );
   nand U25411 ( n25756,n25298,n25762 );
   xor U25412 ( n25762,n25763,n25737 );
   nand U25413 ( n25737,p1_ir_reg_0_,p1_reg2_reg_0_ );
   nand U25414 ( n25763,n25733,n25736 );
   or U25415 ( n25736,n25761,p1_reg2_reg_1_ );
   nand U25416 ( n25733,n25761,p1_reg2_reg_1_ );
   nand U25417 ( n25755,n25283,n25764 );
   xor U25418 ( n25764,n25765,n25766 );
   nand U25419 ( n25766,n25752,n25754 );
   or U25420 ( n25754,n25761,p1_reg1_reg_1_ );
   nand U25421 ( n25752,n25761,p1_reg1_reg_1_ );
   nand U25422 ( n25765,p1_ir_reg_0_,p1_reg1_reg_0_ );
   nand U25423 ( p1_u3243,n25767,n25768,n25769,n25770 );
   nand U25424 ( n25770,p1_ir_reg_0_,n25771 );
   nand U25425 ( n25771,n25772,n25313,n25773 );
   nand U25426 ( n25773,n25298,n24279 );
   not U25427 ( n24279,p1_reg2_reg_0_ );
   nand U25428 ( n25313,n25774,n25264 );
   or U25429 ( n25772,n25567,p1_reg1_reg_0_ );
   nand U25430 ( n25769,n25775,n25746 );
   nand U25431 ( n25775,n25776,n25777 );
   nand U25432 ( n25777,n25283,p1_reg1_reg_0_ );
   nand U25433 ( n25567,n25774,n25743 );
   nand U25434 ( n25776,n25298,p1_reg2_reg_0_ );
   nand U25435 ( n25684,n25742,n25106,n25774 );
   and U25436 ( n25774,n25778,n25279 );
   nand U25437 ( n25778,n25779,n25780 );
   nand U25438 ( n25780,n23566,n25781 );
   nand U25439 ( n25781,n25782,n25783,n23748,n25784 );
   nor U25440 ( n25784,n25012,n25112,n25785,n25266 );
   not U25441 ( n25112,n25269 );
   not U25442 ( n23748,n23652 );
   nand U25443 ( n23652,n25786,n24347 );
   not U25444 ( n25786,n24712 );
   nand U25445 ( n24712,n24346,n24400 );
   nor U25446 ( n24346,n24474,n24672 );
   not U25447 ( n24672,n24397 );
   nand U25448 ( n24397,n23979,n25787,n23989 );
   not U25449 ( n24474,n24403 );
   not U25450 ( n25782,n25267 );
   not U25451 ( n25742,n25743 );
   nand U25452 ( n25768,n25337,p1_addr_reg_0_ );
   not U25453 ( n25337,n25279 );
   nand U25454 ( n25279,n25788,n25789 );
   nand U25455 ( n25788,n25790,n25791 );
   nand U25456 ( n25767,p1_reg3_reg_0_,p1_u3086 );
   nand U25457 ( p1_u3242,n25792,n25793 );
   nand U25458 ( n25793,n25794,n25795 );
   nand U25459 ( n25795,n25796,n25797,n25798,n25799 );
   nand U25460 ( n25799,n23989,n25800,n25801 );
   nand U25461 ( n25800,n25802,n23985 );
   nand U25462 ( n25798,n25803,n25804 );
   or U25463 ( n25803,n25805,n23575 );
   nand U25464 ( n23742,n23978,n23990 );
   or U25465 ( n25797,n25806,n25807,n25808 );
   nand U25466 ( n25796,n25809,n25810 );
   nand U25467 ( n25810,n25811,n25812,n25813 );
   nand U25468 ( n25813,n25814,n25808 );
   nand U25469 ( n25808,n25815,n25816,n25817,n25818 );
   nor U25470 ( n25818,n25819,n25820,n25821,n25822 );
   nand U25471 ( n25822,n24623,n24647,n24674,n24809 );
   nand U25472 ( n24809,n25144,n25141 );
   nand U25473 ( n25141,n24804,n23414 );
   nand U25474 ( n25144,n23741,n23759 );
   nand U25475 ( n24674,n25154,n25184 );
   nand U25476 ( n25184,n23426,n24676 );
   nand U25477 ( n25154,n23796,n23810 );
   nand U25478 ( n24647,n24680,n24681 );
   nand U25479 ( n24681,n24670,n24639 );
   not U25480 ( n24639,n23822 );
   not U25481 ( n24670,n23429 );
   nand U25482 ( n24680,n23429,n23822 );
   or U25483 ( n24623,n24686,n25823 );
   nor U25484 ( n25823,n23432,n24628 );
   nor U25485 ( n24686,n23835,n23820 );
   nand U25486 ( n25821,n24826,n24848,n24874,n24919 );
   nand U25487 ( n24919,n25132,n25134 );
   nand U25488 ( n25134,n23692,n23707 );
   not U25489 ( n23707,n24917 );
   nand U25490 ( n25132,n23402,n24917 );
   nand U25491 ( n24874,n24881,n25139 );
   nand U25492 ( n25139,n23728,n23719 );
   nand U25493 ( n24881,n24876,n23405 );
   nand U25494 ( n24848,n24883,n24886 );
   nand U25495 ( n24886,n23744,n24842 );
   not U25496 ( n24842,n23729 );
   nand U25497 ( n24883,n23729,n23408 );
   not U25498 ( n24826,n24828 );
   nor U25499 ( n24828,n24922,n25824 );
   nor U25500 ( n25824,n23411,n23745 );
   nor U25501 ( n24922,n25185,n24822 );
   not U25502 ( n24822,n23745 );
   not U25503 ( n25185,n23411 );
   nand U25504 ( n25820,n24993,n25010,n25040,n25079 );
   nand U25505 ( n25079,n25120,n25122 );
   not U25506 ( n25122,n25123 );
   nor U25507 ( n25123,n23384,n25089 );
   nand U25508 ( n25120,n23384,n25089 );
   nand U25509 ( n25040,n25094,n25093 );
   nand U25510 ( n25093,n25047,n23387 );
   nand U25511 ( n25094,n23650,n23638 );
   not U25512 ( n23638,n25047 );
   nand U25513 ( n25010,n25052,n25054 );
   nand U25514 ( n25054,n23667,n23649 );
   not U25515 ( n23649,n25194 );
   nand U25516 ( n25052,n25194,n23390 );
   nand U25517 ( n24993,n25056,n25058 );
   nand U25518 ( n25058,n24994,n23393 );
   nand U25519 ( n25056,n23648,n23666 );
   not U25520 ( n23666,n24994 );
   nand U25521 ( n25819,n25118,n24772,n25825,n24540 );
   nand U25522 ( n24540,n24583,n24586 );
   nand U25523 ( n24586,n25230,n23858 );
   not U25524 ( n23858,n25231 );
   not U25525 ( n25230,n23438 );
   nand U25526 ( n24583,n23438,n25231 );
   not U25527 ( n25825,n23977 );
   nor U25528 ( n23977,n25826,n24293 );
   nor U25529 ( n24293,n24278,n23960 );
   not U25530 ( n23960,n23465 );
   not U25531 ( n24278,n23974 );
   nor U25532 ( n25826,n23465,n23974 );
   nand U25533 ( n24772,n24811,n24808 );
   nand U25534 ( n24808,n23766,n23417 );
   nand U25535 ( n24811,n23783,n24745 );
   not U25536 ( n24745,n23766 );
   nand U25537 ( n25118,n25827,n24019 );
   nand U25538 ( n24019,n25828,n24035 );
   not U25539 ( n25827,n24021 );
   nor U25540 ( n24021,n25828,n24035 );
   not U25541 ( n24035,n23609 );
   not U25542 ( n25828,n23381 );
   nor U25543 ( n25817,n25829,n25830 );
   or U25544 ( n25830,n25831,n25832,n24352,n24409 );
   xor U25545 ( n24409,n23450,n24412 );
   not U25546 ( n24352,n24351 );
   xor U25547 ( n24351,n23918,n23934 );
   xor U25548 ( n25832,n23574,n23372 );
   xor U25549 ( n25831,n23375,n23582 );
   or U25550 ( n25829,n24479,n24700,n24725,n24932 );
   xor U25551 ( n24932,n24963,n23693 );
   not U25552 ( n23693,n24934 );
   not U25553 ( n24963,n23399 );
   xor U25554 ( n24725,n23420,n24726 );
   xor U25555 ( n24700,n23423,n23799 );
   not U25556 ( n24479,n24487 );
   xor U25557 ( n24487,n24516,n24482 );
   nor U25558 ( n25816,n24575,n24521,n24441,n24370 );
   nor U25559 ( n24370,n24416,n24415 );
   not U25560 ( n24415,n25170 );
   nand U25561 ( n25170,n23933,n23919 );
   nor U25562 ( n24416,n23919,n23933 );
   and U25563 ( n24441,n24489,n24486 );
   nand U25564 ( n24486,n24446,n23447 );
   nand U25565 ( n24489,n24471,n23897 );
   not U25566 ( n24521,n24510 );
   nand U25567 ( n24510,n25161,n25162 );
   nand U25568 ( n25162,n23857,n23874 );
   not U25569 ( n23874,n24525 );
   nand U25570 ( n25161,n24525,n23441 );
   not U25571 ( n24575,n24584 );
   nand U25572 ( n24584,n25159,n25156 );
   nand U25573 ( n25156,n24578,n23435 );
   nand U25574 ( n25159,n23859,n23847 );
   not U25575 ( n23847,n24578 );
   nor U25576 ( n25815,n24314,n24294,n24030,n24978 );
   not U25577 ( n24978,n24975 );
   xor U25578 ( n24975,n23665,n24979 );
   not U25579 ( n24030,n24017 );
   xor U25580 ( n24017,n23605,n23594 );
   not U25581 ( n23605,n23378 );
   nor U25582 ( n24294,n24320,n25833 );
   nor U25583 ( n25833,n23462,n24296 );
   nor U25584 ( n24320,n23946,n23961 );
   not U25585 ( n23961,n24296 );
   not U25586 ( n23946,n23462 );
   and U25587 ( n24314,n24359,n25179 );
   nand U25588 ( n25179,n24321,n23459 );
   nand U25589 ( n24359,n23962,n23947 );
   nand U25590 ( n25812,n25105,n25804 );
   nand U25591 ( n25811,n25806,n23987,n25801 );
   not U25592 ( n25801,n25804 );
   nand U25593 ( n25804,n25834,n25835,n25836,n25837 );
   nand U25594 ( n25837,n25838,n25839,n25840,n25841 );
   nand U25595 ( n25841,n25842,n25843,n25844 );
   not U25596 ( n25844,n25845 );
   nand U25597 ( n25840,n25846,n25847 );
   nand U25598 ( n25847,n25845,n25848 );
   nand U25599 ( n25848,n25842,n25843 );
   nand U25600 ( n25843,n25849,n25850 );
   nand U25601 ( n25842,n25851,n25852,n25853 );
   or U25602 ( n25853,n25850,n25849 );
   and U25603 ( n25849,n25854,n25855 );
   nand U25604 ( n25855,n25856,n23384 );
   nand U25605 ( n25854,n25857,n25089 );
   nand U25606 ( n25850,n25858,n25859 );
   nand U25607 ( n25859,n25860,n23384 );
   nand U25608 ( n25858,n25861,n25089 );
   nand U25609 ( n25852,n25862,n25863,n25864 );
   nand U25610 ( n25864,n25865,n25866 );
   nand U25611 ( n25863,n25867,n25868,n25869 );
   nand U25612 ( n25869,n25870,n25871 );
   nand U25613 ( n25868,n25872,n25873,n25874 );
   nand U25614 ( n25874,n25875,n25876 );
   nand U25615 ( n25873,n25877,n25878,n25879 );
   nand U25616 ( n25879,n25880,n25881 );
   nand U25617 ( n25878,n25882,n25883,n25884 );
   nand U25618 ( n25884,n25885,n25886 );
   nand U25619 ( n25883,n25887,n25888,n25889 );
   nand U25620 ( n25889,n25890,n25891 );
   nand U25621 ( n25888,n25892,n25893,n25894 );
   nand U25622 ( n25894,n25895,n25896 );
   nand U25623 ( n25893,n25897,n25898,n25899 );
   nand U25624 ( n25899,n25900,n25901 );
   nand U25625 ( n25898,n25902,n25903,n25904 );
   nand U25626 ( n25904,n25905,n25906 );
   nand U25627 ( n25903,n25907,n25908,n25909 );
   nand U25628 ( n25909,n25910,n25911 );
   nand U25629 ( n25908,n25912,n25913,n25914 );
   nand U25630 ( n25914,n25915,n25916 );
   nand U25631 ( n25913,n25917,n25918,n25919 );
   nand U25632 ( n25919,n25920,n25921 );
   nand U25633 ( n25918,n25922,n25923,n25924 );
   nand U25634 ( n25924,n25925,n25926 );
   nand U25635 ( n25923,n25927,n25928,n25929 );
   nand U25636 ( n25929,n25930,n25931 );
   nand U25637 ( n25928,n25932,n25933,n25934 );
   nand U25638 ( n25934,n25935,n25936 );
   nand U25639 ( n25933,n25937,n25938,n25939 );
   nand U25640 ( n25939,n25940,n25941 );
   nand U25641 ( n25938,n25942,n25943,n25944 );
   or U25642 ( n25944,n25941,n25940 );
   and U25643 ( n25940,n25945,n25946 );
   nand U25644 ( n25946,n25860,n23435 );
   nand U25645 ( n25945,n25861,n24578 );
   nand U25646 ( n25941,n25947,n25948 );
   nand U25647 ( n25948,n25856,n23435 );
   nand U25648 ( n25947,n25857,n24578 );
   nand U25649 ( n25943,n25949,n25950,n25951 );
   not U25650 ( n25951,n25952 );
   nand U25651 ( n25942,n25953,n25954 );
   nand U25652 ( n25954,n25952,n25955 );
   nand U25653 ( n25955,n25949,n25950 );
   nand U25654 ( n25950,n25956,n25957,n25958 );
   nand U25655 ( n25958,n25959,n25960 );
   nand U25656 ( n25957,n25961,n25962,n25963 );
   not U25657 ( n25963,n25964 );
   nand U25658 ( n25956,n25965,n25966 );
   nand U25659 ( n25966,n25964,n25967 );
   nand U25660 ( n25967,n25961,n25962 );
   nand U25661 ( n25962,n25968,n25969,n25970 );
   nand U25662 ( n25970,n25971,n25972 );
   nand U25663 ( n25969,n25973,n25974,n25975 );
   not U25664 ( n25975,n25976 );
   nand U25665 ( n25968,n25977,n25978 );
   nand U25666 ( n25978,n25976,n25979 );
   nand U25667 ( n25979,n25973,n25974 );
   nand U25668 ( n25974,n25980,n25981,n25982 );
   nand U25669 ( n25982,n25983,n25984 );
   nand U25670 ( n25981,n25985,n25986,n25987 );
   not U25671 ( n25987,n25988 );
   nand U25672 ( n25980,n25989,n25990 );
   nand U25673 ( n25990,n25988,n25991 );
   nand U25674 ( n25991,n25985,n25986 );
   nand U25675 ( n25986,n25992,n25993,n25994 );
   nand U25676 ( n25994,n25995,n25996 );
   nand U25677 ( n25993,n25997,n25998,n25999 );
   not U25678 ( n25999,n26000 );
   nand U25679 ( n25992,n26001,n26002 );
   nand U25680 ( n26002,n26000,n26003 );
   nand U25681 ( n26003,n25997,n25998 );
   nand U25682 ( n25998,n26004,n26005 );
   nand U25683 ( n26005,n26006,n26007 );
   nand U25684 ( n26007,n23974,n25857 );
   nand U25685 ( n26006,n23465,n25856 );
   nand U25686 ( n26004,n26008,n26009 );
   or U25687 ( n25997,n26009,n26008 );
   or U25688 ( n26008,n25857,n26010 );
   nor U25689 ( n26010,n25809,n23990 );
   nand U25690 ( n26009,n26011,n26012 );
   nand U25691 ( n26012,n25860,n23465 );
   nand U25692 ( n26011,n25861,n23974 );
   nand U25693 ( n26000,n26013,n26014 );
   nand U25694 ( n26014,n25856,n23462 );
   nand U25695 ( n26013,n25857,n24296 );
   nand U25696 ( n26001,n26015,n26016 );
   nand U25697 ( n26016,n25860,n23462 );
   nand U25698 ( n26015,n25861,n24296 );
   or U25699 ( n25985,n25996,n25995 );
   and U25700 ( n25995,n26017,n26018 );
   nand U25701 ( n26018,n25856,n23459 );
   nand U25702 ( n26017,n25857,n24321 );
   nand U25703 ( n25996,n26019,n26020 );
   nand U25704 ( n26020,n25860,n23459 );
   nand U25705 ( n26019,n25861,n24321 );
   nand U25706 ( n25988,n26021,n26022 );
   nand U25707 ( n26022,n25856,n23456 );
   nand U25708 ( n26021,n25857,n23934 );
   nand U25709 ( n25989,n26023,n26024 );
   nand U25710 ( n26024,n25860,n23456 );
   nand U25711 ( n26023,n25861,n23934 );
   or U25712 ( n25973,n25984,n25983 );
   and U25713 ( n25983,n26025,n26026 );
   nand U25714 ( n26026,n25856,n23453 );
   nand U25715 ( n26025,n25857,n24372 );
   nand U25716 ( n25984,n26027,n26028 );
   nand U25717 ( n26028,n25860,n23453 );
   nand U25718 ( n26027,n25861,n24372 );
   nand U25719 ( n25976,n26029,n26030 );
   nand U25720 ( n26030,n25856,n23450 );
   nand U25721 ( n26029,n25857,n24412 );
   nand U25722 ( n25977,n26031,n26032 );
   nand U25723 ( n26032,n25860,n23450 );
   nand U25724 ( n26031,n25861,n24412 );
   or U25725 ( n25961,n25972,n25971 );
   and U25726 ( n25971,n26033,n26034 );
   nand U25727 ( n26034,n25856,n23447 );
   nand U25728 ( n26033,n25857,n24446 );
   nand U25729 ( n25972,n26035,n26036 );
   nand U25730 ( n26036,n25860,n23447 );
   nand U25731 ( n26035,n25861,n24446 );
   nand U25732 ( n25964,n26037,n26038 );
   nand U25733 ( n26038,n25856,n23444 );
   nand U25734 ( n26037,n25857,n24482 );
   nand U25735 ( n25965,n26039,n26040 );
   nand U25736 ( n26040,n25860,n23444 );
   nand U25737 ( n26039,n25861,n24482 );
   or U25738 ( n25949,n25960,n25959 );
   and U25739 ( n25959,n26041,n26042 );
   nand U25740 ( n26042,n25856,n23441 );
   nand U25741 ( n26041,n25857,n24525 );
   nand U25742 ( n25960,n26043,n26044 );
   nand U25743 ( n26044,n25860,n23441 );
   nand U25744 ( n26043,n25861,n24525 );
   nand U25745 ( n25952,n26045,n26046 );
   nand U25746 ( n26046,n25856,n23438 );
   nand U25747 ( n26045,n25857,n25231 );
   nand U25748 ( n25953,n26047,n26048 );
   nand U25749 ( n26048,n25860,n23438 );
   nand U25750 ( n26047,n25861,n25231 );
   or U25751 ( n25937,n25936,n25935 );
   and U25752 ( n25935,n26049,n26050 );
   nand U25753 ( n26050,n25856,n23432 );
   nand U25754 ( n26049,n25857,n24628 );
   nand U25755 ( n25936,n26051,n26052 );
   nand U25756 ( n26052,n25860,n23432 );
   nand U25757 ( n26051,n25861,n24628 );
   or U25758 ( n25932,n25931,n25930 );
   and U25759 ( n25930,n26053,n26054 );
   nand U25760 ( n26054,n25860,n23429 );
   nand U25761 ( n26053,n25861,n23822 );
   nand U25762 ( n25931,n26055,n26056 );
   nand U25763 ( n26056,n25856,n23429 );
   nand U25764 ( n26055,n25857,n23822 );
   or U25765 ( n25927,n25926,n25925 );
   and U25766 ( n25925,n26057,n26058 );
   nand U25767 ( n26058,n25856,n23426 );
   nand U25768 ( n26057,n25857,n24676 );
   nand U25769 ( n25926,n26059,n26060 );
   nand U25770 ( n26060,n25860,n23426 );
   nand U25771 ( n26059,n25861,n24676 );
   or U25772 ( n25922,n25921,n25920 );
   and U25773 ( n25920,n26061,n26062 );
   nand U25774 ( n26062,n25860,n23423 );
   nand U25775 ( n26061,n25861,n23799 );
   nand U25776 ( n25921,n26063,n26064 );
   nand U25777 ( n26064,n25856,n23423 );
   nand U25778 ( n26063,n25857,n23799 );
   or U25779 ( n25917,n25916,n25915 );
   and U25780 ( n25915,n26065,n26066 );
   nand U25781 ( n26066,n25856,n23420 );
   nand U25782 ( n26065,n25857,n24726 );
   nand U25783 ( n25916,n26067,n26068 );
   nand U25784 ( n26068,n25860,n23420 );
   nand U25785 ( n26067,n25861,n24726 );
   or U25786 ( n25912,n25911,n25910 );
   and U25787 ( n25910,n26069,n26070 );
   nand U25788 ( n26070,n25860,n23417 );
   nand U25789 ( n26069,n25861,n23766 );
   nand U25790 ( n25911,n26071,n26072 );
   nand U25791 ( n26072,n25856,n23417 );
   nand U25792 ( n26071,n25857,n23766 );
   or U25793 ( n25907,n25906,n25905 );
   and U25794 ( n25905,n26073,n26074 );
   nand U25795 ( n26074,n25856,n23414 );
   nand U25796 ( n26073,n25857,n24804 );
   nand U25797 ( n25906,n26075,n26076 );
   nand U25798 ( n26076,n25860,n23414 );
   nand U25799 ( n26075,n25861,n24804 );
   or U25800 ( n25902,n25901,n25900 );
   and U25801 ( n25900,n26077,n26078 );
   nand U25802 ( n26078,n25860,n23411 );
   nand U25803 ( n26077,n25861,n23745 );
   nand U25804 ( n25901,n26079,n26080 );
   nand U25805 ( n26080,n25856,n23411 );
   nand U25806 ( n26079,n25857,n23745 );
   or U25807 ( n25897,n25896,n25895 );
   and U25808 ( n25895,n26081,n26082 );
   nand U25809 ( n26082,n25856,n23408 );
   nand U25810 ( n26081,n25857,n23729 );
   nand U25811 ( n25896,n26083,n26084 );
   nand U25812 ( n26084,n25860,n23408 );
   nand U25813 ( n26083,n25861,n23729 );
   or U25814 ( n25892,n25891,n25890 );
   and U25815 ( n25890,n26085,n26086 );
   nand U25816 ( n26086,n25860,n23405 );
   nand U25817 ( n26085,n25861,n24876 );
   nand U25818 ( n25891,n26087,n26088 );
   nand U25819 ( n26088,n25856,n23405 );
   nand U25820 ( n26087,n25857,n24876 );
   or U25821 ( n25887,n25886,n25885 );
   and U25822 ( n25885,n26089,n26090 );
   nand U25823 ( n26090,n25856,n23402 );
   nand U25824 ( n26089,n25857,n24917 );
   nand U25825 ( n25886,n26091,n26092 );
   nand U25826 ( n26092,n25860,n23402 );
   nand U25827 ( n26091,n25861,n24917 );
   or U25828 ( n25882,n25881,n25880 );
   and U25829 ( n25880,n26093,n26094 );
   nand U25830 ( n26094,n25860,n23399 );
   nand U25831 ( n26093,n25861,n24934 );
   nand U25832 ( n25881,n26095,n26096 );
   nand U25833 ( n26096,n25856,n23399 );
   nand U25834 ( n26095,n25857,n24934 );
   or U25835 ( n25877,n25876,n25875 );
   and U25836 ( n25875,n26097,n26098 );
   nand U25837 ( n26098,n25856,n23396 );
   nand U25838 ( n26097,n25857,n24979 );
   nand U25839 ( n25876,n26099,n26100 );
   nand U25840 ( n26100,n25860,n23396 );
   nand U25841 ( n26099,n25861,n24979 );
   or U25842 ( n25872,n25871,n25870 );
   and U25843 ( n25870,n26101,n26102 );
   nand U25844 ( n26102,n25860,n23393 );
   nand U25845 ( n26101,n25861,n24994 );
   nand U25846 ( n25871,n26103,n26104 );
   nand U25847 ( n26104,n25856,n23393 );
   nand U25848 ( n26103,n25857,n24994 );
   or U25849 ( n25867,n25866,n25865 );
   and U25850 ( n25865,n26105,n26106 );
   nand U25851 ( n26106,n25856,n23390 );
   nand U25852 ( n26105,n25857,n25194 );
   nand U25853 ( n25866,n26107,n26108 );
   nand U25854 ( n26108,n25860,n23390 );
   nand U25855 ( n26107,n25861,n25194 );
   nand U25856 ( n25862,n26109,n26110 );
   or U25857 ( n25851,n26110,n26109 );
   and U25858 ( n26109,n26111,n26112 );
   nand U25859 ( n26112,n25856,n23387 );
   nand U25860 ( n26111,n25857,n25047 );
   nand U25861 ( n26110,n26113,n26114 );
   nand U25862 ( n26114,n25860,n23387 );
   nand U25863 ( n26113,n25861,n25047 );
   nand U25864 ( n25845,n26115,n26116 );
   nand U25865 ( n26116,n25860,n23381 );
   nand U25866 ( n26115,n25861,n23609 );
   nand U25867 ( n25846,n26117,n26118 );
   nand U25868 ( n26118,n25856,n23381 );
   nand U25869 ( n26117,n25857,n23609 );
   or U25870 ( n25839,n26119,n26120 );
   nand U25871 ( n25836,n26121,n26122,n26123 );
   nand U25872 ( n26123,n26124,n23372 );
   nand U25873 ( n25835,n25838,n26119,n26120 );
   and U25874 ( n26120,n26125,n26126 );
   nand U25875 ( n26126,n25856,n23378 );
   nand U25876 ( n26125,n25857,n23594 );
   nand U25877 ( n26119,n26129,n26130 );
   nand U25878 ( n26130,n25860,n23378 );
   nand U25879 ( n26132,n26133,n23987 );
   nand U25880 ( n26129,n25861,n23594 );
   nand U25881 ( n23594,n26134,n26135 );
   nand U25882 ( n26135,n26136,n20860 );
   xor U25883 ( n20860,n26137,n26138 );
   xor U25884 ( n26138,si_29_,n26139 );
   nand U25885 ( n26134,n26140,p2_datao_reg_29_ );
   and U25886 ( n25838,n26141,n26142 );
   or U25887 ( n26142,n26143,n26144 );
   nand U25888 ( n25834,n26143,n26141,n26144 );
   and U25889 ( n26144,n26145,n26146 );
   nand U25890 ( n26146,n25857,n23582 );
   nand U25891 ( n26145,n26147,n23375 );
   nand U25892 ( n26141,n26148,n26149 );
   nand U25893 ( n26149,n26150,n26121 );
   nand U25894 ( n26121,n23574,n25861 );
   not U25895 ( n26148,n26122 );
   nand U25896 ( n26122,n26151,n26152 );
   nand U25897 ( n26152,n25857,n23574 );
   nand U25898 ( n23574,n26153,n26154 );
   nand U25899 ( n26154,n26136,n24253 );
   not U25900 ( n24253,n21927 );
   nand U25901 ( n21927,n26155,n26156 );
   nand U25902 ( n26156,n26157,n26158 );
   nand U25903 ( n26158,n26159,n26160 );
   nand U25904 ( n26160,si_30_,n26161 );
   nand U25905 ( n26155,n26162,n26163 );
   nand U25906 ( n26163,n26161,n26164 );
   nand U25907 ( n26164,n26159,n26165 );
   not U25908 ( n26162,n26157 );
   xor U25909 ( n26157,n26166,si_31_ );
   nor U25910 ( n26166,n26167,n26168 );
   nor U25911 ( n26168,p1_datao_reg_31_,n16576 );
   nor U25912 ( n26167,p2_datao_reg_31_,n16572 );
   nand U25913 ( n26153,n26140,p2_datao_reg_31_ );
   nand U25914 ( n26151,n26147,n23372 );
   not U25915 ( n26147,n26128 );
   nand U25916 ( n26128,n25861,n26169 );
   nand U25917 ( n26169,n25783,n26150,n26170,n26171 );
   nand U25918 ( n26143,n26172,n26173 );
   nand U25919 ( n26173,n26124,n23375 );
   nand U25920 ( n23375,n26174,n26175,n26176 );
   nand U25921 ( n26176,p1_reg2_reg_30_,n26177 );
   nand U25922 ( n26175,p1_reg0_reg_30_,n26178 );
   nand U25923 ( n26174,p1_reg1_reg_30_,n26179 );
   not U25924 ( n26124,n26131 );
   nand U25925 ( n26131,n25857,n26180 );
   nand U25926 ( n26180,n26181,n23975,n26150 );
   not U25927 ( n26150,n23372 );
   nand U25928 ( n23372,n26182,n26183,n26184 );
   nand U25929 ( n26184,p1_reg2_reg_31_,n26177 );
   nand U25930 ( n26183,p1_reg0_reg_31_,n26178 );
   nand U25931 ( n26182,p1_reg1_reg_31_,n26179 );
   nand U25932 ( n23975,n23987,n25814 );
   nand U25933 ( n26181,n25787,n25291 );
   or U25934 ( n26186,n25787,n26187 );
   or U25935 ( n26185,n23985,n23979 );
   nand U25936 ( n23985,n23990,n25787 );
   nand U25937 ( n26172,n25861,n23582 );
   nand U25938 ( n23582,n26189,n26190 );
   nand U25939 ( n26190,n26136,n20869 );
   nand U25940 ( n20869,n26191,n26192 );
   nand U25941 ( n26192,si_30_,n26193 );
   nand U25942 ( n26193,n26161,n26159 );
   or U25943 ( n26159,n26194,n26195 );
   nand U25944 ( n26161,n26195,n26194 );
   nand U25945 ( n26191,n26196,n26165 );
   not U25946 ( n26165,si_30_ );
   xor U25947 ( n26196,n26195,n26194 );
   nand U25948 ( n26194,n26197,n26198 );
   nand U25949 ( n26198,n26199,n26200 );
   not U25950 ( n26200,si_29_ );
   or U25951 ( n26199,n26139,n26137 );
   nand U25952 ( n26197,n26137,n26139 );
   nand U25953 ( n26139,n26201,n26202 );
   nand U25954 ( n26202,n26203,n26204 );
   not U25955 ( n26204,si_28_ );
   or U25956 ( n26203,n26205,n26206 );
   nand U25957 ( n26201,n26206,n26205 );
   nand U25958 ( n26137,n26207,n26208 );
   nand U25959 ( n26208,n16576,n17678 );
   not U25960 ( n17678,p2_datao_reg_29_ );
   nand U25961 ( n26207,n16572,n17679 );
   not U25962 ( n17679,p1_datao_reg_29_ );
   and U25963 ( n26195,n26209,n26210 );
   nand U25964 ( n26210,n16572,p1_datao_reg_30_ );
   nand U25965 ( n26209,n16576,p2_datao_reg_30_ );
   nand U25966 ( n26189,n26140,p2_datao_reg_30_ );
   and U25967 ( n26211,n26170,n25783 );
   nand U25968 ( n25792,n26212,n26213,p1_b_reg );
   or U25969 ( n26213,n25743,n25264,n26214 );
   nand U25970 ( n26212,n25794,n23987 );
   nand U25971 ( p1_u3241,n26215,n26216,n26217,n26218 );
   nor U25972 ( n26218,n26219,n26220,n26221 );
   nor U25973 ( n26221,n23783,n26222 );
   not U25974 ( n23783,n23417 );
   and U25975 ( n26220,n26223,n24736 );
   nor U25976 ( n26219,p1_state_reg,n26224 );
   nand U25977 ( n26217,n26225,n24726 );
   or U25978 ( n26216,n26226,n26227 );
   xor U25979 ( n26226,n26228,n26229 );
   xor U25980 ( n26229,n26230,n26231 );
   nand U25981 ( n26215,n26232,n23423 );
   nand U25982 ( p1_u3240,n26233,n26234,n26235,n26236 );
   nor U25983 ( n26236,n26237,n26238,n26239 );
   nor U25984 ( n26239,n26240,n25024 );
   nor U25985 ( n26238,n23607,n26222 );
   nor U25986 ( n26237,p1_state_reg,n26241 );
   nand U25987 ( n26235,n26232,n23390 );
   nand U25988 ( n26234,n26242,n26243,n26244 );
   nand U25989 ( n26243,n26245,n26246,n26247 );
   nand U25990 ( n26247,n26248,n26249 );
   nand U25991 ( n26245,n26250,n26251 );
   nand U25992 ( n26242,n26252,n26248,n26253 );
   nand U25993 ( n26252,n26254,n26246 );
   nand U25994 ( n26233,n26225,n25047 );
   nand U25995 ( p1_u3239,n26255,n26256,n26257,n26258 );
   nor U25996 ( n26258,n25617,n26259,n26260 );
   nor U25997 ( n26260,n23920,n26261 );
   nor U25998 ( n26259,n24516,n26222 );
   nor U25999 ( n25617,p1_state_reg,n26262 );
   nand U26000 ( n26257,n26263,n26223 );
   or U26001 ( n26256,n26264,n26227 );
   xor U26002 ( n26264,n26265,n26266 );
   xor U26003 ( n26265,n26267,n26268 );
   nand U26004 ( n26255,n26225,n24446 );
   nand U26005 ( p1_u3238,n26269,n26270,n26271,n26272 );
   nor U26006 ( n26272,n26273,n26274,n26275 );
   nor U26007 ( n26275,n23744,n26222 );
   not U26008 ( n23744,n23408 );
   nor U26009 ( n26274,n23741,n26261 );
   nor U26010 ( n26273,p1_state_reg,n26276 );
   nand U26011 ( n26271,n26277,n26223 );
   or U26012 ( n26270,n26278,n26227 );
   xor U26013 ( n26278,n26279,n26280 );
   xor U26014 ( n26279,n26281,n26282 );
   nand U26015 ( n26269,n26225,n23745 );
   nand U26016 ( p1_u3237,n26283,n26284,n26285 );
   nor U26017 ( n26285,n26286,n26287,n26288 );
   nor U26018 ( n26288,n26289,n25727 );
   not U26019 ( n25727,p1_reg3_reg_2_ );
   nor U26020 ( n26287,n26227,n26290,n26291 );
   and U26021 ( n26291,n26292,n26293,n26294 );
   nor U26022 ( n26290,n26292,n26295 );
   xor U26023 ( n26295,n26296,n26297 );
   nor U26024 ( n26286,n23947,n26298 );
   not U26025 ( n23947,n24321 );
   nand U26026 ( n26284,n26299,n23456 );
   nand U26027 ( n26283,n26232,n23462 );
   nand U26028 ( p1_u3236,n26300,n26301,n26302,n26303 );
   nor U26029 ( n26303,n26304,n26305,n26306 );
   nor U26030 ( n26306,n26240,n24596 );
   not U26031 ( n24596,n26307 );
   nor U26032 ( n26305,n23835,n26298 );
   not U26033 ( n23835,n24628 );
   and U26034 ( n26304,p1_u3086,p1_reg3_reg_11_ );
   nand U26035 ( n26302,n26299,n23429 );
   nand U26036 ( n26301,n26308,n26244 );
   xor U26037 ( n26308,n26309,n26310 );
   xor U26038 ( n26310,n26311,n26312 );
   nand U26039 ( n26300,n26232,n23435 );
   nand U26040 ( p1_u3235,n26313,n26314,n26315,n26316 );
   nor U26041 ( n26316,n26317,n26318,n26319 );
   nor U26042 ( n26319,n23665,n26222 );
   not U26043 ( n23665,n23396 );
   nor U26044 ( n26318,n23692,n26261 );
   not U26045 ( n23692,n23402 );
   nor U26046 ( n26317,p1_state_reg,n26320 );
   nand U26047 ( n26315,n24945,n26223 );
   or U26048 ( n26314,n26227,n26321 );
   xor U26049 ( n26321,n26322,n26323 );
   xor U26050 ( n26323,n26324,n26325 );
   nand U26051 ( n26313,n26225,n24934 );
   nand U26052 ( p1_u3234,n26326,n26327,n26328,n26329 );
   nor U26053 ( n26329,n25446,n26330,n26331 );
   nor U26054 ( n26331,n26240,n24658 );
   nor U26055 ( n26330,n23810,n26298 );
   not U26056 ( n23810,n24676 );
   nor U26057 ( n25446,p1_state_reg,n26332 );
   nand U26058 ( n26328,n26232,n23429 );
   nand U26059 ( n26327,n26333,n26334,n26244 );
   nand U26060 ( n26334,n26335,n26336 );
   nand U26061 ( n26336,n26337,n26338 );
   nand U26062 ( n26333,n26337,n26338,n26339 );
   nand U26063 ( n26326,n26299,n23423 );
   nand U26064 ( p1_u3233,n26340,n26341,n26342,n26343 );
   nor U26065 ( n26343,n26344,n26345,n26346 );
   nor U26066 ( n26346,n26240,n24861 );
   not U26067 ( n24861,n26347 );
   nor U26068 ( n26345,n23719,n26298 );
   not U26069 ( n23719,n24876 );
   nor U26070 ( n26344,p1_state_reg,n26348 );
   nand U26071 ( n26342,n26232,n23408 );
   nand U26072 ( n26341,n26349,n26350,n26244 );
   or U26073 ( n26350,n26351,n26352 );
   xor U26074 ( n26351,n26353,n26354 );
   nand U26075 ( n26349,n26355,n26356,n26352 );
   nand U26076 ( n26340,n26299,n23402 );
   nand U26077 ( p1_u3232,n26357,n26358,n26359,n26360 );
   nand U26078 ( n26360,p1_reg3_reg_0_,n26361 );
   nand U26079 ( n26359,n26244,n25744 );
   xor U26080 ( n25744,n26362,n26363 );
   xor U26081 ( n26363,n26364,n26365 );
   nand U26082 ( n26358,n26225,n23974 );
   nand U26083 ( n26357,n26299,n23462 );
   nand U26084 ( p1_u3231,n26366,n26367,n26368,n26369 );
   nor U26085 ( n26369,n25538,n26370,n26371 );
   nor U26086 ( n26371,n23857,n26261 );
   nor U26087 ( n26370,n23859,n26222 );
   not U26088 ( n23859,n23435 );
   nor U26089 ( n25538,p1_state_reg,n26372 );
   nand U26090 ( n26368,n24537,n26223 );
   or U26091 ( n26367,n26373,n26227 );
   xor U26092 ( n26373,n26374,n26375 );
   xor U26093 ( n26375,n26376,n26377 );
   nand U26094 ( n26366,n26225,n25231 );
   nand U26095 ( p1_u3230,n26378,n26379,n26380,n26381 );
   nor U26096 ( n26381,n26382,n26383,n26384 );
   nor U26097 ( n26384,n23918,n26261 );
   not U26098 ( n23918,n23456 );
   nor U26099 ( n26383,n23920,n26222 );
   not U26100 ( n23920,n23450 );
   nor U26101 ( n26382,p1_state_reg,n26385 );
   nand U26102 ( n26380,n26225,n24372 );
   nand U26103 ( n26379,n26386,n26223 );
   or U26104 ( n26378,n26387,n26227 );
   xor U26105 ( n26387,n26388,n26389 );
   xor U26106 ( n26388,n26390,n26391 );
   nand U26107 ( p1_u3229,n26392,n26393,n26394,n26395 );
   nor U26108 ( n26395,n26396,n26397,n26398 );
   nor U26109 ( n26398,n23667,n26222 );
   not U26110 ( n23667,n23390 );
   nor U26111 ( n26397,n26240,n24989 );
   nor U26112 ( n26396,p1_state_reg,n26399 );
   nand U26113 ( n26394,n26225,n24994 );
   nand U26114 ( n26393,n26244,n26400 );
   xor U26115 ( n26400,n26401,n26402 );
   nand U26116 ( n26401,n26403,n26404 );
   nand U26117 ( n26392,n26232,n23396 );
   nand U26118 ( p1_u3228,n26405,n26406,n26407,n26408 );
   nor U26119 ( n26408,n25343,n26409,n26410 );
   nor U26120 ( n26410,n26240,n24788 );
   nor U26121 ( n26409,n23759,n26298 );
   not U26122 ( n23759,n24804 );
   nor U26123 ( n25343,p1_state_reg,n26411 );
   not U26124 ( n26411,p1_reg3_reg_17_ );
   nand U26125 ( n26407,n26232,n23417 );
   nand U26126 ( n26406,n26412,n26413,n26244 );
   nand U26127 ( n26413,n26414,n26415 );
   nand U26128 ( n26415,n26416,n26417 );
   nand U26129 ( n26412,n26416,n26417,n26418 );
   nand U26130 ( n26405,n26299,n23411 );
   nand U26131 ( p1_u3227,n26419,n26420,n26421,n26422 );
   nor U26132 ( n26422,n25646,n26423,n26424 );
   nor U26133 ( n26424,n23933,n26261 );
   nor U26134 ( n26423,n24471,n26222 );
   nor U26135 ( n25646,p1_state_reg,n26425 );
   nand U26136 ( n26421,n24385,n26223 );
   nand U26137 ( n26420,n26426,n26244 );
   xor U26138 ( n26426,n26427,n26428 );
   xor U26139 ( n26427,n26429,n26430 );
   nand U26140 ( n26419,n26225,n24412 );
   nand U26141 ( p1_u3226,n26431,n26432,n26433,n26434 );
   nor U26142 ( n26434,n26435,n26436,n26437 );
   nor U26143 ( n26437,n23741,n26222 );
   not U26144 ( n23741,n23414 );
   nor U26145 ( n26436,n26240,n24746 );
   nor U26146 ( n26435,p1_state_reg,n26438 );
   nand U26147 ( n26433,n26225,n23766 );
   nand U26148 ( n26432,n26439,n26244 );
   xor U26149 ( n26439,n26440,n26441 );
   xor U26150 ( n26441,n26442,n26443 );
   nand U26151 ( n26431,n26232,n23420 );
   nand U26152 ( p1_u3225,n26444,n26445,n26446,n26447 );
   nor U26153 ( n26447,n26448,n26449,n26450 );
   nor U26154 ( n26450,n23650,n26222 );
   nor U26155 ( n26449,n26240,n25006 );
   and U26156 ( n26448,p1_u3086,p1_reg3_reg_25_ );
   nand U26157 ( n26446,n26225,n25194 );
   nand U26158 ( n26445,n26244,n26451 );
   nand U26159 ( n26451,n26452,n26453,n26454 );
   or U26160 ( n26454,n26246,n26254 );
   nand U26161 ( n26453,n26254,n26455,n26456 );
   nand U26162 ( n26452,n26457,n26458 );
   xor U26163 ( n26457,n26254,n26455 );
   not U26164 ( n26254,n26251 );
   nand U26165 ( n26251,n26403,n26459 );
   nand U26166 ( n26444,n26232,n23393 );
   nand U26167 ( p1_u3224,n26460,n26461,n26462,n26463 );
   nor U26168 ( n26463,n25466,n26464,n26465 );
   nor U26169 ( n26465,n23796,n26222 );
   nor U26170 ( n26464,n23820,n26261 );
   nor U26171 ( n25466,p1_state_reg,n26466 );
   nand U26172 ( n26462,n26467,n26223 );
   nand U26173 ( n26461,n26244,n26468 );
   xor U26174 ( n26468,n26469,n26470 );
   xor U26175 ( n26469,n26471,n26472 );
   nand U26176 ( n26460,n26225,n23822 );
   nand U26177 ( p1_u3223,n26473,n26474,n26475,n26476 );
   nor U26178 ( n26476,n26477,n26478,n26479 );
   nor U26179 ( n26479,n23728,n26261 );
   nor U26180 ( n26478,n26240,n24895 );
   not U26181 ( n24895,n26480 );
   and U26182 ( n26477,p1_u3086,p1_reg3_reg_21_ );
   nand U26183 ( n26475,n26225,n24917 );
   nand U26184 ( n26474,n26481,n26482,n26244 );
   nand U26185 ( n26482,n26483,n26356,n26484 );
   nand U26186 ( n26484,n26485,n26486 );
   nand U26187 ( n26483,n26352,n26355 );
   not U26188 ( n26352,n26487 );
   nand U26189 ( n26481,n26488,n26485,n26489 );
   nand U26190 ( n26488,n26487,n26356 );
   nand U26191 ( n26487,n26490,n26491 );
   nand U26192 ( n26491,n26492,n26493 );
   nand U26193 ( n26473,n26299,n23399 );
   nand U26194 ( p1_u3222,n26494,n26495,n26496,n26497 );
   nand U26195 ( n26497,n26225,n24296 );
   nor U26196 ( n26496,n26498,n26499 );
   nor U26197 ( n26499,n26289,n24301 );
   not U26198 ( n24301,p1_reg3_reg_1_ );
   not U26199 ( n26289,n26361 );
   nand U26200 ( n26361,n26240,p1_state_reg );
   nor U26201 ( n26498,n26500,n26227 );
   xor U26202 ( n26500,n26501,n26502 );
   xor U26203 ( n26501,n26503,n26504 );
   nand U26204 ( n26495,n26299,n23459 );
   nand U26205 ( n26494,n26232,n23465 );
   nand U26206 ( p1_u3221,n26505,n26506,n26507,n26508 );
   nor U26207 ( n26508,n25564,n26509,n26510 );
   nor U26208 ( n26510,n24516,n26261 );
   not U26209 ( n24516,n23444 );
   nor U26210 ( n26509,n26240,n24499 );
   nor U26211 ( n25564,p1_state_reg,n26511 );
   nand U26212 ( n26507,n26299,n23438 );
   or U26213 ( n26506,n26512,n26227 );
   xor U26214 ( n26512,n26513,n26514 );
   xor U26215 ( n26513,n26515,n26516 );
   nand U26216 ( n26505,n26225,n24525 );
   nand U26217 ( p1_u3220,n26517,n26518,n26519,n26520 );
   nor U26218 ( n26520,n26521,n26522,n26523 );
   nor U26219 ( n26523,n23607,n26261 );
   not U26220 ( n23607,n23384 );
   nor U26221 ( n26522,n26240,n25111 );
   nor U26222 ( n26521,p1_state_reg,n26524 );
   nand U26223 ( n26519,n26225,n23609 );
   nand U26224 ( n26518,n26525,n26526,n26244 );
   nand U26225 ( n26526,n26527,n26528 );
   nand U26226 ( n26528,n26529,n26530 );
   or U26227 ( n26530,n26531,n26532 );
   not U26228 ( n26527,n26533 );
   nand U26229 ( n26525,n26533,n26534 );
   nand U26230 ( n26534,n26535,n26536 );
   nand U26231 ( n26536,n26531,n26529 );
   not U26232 ( n26529,n26537 );
   xor U26233 ( n26533,n26538,n26539 );
   nand U26234 ( n26539,n26540,n26541 );
   nand U26235 ( n26541,n26542,n23609 );
   nand U26236 ( n26540,n26543,n23381 );
   xor U26237 ( n26538,n26544,n26364 );
   nand U26238 ( n26544,n26545,n26546 );
   nand U26239 ( n26546,n26547,n23609 );
   nand U26240 ( n23609,n26548,n26549 );
   nand U26241 ( n26549,n26136,n20853 );
   xor U26242 ( n20853,n26206,n26550 );
   xor U26243 ( n26550,si_28_,n26205 );
   nand U26244 ( n26205,n26551,n26552 );
   nand U26245 ( n26552,n26553,n26554 );
   not U26246 ( n26554,si_27_ );
   or U26247 ( n26553,n26555,n26556 );
   nand U26248 ( n26551,n26556,n26555 );
   nand U26249 ( n26206,n26557,n26558 );
   or U26250 ( n26558,n16572,p2_datao_reg_28_ );
   nand U26251 ( n26557,n16572,n17683 );
   not U26252 ( n17683,p1_datao_reg_28_ );
   nand U26253 ( n26548,n26140,p2_datao_reg_28_ );
   nand U26254 ( n26545,n26542,n23381 );
   nand U26255 ( n26517,n26299,n23378 );
   nand U26256 ( n23378,n26559,n26560,n26561,n26562 );
   nand U26257 ( n26562,n26563,n24007 );
   nor U26258 ( n24007,n26564,n26565,n26524 );
   nand U26259 ( n26561,p1_reg0_reg_29_,n26178 );
   nand U26260 ( n26560,p1_reg1_reg_29_,n26179 );
   nand U26261 ( n26559,p1_reg2_reg_29_,n26177 );
   nand U26262 ( p1_u3219,n26566,n26567,n26568,n26569 );
   nor U26263 ( n26569,n25278,n26570,n26571 );
   nor U26264 ( n26571,n23728,n26222 );
   not U26265 ( n23728,n23405 );
   nor U26266 ( n26570,n26240,n24843 );
   nor U26267 ( n25278,p1_state_reg,n26572 );
   nand U26268 ( n26568,n26225,n23729 );
   nand U26269 ( n26567,n26244,n26573 );
   nand U26270 ( n26573,n26574,n26575,n26576 );
   nand U26271 ( n26576,n26577,n26578 );
   nand U26272 ( n26575,n26493,n26579,n26580 );
   nand U26273 ( n26574,n26581,n26582 );
   xor U26274 ( n26581,n26493,n26579 );
   nand U26275 ( n26566,n26232,n23411 );
   nand U26276 ( p1_u3218,n26583,n26584,n26585,n26586 );
   nor U26277 ( n26586,n26587,n25706,n26588 );
   nor U26278 ( n26588,p1_reg3_reg_3_,n26240 );
   nor U26279 ( n25706,p1_state_reg,n26589 );
   nor U26280 ( n26587,n23962,n26261 );
   not U26281 ( n23962,n23459 );
   nand U26282 ( n26585,n26299,n23453 );
   nand U26283 ( n26584,n26590,n26591,n26244 );
   nand U26284 ( n26591,n26592,n26293,n26593,n26594 );
   nand U26285 ( n26592,n26595,n26294 );
   nand U26286 ( n26590,n26596,n26597 );
   nand U26287 ( n26597,n26593,n26594 );
   nand U26288 ( n26583,n26225,n23934 );
   nand U26289 ( p1_u3217,n26598,n26599,n26600,n26601 );
   nor U26290 ( n26601,n25518,n26602,n26603 );
   nor U26291 ( n26603,n23820,n26222 );
   not U26292 ( n23820,n23432 );
   nor U26293 ( n26602,n26240,n24558 );
   not U26294 ( n24558,n26604 );
   nor U26295 ( n25518,p1_state_reg,n26605 );
   nand U26296 ( n26600,n26225,n24578 );
   or U26297 ( n26599,n26606,n26227 );
   xor U26298 ( n26606,n26607,n26608 );
   xor U26299 ( n26608,n26609,n26610 );
   nand U26300 ( n26598,n26232,n23438 );
   nand U26301 ( p1_u3216,n26611,n26612,n26613,n26614 );
   nor U26302 ( n26614,n26615,n26616,n26617 );
   nor U26303 ( n26617,n23648,n26222 );
   not U26304 ( n23648,n23393 );
   nor U26305 ( n26616,n26240,n24954 );
   and U26306 ( n26615,p1_u3086,p1_reg3_reg_23_ );
   nand U26307 ( n26613,n26225,n24979 );
   or U26308 ( n26612,n26618,n26227 );
   xor U26309 ( n26618,n26619,n26620 );
   xor U26310 ( n26620,n26621,n26622 );
   nand U26311 ( n26611,n26232,n23399 );
   nand U26312 ( p1_u3215,n26623,n26624,n26625,n26626 );
   nor U26313 ( n26626,n26627,n26628,n26629 );
   nor U26314 ( n26629,n23795,n26222 );
   not U26315 ( n23795,n23420 );
   nor U26316 ( n26628,n23796,n26261 );
   not U26317 ( n23796,n23426 );
   nor U26318 ( n26627,p1_state_reg,n26630 );
   nand U26319 ( n26625,n26631,n26223 );
   or U26320 ( n26624,n26632,n26227 );
   xor U26321 ( n26632,n26633,n26634 );
   xor U26322 ( n26633,n26635,n26636 );
   nand U26323 ( n26623,n26225,n23799 );
   nand U26324 ( p1_u3214,n26637,n26638,n26639,n26640 );
   nor U26325 ( n26640,n26641,n26642,n26643 );
   nor U26326 ( n26643,n23650,n26261 );
   not U26327 ( n23650,n23387 );
   nor U26328 ( n26642,n26240,n25067 );
   nor U26329 ( n26641,p1_state_reg,n26564 );
   nand U26330 ( n26639,n26225,n25089 );
   nand U26331 ( n26638,n26644,n26244 );
   xor U26332 ( n26644,n26645,n26531 );
   nand U26333 ( n26531,n26248,n26646 );
   nand U26334 ( n26646,n26253,n26647 );
   nand U26335 ( n26647,n26246,n26403,n26459 );
   nand U26336 ( n26459,n26648,n26404 );
   nand U26337 ( n26404,n26649,n26650 );
   not U26338 ( n26650,n26651 );
   xor U26339 ( n26649,n26652,n26653 );
   not U26340 ( n26648,n26402 );
   nand U26341 ( n26402,n26654,n26655 );
   nand U26342 ( n26655,n26619,n26656 );
   or U26343 ( n26656,n26622,n26621 );
   xor U26344 ( n26619,n26652,n26657 );
   nand U26345 ( n26657,n26658,n26659 );
   nand U26346 ( n26659,n26547,n24979 );
   nand U26347 ( n26658,n26542,n23396 );
   nand U26348 ( n26654,n26621,n26622 );
   nand U26349 ( n26622,n26660,n26661 );
   nand U26350 ( n26661,n26325,n26662 );
   nand U26351 ( n26662,n26322,n26324 );
   and U26352 ( n26325,n26663,n26485,n26664 );
   nand U26353 ( n26664,n26665,n26486 );
   not U26354 ( n26665,n26356 );
   nand U26355 ( n26356,n26354,n26353 );
   nand U26356 ( n26485,n26666,n26667 );
   xor U26357 ( n26666,n26668,n26364 );
   nand U26358 ( n26663,n26489,n26669 );
   nand U26359 ( n26669,n26492,n26670 );
   nand U26360 ( n26670,n26578,n26490 );
   not U26361 ( n26490,n26577 );
   nor U26362 ( n26577,n26579,n26582 );
   not U26363 ( n26578,n26493 );
   nand U26364 ( n26493,n26671,n26672 );
   nand U26365 ( n26672,n26673,n26282 );
   nand U26366 ( n26282,n26674,n26417 );
   nand U26367 ( n26417,n26675,n26676 );
   not U26368 ( n26676,n26677 );
   xor U26369 ( n26675,n26652,n26678 );
   nand U26370 ( n26674,n26414,n26416 );
   nand U26371 ( n26416,n26679,n26677 );
   nand U26372 ( n26677,n26680,n26681 );
   nand U26373 ( n26681,n26542,n24804 );
   nand U26374 ( n26680,n26543,n23414 );
   xor U26375 ( n26679,n26678,n26364 );
   nand U26376 ( n26678,n26682,n26683 );
   nand U26377 ( n26683,n26547,n24804 );
   nand U26378 ( n24804,n26684,n26685,n26686 );
   nand U26379 ( n26686,n26140,p2_datao_reg_17_ );
   nand U26380 ( n26685,n25344,n25265 );
   not U26381 ( n25344,n25327 );
   nand U26382 ( n25327,n26687,n26688,n24163 );
   nand U26383 ( n26688,n24155,n24254 );
   nand U26384 ( n26687,p1_ir_reg_17_,n24147,p1_ir_reg_31_ );
   nand U26385 ( n26684,n26136,n20761 );
   not U26386 ( n20761,n22955 );
   xor U26387 ( n22955,n26689,n26690 );
   xor U26388 ( n26689,n26691,n26692 );
   nand U26389 ( n26682,n26542,n23414 );
   nand U26390 ( n23414,n26693,n26694,n26695,n26696 );
   nand U26391 ( n26696,n26563,n26697 );
   not U26392 ( n26697,n24788 );
   xor U26393 ( n24788,p1_reg3_reg_17_,n26698 );
   nand U26394 ( n26695,p1_reg0_reg_17_,n26178 );
   nand U26395 ( n26694,p1_reg1_reg_17_,n26179 );
   nand U26396 ( n26693,p1_reg2_reg_17_,n26177 );
   not U26397 ( n26414,n26418 );
   nand U26398 ( n26418,n26699,n26700 );
   nand U26399 ( n26700,n26440,n26701 );
   nand U26400 ( n26701,n26442,n26443 );
   xor U26401 ( n26440,n26364,n26702 );
   nand U26402 ( n26702,n26703,n26704 );
   nand U26403 ( n26704,n26547,n23766 );
   nand U26404 ( n26703,n26542,n23417 );
   or U26405 ( n26699,n26443,n26442 );
   and U26406 ( n26442,n26705,n26706 );
   nand U26407 ( n26706,n26542,n23766 );
   nand U26408 ( n23766,n26707,n26708,n26709 );
   nand U26409 ( n26709,n26140,p2_datao_reg_16_ );
   nand U26410 ( n26708,n25354,n25265 );
   not U26411 ( n25354,n25355 );
   nand U26412 ( n25355,n26710,n26711 );
   or U26413 ( n26711,p1_ir_reg_16_,p1_ir_reg_31_ );
   nand U26414 ( n26710,p1_ir_reg_31_,n26712 );
   nand U26415 ( n26712,n24146,n24147 );
   not U26416 ( n24147,n24154 );
   nand U26417 ( n24146,p1_ir_reg_16_,n26713 );
   nand U26418 ( n26713,n24139,n24141 );
   not U26419 ( n24141,p1_ir_reg_15_ );
   nand U26420 ( n26707,n26136,n20751 );
   not U26421 ( n20751,n23101 );
   xor U26422 ( n23101,n26714,n26715 );
   xor U26423 ( n26714,n26716,n26717 );
   nand U26424 ( n26705,n26543,n23417 );
   nand U26425 ( n23417,n26718,n26719,n26720,n26721 );
   nand U26426 ( n26721,n26722,n26563 );
   not U26427 ( n26722,n24746 );
   nand U26428 ( n24746,n26723,n26698 );
   nand U26429 ( n26723,n26438,n26724 );
   nand U26430 ( n26724,p1_reg3_reg_15_,n26725 );
   not U26431 ( n26438,p1_reg3_reg_16_ );
   nand U26432 ( n26720,p1_reg0_reg_16_,n26178 );
   nand U26433 ( n26719,p1_reg1_reg_16_,n26179 );
   nand U26434 ( n26718,p1_reg2_reg_16_,n26177 );
   nand U26435 ( n26443,n26726,n26727 );
   nand U26436 ( n26727,n26228,n26728 );
   nand U26437 ( n26728,n26231,n26230 );
   xor U26438 ( n26228,n26652,n26729 );
   nand U26439 ( n26729,n26730,n26731 );
   nand U26440 ( n26731,n26547,n24726 );
   nand U26441 ( n26730,n26542,n23420 );
   or U26442 ( n26726,n26230,n26231 );
   and U26443 ( n26231,n26732,n26733 );
   nand U26444 ( n26733,n26734,n26636 );
   nand U26445 ( n26636,n26735,n26338 );
   nand U26446 ( n26338,n26736,n26737 );
   not U26447 ( n26737,n26738 );
   xor U26448 ( n26736,n26652,n26739 );
   nand U26449 ( n26735,n26335,n26337 );
   nand U26450 ( n26337,n26740,n26738 );
   nand U26451 ( n26738,n26741,n26742 );
   nand U26452 ( n26742,n26542,n24676 );
   nand U26453 ( n26741,n26543,n23426 );
   xor U26454 ( n26740,n26739,n26364 );
   nand U26455 ( n26739,n26743,n26744 );
   nand U26456 ( n26744,n26547,n24676 );
   nand U26457 ( n24676,n26745,n26746,n26747 );
   nand U26458 ( n26747,n26140,p2_datao_reg_13_ );
   nand U26459 ( n26746,n25447,n25265 );
   not U26460 ( n25447,n25454 );
   nand U26461 ( n25454,n26748,n26749,n26750 );
   nand U26462 ( n26749,n24126,n24254 );
   nand U26463 ( n26748,p1_ir_reg_13_,n24118,p1_ir_reg_31_ );
   nand U26464 ( n26745,n26136,n20727 );
   xor U26465 ( n20727,n26751,n26752 );
   nand U26466 ( n26752,n26753,n26754,n26755 );
   and U26467 ( n26751,n26756,n26757 );
   nand U26468 ( n26743,n26542,n23426 );
   nand U26469 ( n23426,n26758,n26759,n26760,n26761 );
   nand U26470 ( n26761,n26563,n26762 );
   not U26471 ( n26762,n24658 );
   xor U26472 ( n24658,p1_reg3_reg_13_,n26763 );
   nand U26473 ( n26760,p1_reg0_reg_13_,n26178 );
   nand U26474 ( n26759,p1_reg1_reg_13_,n26179 );
   nand U26475 ( n26758,p1_reg2_reg_13_,n26177 );
   not U26476 ( n26335,n26339 );
   nand U26477 ( n26339,n26764,n26765 );
   nand U26478 ( n26765,n26766,n26472 );
   nand U26479 ( n26472,n26767,n26768 );
   nand U26480 ( n26768,n26542,n23822 );
   nand U26481 ( n26767,n26543,n23429 );
   nand U26482 ( n26766,n26471,n26470 );
   or U26483 ( n26764,n26470,n26471 );
   and U26484 ( n26471,n26769,n26770 );
   nand U26485 ( n26770,n26312,n26771 );
   or U26486 ( n26771,n26311,n26309 );
   and U26487 ( n26312,n26772,n26773 );
   nand U26488 ( n26773,n26607,n26774 );
   or U26489 ( n26774,n26610,n26609 );
   xor U26490 ( n26607,n26652,n26775 );
   nand U26491 ( n26775,n26776,n26777 );
   nand U26492 ( n26777,n26547,n24578 );
   nand U26493 ( n26776,n26542,n23435 );
   nand U26494 ( n26772,n26609,n26610 );
   nand U26495 ( n26610,n26778,n26779 );
   nand U26496 ( n26779,n26374,n26780 );
   or U26497 ( n26780,n26377,n26376 );
   xor U26498 ( n26374,n26652,n26781 );
   nand U26499 ( n26781,n26782,n26783 );
   nand U26500 ( n26783,n26547,n25231 );
   nand U26501 ( n26782,n26542,n23438 );
   nand U26502 ( n26778,n26376,n26377 );
   nand U26503 ( n26377,n26784,n26785 );
   nand U26504 ( n26785,n26786,n26516 );
   nand U26505 ( n26516,n26787,n26788 );
   nand U26506 ( n26787,n26789,n26790 );
   nand U26507 ( n26786,n26514,n26515 );
   or U26508 ( n26784,n26515,n26514 );
   xor U26509 ( n26514,n26364,n26791 );
   nand U26510 ( n26791,n26792,n26793 );
   nand U26511 ( n26793,n26547,n24525 );
   nand U26512 ( n26792,n26542,n23441 );
   nand U26513 ( n26515,n26794,n26795 );
   nand U26514 ( n26795,n26542,n24525 );
   nand U26515 ( n24525,n26796,n26797,n26798 );
   nand U26516 ( n26798,n26140,p2_datao_reg_8_ );
   nand U26517 ( n26797,n25565,n25265 );
   not U26518 ( n25565,n25583 );
   nand U26519 ( n25583,n26799,n26800 );
   or U26520 ( n26800,p1_ir_reg_31_,p1_ir_reg_8_ );
   nand U26521 ( n26799,p1_ir_reg_31_,n26801 );
   nand U26522 ( n26801,n24095,n24096 );
   nand U26523 ( n24095,p1_ir_reg_8_,n26802 );
   nand U26524 ( n26802,n24089,n24090 );
   not U26525 ( n24090,p1_ir_reg_7_ );
   nand U26526 ( n26796,n26136,n20684 );
   xor U26527 ( n20684,n26803,n26804 );
   nand U26528 ( n26804,n26805,n26806 );
   nand U26529 ( n26806,n26807,n26808 );
   and U26530 ( n26803,n26809,n26810 );
   nand U26531 ( n26794,n26543,n23441 );
   and U26532 ( n26376,n26811,n26812 );
   nand U26533 ( n26812,n26543,n23438 );
   nand U26534 ( n23438,n26813,n26814,n26815,n26816 );
   nand U26535 ( n26816,n26563,n24537 );
   xor U26536 ( n24537,n26372,n26817 );
   nand U26537 ( n26815,p1_reg0_reg_9_,n26178 );
   nand U26538 ( n26814,p1_reg1_reg_9_,n26179 );
   nand U26539 ( n26813,p1_reg2_reg_9_,n26177 );
   nand U26540 ( n26811,n26542,n25231 );
   nand U26541 ( n25231,n26818,n26819,n26820 );
   nand U26542 ( n26820,n26140,p2_datao_reg_9_ );
   nand U26543 ( n26819,n25539,n25265 );
   and U26544 ( n25539,n26821,n26822 );
   nand U26545 ( n26822,n24254,n26823 );
   or U26546 ( n26821,n24101,n24254 );
   xor U26547 ( n24101,p1_ir_reg_9_,n24096 );
   nand U26548 ( n26818,n26136,n20693 );
   xor U26549 ( n20693,n26824,n26825 );
   and U26550 ( n26824,n26826,n26827 );
   and U26551 ( n26609,n26828,n26829 );
   nand U26552 ( n26829,n26543,n23435 );
   nand U26553 ( n23435,n26830,n26831,n26832,n26833 );
   nand U26554 ( n26833,n26604,n26563 );
   nor U26555 ( n26604,n26834,n26835 );
   and U26556 ( n26834,n26605,n26836 );
   nand U26557 ( n26836,p1_reg3_reg_9_,n26837 );
   not U26558 ( n26837,n26817 );
   nand U26559 ( n26832,p1_reg0_reg_10_,n26178 );
   nand U26560 ( n26831,p1_reg1_reg_10_,n26179 );
   nand U26561 ( n26830,p1_reg2_reg_10_,n26177 );
   nand U26562 ( n26828,n26542,n24578 );
   nand U26563 ( n24578,n26838,n26839,n26840 );
   nand U26564 ( n26840,n26140,p2_datao_reg_10_ );
   nand U26565 ( n26839,n25519,n25265 );
   not U26566 ( n25519,n25525 );
   nand U26567 ( n25525,n26841,n26842 );
   or U26568 ( n26842,p1_ir_reg_10_,p1_ir_reg_31_ );
   nand U26569 ( n26841,p1_ir_reg_31_,n24107 );
   nand U26570 ( n24107,n26843,n26844 );
   nand U26571 ( n26844,p1_ir_reg_10_,n26845 );
   nand U26572 ( n26845,n26846,n26823 );
   not U26573 ( n26823,p1_ir_reg_9_ );
   nand U26574 ( n26838,n26136,n20700 );
   xor U26575 ( n20700,n26847,n26848 );
   xor U26576 ( n26848,si_10_,n26849 );
   nand U26577 ( n26769,n26309,n26311 );
   nand U26578 ( n26311,n26850,n26851 );
   nand U26579 ( n26851,n26543,n23432 );
   nand U26580 ( n26850,n26542,n24628 );
   xor U26581 ( n26309,n26364,n26852 );
   nand U26582 ( n26852,n26853,n26854 );
   nand U26583 ( n26854,n26547,n24628 );
   nand U26584 ( n24628,n26855,n26856,n26857 );
   nand U26585 ( n26857,n26140,p2_datao_reg_11_ );
   nand U26586 ( n26856,n25481,n25265 );
   not U26587 ( n25481,n25479 );
   nand U26588 ( n25479,n26858,n26859 );
   nand U26589 ( n26859,n26860,n24254 );
   or U26590 ( n26858,n24112,n24254 );
   xor U26591 ( n24112,p1_ir_reg_11_,n26843 );
   nand U26592 ( n26855,n26136,n20710 );
   xor U26593 ( n20710,n26861,n26862 );
   nor U26594 ( n26861,n26863,n26864 );
   nand U26595 ( n26853,n26542,n23432 );
   nand U26596 ( n23432,n26865,n26866,n26867,n26868 );
   nand U26597 ( n26868,n26563,n26307 );
   xor U26598 ( n26307,p1_reg3_reg_11_,n26835 );
   nand U26599 ( n26867,p1_reg0_reg_11_,n26178 );
   nand U26600 ( n26866,p1_reg1_reg_11_,n26179 );
   nand U26601 ( n26865,p1_reg2_reg_11_,n26177 );
   xor U26602 ( n26470,n26652,n26869 );
   nand U26603 ( n26869,n26870,n26871 );
   nand U26604 ( n26871,n26547,n23822 );
   nand U26605 ( n23822,n26872,n26873,n26874 );
   nand U26606 ( n26874,n26140,p2_datao_reg_12_ );
   nand U26607 ( n26873,n25467,n25265 );
   not U26608 ( n25467,n25484 );
   nand U26609 ( n25484,n26875,n26876 );
   or U26610 ( n26876,p1_ir_reg_12_,p1_ir_reg_31_ );
   nand U26611 ( n26875,p1_ir_reg_31_,n26877 );
   nand U26612 ( n26877,n24117,n24118 );
   not U26613 ( n24118,n24125 );
   nand U26614 ( n24117,p1_ir_reg_12_,n26878 );
   nand U26615 ( n26878,n26879,n26860 );
   not U26616 ( n26860,p1_ir_reg_11_ );
   nand U26617 ( n26872,n26136,n20717 );
   xor U26618 ( n20717,n26880,n26881 );
   nand U26619 ( n26881,n26882,n26883 );
   nand U26620 ( n26883,n26884,n26862 );
   and U26621 ( n26880,n26754,n26885 );
   nand U26622 ( n26870,n26542,n23429 );
   nand U26623 ( n23429,n26886,n26887,n26888,n26889 );
   nand U26624 ( n26889,n26467,n26563 );
   not U26625 ( n26467,n24640 );
   nand U26626 ( n24640,n26890,n26763 );
   nand U26627 ( n26890,n26466,n26891 );
   nand U26628 ( n26891,p1_reg3_reg_11_,n26835 );
   not U26629 ( n26466,p1_reg3_reg_12_ );
   nand U26630 ( n26888,p1_reg0_reg_12_,n26178 );
   nand U26631 ( n26887,p1_reg1_reg_12_,n26179 );
   nand U26632 ( n26886,p1_reg2_reg_12_,n26177 );
   nand U26633 ( n26734,n26634,n26635 );
   or U26634 ( n26732,n26635,n26634 );
   xor U26635 ( n26634,n26364,n26892 );
   nand U26636 ( n26892,n26893,n26894 );
   nand U26637 ( n26894,n26547,n23799 );
   nand U26638 ( n26893,n26542,n23423 );
   nand U26639 ( n26635,n26895,n26896 );
   nand U26640 ( n26896,n26542,n23799 );
   nand U26641 ( n23799,n26897,n26898,n26899 );
   nand U26642 ( n26899,n26140,p2_datao_reg_14_ );
   nand U26643 ( n26898,n25425,n25265 );
   not U26644 ( n25425,n25409 );
   nand U26645 ( n25409,n26900,n26901 );
   or U26646 ( n26901,p1_ir_reg_14_,p1_ir_reg_31_ );
   nand U26647 ( n26900,p1_ir_reg_31_,n24132 );
   nand U26648 ( n24132,n24140,n26902 );
   nand U26649 ( n26902,p1_ir_reg_14_,n26750 );
   nand U26650 ( n26897,n26136,n20734 );
   nand U26651 ( n20734,n26903,n26904,n26905 );
   nand U26652 ( n26905,n26906,n26907 );
   or U26653 ( n26904,n26907,n26908,si_14_ );
   nand U26654 ( n26903,n26909,si_14_ );
   xor U26655 ( n26909,n26908,n26907 );
   nand U26656 ( n26907,n26910,n26911 );
   nand U26657 ( n26911,n26912,n26757 );
   nand U26658 ( n26895,n26543,n23423 );
   nand U26659 ( n23423,n26913,n26914,n26915,n26916 );
   nand U26660 ( n26916,n26631,n26563 );
   not U26661 ( n26631,n24704 );
   nand U26662 ( n24704,n26917,n26918 );
   nand U26663 ( n26917,n26630,n26919 );
   or U26664 ( n26919,n26332,n26763 );
   nand U26665 ( n26915,p1_reg0_reg_14_,n26178 );
   nand U26666 ( n26914,p1_reg1_reg_14_,n26179 );
   nand U26667 ( n26913,p1_reg2_reg_14_,n26177 );
   nand U26668 ( n26230,n26920,n26921 );
   nand U26669 ( n26921,n26543,n23420 );
   nand U26670 ( n23420,n26922,n26923,n26924,n26925 );
   nand U26671 ( n26925,n26563,n24736 );
   xor U26672 ( n24736,n26224,n26918 );
   not U26673 ( n26918,n26725 );
   not U26674 ( n26224,p1_reg3_reg_15_ );
   nand U26675 ( n26924,p1_reg0_reg_15_,n26178 );
   nand U26676 ( n26923,p1_reg1_reg_15_,n26179 );
   nand U26677 ( n26922,p1_reg2_reg_15_,n26177 );
   nand U26678 ( n26920,n26542,n24726 );
   nand U26679 ( n24726,n26926,n26927,n26928 );
   nand U26680 ( n26928,n26140,p2_datao_reg_15_ );
   nand U26681 ( n26927,n25265,n25394 );
   not U26682 ( n25394,n25383 );
   xor U26683 ( n25383,p1_ir_reg_15_,n26929 );
   nand U26684 ( n26929,p1_ir_reg_31_,n24140 );
   nand U26685 ( n26926,n26136,n20744 );
   xor U26686 ( n20744,n26930,n26931 );
   xor U26687 ( n26930,n26932,n26933 );
   nand U26688 ( n26932,n26934,n26935 );
   nand U26689 ( n26935,n26757,n26936,n26912 );
   nand U26690 ( n26673,n26280,n26281 );
   or U26691 ( n26671,n26281,n26280 );
   xor U26692 ( n26280,n26364,n26937 );
   nand U26693 ( n26937,n26938,n26939 );
   nand U26694 ( n26939,n26547,n23745 );
   nand U26695 ( n26938,n26542,n23411 );
   nand U26696 ( n26281,n26940,n26941 );
   nand U26697 ( n26941,n26542,n23745 );
   nand U26698 ( n23745,n26942,n26943,n26944 );
   nand U26699 ( n26944,n26140,p2_datao_reg_18_ );
   nand U26700 ( n26943,n25294,n25265 );
   not U26701 ( n25294,n25293 );
   nand U26702 ( n25293,n26945,n26946,n26947 );
   nand U26703 ( n26946,n24164,n24254 );
   nand U26704 ( n26945,p1_ir_reg_18_,n24163,p1_ir_reg_31_ );
   nand U26705 ( n26942,n26136,n20768 );
   not U26706 ( n20768,n23123 );
   xor U26707 ( n23123,n26948,n26949 );
   xor U26708 ( n26948,n26950,n26951 );
   nand U26709 ( n26940,n26543,n23411 );
   nand U26710 ( n23411,n26952,n26953,n26954,n26955 );
   nand U26711 ( n26955,n26277,n26563 );
   not U26712 ( n26277,n24823 );
   nand U26713 ( n24823,n26956,n26957 );
   nand U26714 ( n26956,n26276,n26958 );
   nand U26715 ( n26958,p1_reg3_reg_17_,n26959 );
   not U26716 ( n26276,p1_reg3_reg_18_ );
   nand U26717 ( n26954,p1_reg0_reg_18_,n26178 );
   nand U26718 ( n26953,p1_reg1_reg_18_,n26179 );
   nand U26719 ( n26952,p1_reg2_reg_18_,n26177 );
   nand U26720 ( n26492,n26582,n26579 );
   nand U26721 ( n26579,n26960,n26961 );
   nand U26722 ( n26961,n26542,n23729 );
   nand U26723 ( n26960,n26543,n23408 );
   not U26724 ( n26582,n26580 );
   xor U26725 ( n26580,n26652,n26962 );
   nand U26726 ( n26962,n26963,n26964 );
   nand U26727 ( n26964,n26547,n23729 );
   nand U26728 ( n23729,n26965,n26966,n26967 );
   nand U26729 ( n26967,n25265,n23979 );
   nand U26730 ( n26966,n26136,n20778 );
   xor U26731 ( n20778,n26968,n26969 );
   xor U26732 ( n26969,si_19_,n26970 );
   nand U26733 ( n26965,n26140,p2_datao_reg_19_ );
   nand U26734 ( n26963,n26542,n23408 );
   nand U26735 ( n23408,n26971,n26972,n26973,n26974 );
   nand U26736 ( n26974,n26563,n26975 );
   not U26737 ( n26975,n24843 );
   xor U26738 ( n24843,p1_reg3_reg_19_,n26957 );
   nand U26739 ( n26973,p1_reg0_reg_19_,n26178 );
   nand U26740 ( n26972,p1_reg1_reg_19_,n26179 );
   nand U26741 ( n26971,p1_reg2_reg_19_,n26177 );
   and U26742 ( n26489,n26486,n26355 );
   or U26743 ( n26355,n26353,n26354 );
   xor U26744 ( n26354,n26364,n26976 );
   nand U26745 ( n26976,n26977,n26978 );
   nand U26746 ( n26978,n26547,n24876 );
   nand U26747 ( n26977,n26542,n23405 );
   nand U26748 ( n26353,n26979,n26980 );
   nand U26749 ( n26980,n26542,n24876 );
   nand U26750 ( n24876,n26981,n26982 );
   nand U26751 ( n26982,n26136,n20785 );
   xor U26752 ( n20785,n26983,n26984 );
   xor U26753 ( n26984,si_20_,n26985 );
   nand U26754 ( n26981,n26140,p2_datao_reg_20_ );
   nand U26755 ( n26979,n26543,n23405 );
   nand U26756 ( n23405,n26986,n26987,n26988,n26989 );
   nand U26757 ( n26989,n26347,n26563 );
   nor U26758 ( n26347,n26990,n26991 );
   and U26759 ( n26990,n26348,n26992 );
   nand U26760 ( n26992,p1_reg3_reg_19_,n26993 );
   not U26761 ( n26993,n26957 );
   nand U26762 ( n26988,p1_reg0_reg_20_,n26178 );
   nand U26763 ( n26987,p1_reg1_reg_20_,n26179 );
   nand U26764 ( n26986,p1_reg2_reg_20_,n26177 );
   nand U26765 ( n26486,n26994,n26995 );
   not U26766 ( n26995,n26667 );
   nand U26767 ( n26667,n26996,n26997 );
   nand U26768 ( n26997,n26542,n24917 );
   nand U26769 ( n26996,n26543,n23402 );
   xor U26770 ( n26994,n26652,n26668 );
   nand U26771 ( n26668,n26998,n26999 );
   nand U26772 ( n26999,n26547,n24917 );
   nand U26773 ( n24917,n27000,n27001 );
   nand U26774 ( n27001,n26136,n20794 );
   xor U26775 ( n20794,n27002,n27003 );
   xor U26776 ( n27003,si_21_,n27004 );
   nand U26777 ( n27000,n26140,p2_datao_reg_21_ );
   nand U26778 ( n26998,n26542,n23402 );
   nand U26779 ( n23402,n27005,n27006,n27007,n27008 );
   nand U26780 ( n27008,n26563,n26480 );
   xor U26781 ( n26480,p1_reg3_reg_21_,n26991 );
   nand U26782 ( n27007,p1_reg0_reg_21_,n26178 );
   nand U26783 ( n27006,p1_reg1_reg_21_,n26179 );
   nand U26784 ( n27005,p1_reg2_reg_21_,n26177 );
   or U26785 ( n26660,n26324,n26322 );
   xor U26786 ( n26322,n26364,n27009 );
   nand U26787 ( n27009,n27010,n27011 );
   nand U26788 ( n27011,n26547,n24934 );
   nand U26789 ( n27010,n26542,n23399 );
   nand U26790 ( n26324,n27012,n27013 );
   nand U26791 ( n27013,n26543,n23399 );
   nand U26792 ( n23399,n27014,n27015,n27016,n27017 );
   nand U26793 ( n27017,n24945,n26563 );
   and U26794 ( n24945,n27018,n27019 );
   nand U26795 ( n27018,n26320,n27020 );
   nand U26796 ( n27020,p1_reg3_reg_21_,n26991 );
   not U26797 ( n26320,p1_reg3_reg_22_ );
   nand U26798 ( n27016,p1_reg0_reg_22_,n26178 );
   nand U26799 ( n27015,p1_reg1_reg_22_,n26179 );
   nand U26800 ( n27014,p1_reg2_reg_22_,n26177 );
   nand U26801 ( n27012,n26542,n24934 );
   nand U26802 ( n24934,n27021,n27022 );
   nand U26803 ( n27022,n26136,n20804 );
   xor U26804 ( n20804,n27023,n27024 );
   xor U26805 ( n27024,si_22_,n27025 );
   nand U26806 ( n27021,n26140,p2_datao_reg_22_ );
   and U26807 ( n26621,n27026,n27027 );
   nand U26808 ( n27027,n26543,n23396 );
   nand U26809 ( n23396,n27028,n27029,n27030,n27031 );
   nand U26810 ( n27031,n26563,n27032 );
   not U26811 ( n27032,n24954 );
   xor U26812 ( n24954,p1_reg3_reg_23_,n27019 );
   nand U26813 ( n27030,p1_reg0_reg_23_,n26178 );
   nand U26814 ( n27029,p1_reg1_reg_23_,n26179 );
   nand U26815 ( n27028,p1_reg2_reg_23_,n26177 );
   nand U26816 ( n27026,n26542,n24979 );
   nand U26817 ( n24979,n27033,n27034 );
   nand U26818 ( n27034,n26136,n20811 );
   xor U26819 ( n20811,n27035,n27036 );
   xor U26820 ( n27036,si_23_,n27037 );
   nand U26821 ( n27033,n26140,p2_datao_reg_23_ );
   nand U26822 ( n26403,n27038,n26651 );
   nand U26823 ( n26651,n27039,n27040 );
   nand U26824 ( n27040,n26542,n24994 );
   nand U26825 ( n27039,n26543,n23393 );
   xor U26826 ( n27038,n26653,n26364 );
   nand U26827 ( n26653,n27041,n27042 );
   nand U26828 ( n27042,n26547,n24994 );
   nand U26829 ( n24994,n27043,n27044 );
   nand U26830 ( n27044,n26136,n20818 );
   xor U26831 ( n20818,n27045,n27046 );
   xor U26832 ( n27046,si_24_,n27047 );
   nand U26833 ( n27043,n26140,p2_datao_reg_24_ );
   nand U26834 ( n27041,n26542,n23393 );
   nand U26835 ( n23393,n27048,n27049,n27050,n27051 );
   nand U26836 ( n27051,n27052,n26563 );
   not U26837 ( n27052,n24989 );
   nand U26838 ( n24989,n27053,n27054 );
   nand U26839 ( n27053,n26399,n27055 );
   nand U26840 ( n27055,p1_reg3_reg_23_,n27056 );
   not U26841 ( n26399,p1_reg3_reg_24_ );
   nand U26842 ( n27050,p1_reg0_reg_24_,n26178 );
   nand U26843 ( n27049,p1_reg1_reg_24_,n26179 );
   nand U26844 ( n27048,p1_reg2_reg_24_,n26177 );
   nand U26845 ( n26246,n27057,n26456 );
   not U26846 ( n27057,n26455 );
   and U26847 ( n26253,n26249,n26250 );
   nand U26848 ( n26250,n26458,n26455 );
   xor U26849 ( n26455,n26652,n27058 );
   nand U26850 ( n27058,n27059,n27060 );
   nand U26851 ( n27060,n26547,n25194 );
   nand U26852 ( n27059,n26542,n23390 );
   not U26853 ( n26458,n26456 );
   nand U26854 ( n26456,n27061,n27062 );
   nand U26855 ( n27062,n26542,n25194 );
   nand U26856 ( n25194,n27063,n27064 );
   nand U26857 ( n27064,n26136,n20827 );
   xor U26858 ( n20827,n27065,n27066 );
   xor U26859 ( n27066,si_25_,n27067 );
   nand U26860 ( n27063,n26140,p2_datao_reg_25_ );
   nand U26861 ( n27061,n26543,n23390 );
   nand U26862 ( n23390,n27068,n27069,n27070,n27071 );
   nand U26863 ( n27071,n26563,n27072 );
   not U26864 ( n27072,n25006 );
   xor U26865 ( n25006,p1_reg3_reg_25_,n27054 );
   nand U26866 ( n27070,p1_reg0_reg_25_,n26178 );
   nand U26867 ( n27069,p1_reg1_reg_25_,n26179 );
   nand U26868 ( n27068,p1_reg2_reg_25_,n26177 );
   nand U26869 ( n26249,n27073,n27074,n27075 );
   xor U26870 ( n27075,n26652,n27076 );
   nand U26871 ( n26248,n27077,n27078 );
   nand U26872 ( n27078,n27073,n27074 );
   nand U26873 ( n27074,n26542,n25047 );
   nand U26874 ( n27073,n26543,n23387 );
   xor U26875 ( n27077,n27076,n26364 );
   nand U26876 ( n27076,n27079,n27080 );
   nand U26877 ( n27080,n26547,n25047 );
   nand U26878 ( n25047,n27081,n27082 );
   nand U26879 ( n27082,n26136,n20834 );
   xor U26880 ( n20834,n27083,n27084 );
   xor U26881 ( n27084,si_26_,n27085 );
   nand U26882 ( n27081,n26140,p2_datao_reg_26_ );
   nand U26883 ( n27079,n26542,n23387 );
   nand U26884 ( n23387,n27086,n27087,n27088,n27089 );
   nand U26885 ( n27089,n27090,n26563 );
   not U26886 ( n27090,n25024 );
   nand U26887 ( n25024,n26565,n27091 );
   nand U26888 ( n27091,n27092,n26241 );
   nand U26889 ( n27088,p1_reg0_reg_26_,n26178 );
   nand U26890 ( n27087,p1_reg1_reg_26_,n26179 );
   nand U26891 ( n27086,p1_reg2_reg_26_,n26177 );
   nor U26892 ( n26645,n26532,n26537 );
   nor U26893 ( n26537,n27093,n27094 );
   not U26894 ( n26532,n26535 );
   nand U26895 ( n26535,n27094,n27093 );
   nand U26896 ( n27093,n27095,n27096 );
   nand U26897 ( n27096,n26542,n25089 );
   nand U26898 ( n27095,n26543,n23384 );
   xor U26899 ( n27094,n26364,n27097 );
   nand U26900 ( n27097,n27098,n27099 );
   nand U26901 ( n27099,n26547,n25089 );
   nand U26902 ( n25089,n27100,n27101 );
   nand U26903 ( n27101,n26136,n20843 );
   xor U26904 ( n20843,n26556,n27102 );
   xor U26905 ( n27102,si_27_,n26555 );
   nand U26906 ( n26555,n27103,n27104 );
   nand U26907 ( n27104,n27105,n27106 );
   not U26908 ( n27106,si_26_ );
   or U26909 ( n27105,n27085,n27083 );
   nand U26910 ( n27103,n27083,n27085 );
   nand U26911 ( n27085,n27107,n27108 );
   nand U26912 ( n27108,n27109,n27110 );
   not U26913 ( n27110,si_25_ );
   or U26914 ( n27109,n27067,n27065 );
   nand U26915 ( n27107,n27065,n27067 );
   nand U26916 ( n27067,n27111,n27112 );
   nand U26917 ( n27112,n27113,n27114 );
   not U26918 ( n27114,si_24_ );
   or U26919 ( n27113,n27047,n27045 );
   nand U26920 ( n27111,n27045,n27047 );
   nand U26921 ( n27047,n27115,n27116 );
   nand U26922 ( n27116,n27117,n27118 );
   not U26923 ( n27118,si_23_ );
   or U26924 ( n27117,n27037,n27035 );
   nand U26925 ( n27115,n27035,n27037 );
   nand U26926 ( n27037,n27119,n27120 );
   nand U26927 ( n27120,n27121,n27122 );
   not U26928 ( n27122,si_22_ );
   or U26929 ( n27121,n27025,n27023 );
   nand U26930 ( n27119,n27023,n27025 );
   nand U26931 ( n27025,n27123,n27124 );
   nand U26932 ( n27124,n27125,n27126 );
   not U26933 ( n27126,si_21_ );
   or U26934 ( n27125,n27004,n27002 );
   nand U26935 ( n27123,n27002,n27004 );
   nand U26936 ( n27004,n27127,n27128 );
   nand U26937 ( n27128,n27129,n27130 );
   not U26938 ( n27130,si_20_ );
   or U26939 ( n27129,n26985,n26983 );
   nand U26940 ( n27127,n26983,n26985 );
   nand U26941 ( n26985,n27131,n27132 );
   nand U26942 ( n27132,n27133,n27134 );
   not U26943 ( n27134,si_19_ );
   or U26944 ( n27133,n26970,n26968 );
   nand U26945 ( n27131,n26968,n26970 );
   nand U26946 ( n26970,n27135,n27136 );
   nand U26947 ( n27136,n27137,n26951 );
   not U26948 ( n26951,si_18_ );
   or U26949 ( n27137,n26950,n26949 );
   nand U26950 ( n27135,n26949,n26950 );
   nand U26951 ( n26950,n27138,n27139 );
   nand U26952 ( n27139,n27140,n26692 );
   not U26953 ( n26692,si_17_ );
   or U26954 ( n27140,n26691,n26690 );
   nand U26955 ( n27138,n26690,n26691 );
   nand U26956 ( n26691,n27141,n27142 );
   nand U26957 ( n27142,n27143,n26717 );
   not U26958 ( n26717,si_16_ );
   nand U26959 ( n27143,n26715,n26716 );
   or U26960 ( n27141,n26716,n26715 );
   nand U26961 ( n26715,n27144,n27145 );
   nand U26962 ( n27145,n16572,p1_datao_reg_16_ );
   nand U26963 ( n27144,n16576,p2_datao_reg_16_ );
   nand U26964 ( n26716,n27146,n27147,n27148 );
   or U26965 ( n27148,n26934,n26931 );
   nand U26966 ( n27147,n26912,n27149,n26757,n26936 );
   nand U26967 ( n27149,n26931,n26933 );
   not U26968 ( n26933,si_15_ );
   not U26969 ( n26912,n26755 );
   nand U26970 ( n26755,n26862,n26885,n26884 );
   not U26971 ( n26884,n26863 );
   nor U26972 ( n26863,n27150,si_11_ );
   nand U26973 ( n26862,n27151,n27152 );
   nand U26974 ( n27152,si_10_,n27153 );
   or U26975 ( n27153,n26849,n26847 );
   nand U26976 ( n27151,n26847,n26849 );
   nand U26977 ( n26849,n26826,n27154 );
   nand U26978 ( n27154,n26825,n26827 );
   nand U26979 ( n26827,n27155,n27156,n27157 );
   not U26980 ( n27157,si_9_ );
   nand U26981 ( n27156,n16572,p1_datao_reg_9_ );
   nand U26982 ( n27155,n16576,p2_datao_reg_9_ );
   nand U26983 ( n26825,n27158,n26809,n27159 );
   nand U26984 ( n27159,n27160,n26810 );
   nand U26985 ( n26809,n27161,n27162,si_8_ );
   nand U26986 ( n27162,n16576,n19258 );
   not U26987 ( n19258,p2_datao_reg_8_ );
   nand U26988 ( n27161,n16572,n19259 );
   not U26989 ( n19259,p1_datao_reg_8_ );
   nand U26990 ( n27158,n26807,n26808,n26810 );
   nand U26991 ( n26810,n27163,n27164,n27165 );
   not U26992 ( n27165,si_8_ );
   nand U26993 ( n27164,n16572,p1_datao_reg_8_ );
   nand U26994 ( n27163,n16576,p2_datao_reg_8_ );
   not U26995 ( n26808,n27166 );
   nand U26996 ( n26826,n27167,n27168,si_9_ );
   or U26997 ( n27168,n16572,p2_datao_reg_9_ );
   nand U26998 ( n27167,n16572,n19253 );
   not U26999 ( n19253,p1_datao_reg_9_ );
   and U27000 ( n26847,n27169,n27170 );
   nand U27001 ( n27170,n16576,n19252 );
   not U27002 ( n19252,p2_datao_reg_10_ );
   nand U27003 ( n27169,n16572,n19027 );
   not U27004 ( n19027,p1_datao_reg_10_ );
   nand U27005 ( n27146,si_15_,n27171 );
   nand U27006 ( n27171,n26931,n26934 );
   nand U27007 ( n26934,n26936,n27172 );
   nand U27008 ( n27172,n26910,n27173 );
   nand U27009 ( n27173,n27174,si_14_ );
   and U27010 ( n26910,n27175,n26756 );
   nand U27011 ( n26756,n27176,n27177,si_13_ );
   or U27012 ( n27177,n16572,p2_datao_reg_13_ );
   nand U27013 ( n27176,n16572,n19070 );
   not U27014 ( n19070,p1_datao_reg_13_ );
   nand U27015 ( n27175,n26757,n27178 );
   nand U27016 ( n27178,n26753,n26754 );
   nand U27017 ( n26754,n27179,n27180,si_12_ );
   nand U27018 ( n27180,n16576,n19244 );
   not U27019 ( n19244,p2_datao_reg_12_ );
   nand U27020 ( n27179,n16572,n19245 );
   not U27021 ( n19245,p1_datao_reg_12_ );
   nand U27022 ( n26753,n26864,n26885 );
   nand U27023 ( n26885,n27181,n27182,n27183 );
   not U27024 ( n27183,si_12_ );
   nand U27025 ( n27182,n16572,p1_datao_reg_12_ );
   nand U27026 ( n27181,n16576,p2_datao_reg_12_ );
   not U27027 ( n26864,n26882 );
   nand U27028 ( n26882,si_11_,n27150 );
   nand U27029 ( n27150,n27184,n27185 );
   nand U27030 ( n27185,n16572,p1_datao_reg_11_ );
   nand U27031 ( n27184,n16576,p2_datao_reg_11_ );
   nand U27032 ( n26757,n27186,n27187,n27188 );
   not U27033 ( n27188,si_13_ );
   nand U27034 ( n27187,n16572,p1_datao_reg_13_ );
   nand U27035 ( n27186,n16576,p2_datao_reg_13_ );
   not U27036 ( n26936,n26906 );
   nor U27037 ( n26906,n27174,si_14_ );
   not U27038 ( n27174,n26908 );
   nand U27039 ( n26908,n27189,n27190 );
   or U27040 ( n27190,n16572,p2_datao_reg_14_ );
   nand U27041 ( n27189,n16572,n19237 );
   not U27042 ( n19237,p1_datao_reg_14_ );
   nand U27043 ( n26931,n27191,n27192 );
   or U27044 ( n27192,n16572,p2_datao_reg_15_ );
   nand U27045 ( n27191,n16572,n19233 );
   not U27046 ( n19233,p1_datao_reg_15_ );
   nand U27047 ( n26690,n27193,n27194 );
   or U27048 ( n27194,n16572,p2_datao_reg_17_ );
   nand U27049 ( n27193,n16572,n19225 );
   not U27050 ( n19225,p1_datao_reg_17_ );
   nand U27051 ( n26949,n27195,n27196 );
   or U27052 ( n27196,n16572,p2_datao_reg_18_ );
   nand U27053 ( n27195,n16572,n19221 );
   not U27054 ( n19221,p1_datao_reg_18_ );
   nand U27055 ( n26968,n27197,n27198 );
   or U27056 ( n27198,n16572,p2_datao_reg_19_ );
   nand U27057 ( n27197,n16572,n19217 );
   not U27058 ( n19217,p1_datao_reg_19_ );
   nand U27059 ( n26983,n27199,n27200 );
   or U27060 ( n27200,n16572,p2_datao_reg_20_ );
   nand U27061 ( n27199,n16572,n19213 );
   not U27062 ( n19213,p1_datao_reg_20_ );
   nand U27063 ( n27002,n27201,n27202 );
   or U27064 ( n27202,n16572,p2_datao_reg_21_ );
   nand U27065 ( n27201,n16572,n19209 );
   not U27066 ( n19209,p1_datao_reg_21_ );
   nand U27067 ( n27023,n27203,n27204 );
   or U27068 ( n27204,n16572,p2_datao_reg_22_ );
   nand U27069 ( n27203,n16572,n19205 );
   not U27070 ( n19205,p1_datao_reg_22_ );
   nand U27071 ( n27035,n27205,n27206 );
   or U27072 ( n27206,n16572,p2_datao_reg_23_ );
   nand U27073 ( n27205,n16572,n19201 );
   not U27074 ( n19201,p1_datao_reg_23_ );
   nand U27075 ( n27045,n27207,n27208 );
   or U27076 ( n27208,n16572,p2_datao_reg_24_ );
   nand U27077 ( n27207,n16572,n19197 );
   not U27078 ( n19197,p1_datao_reg_24_ );
   nand U27079 ( n27065,n27209,n27210 );
   or U27080 ( n27210,n16572,p2_datao_reg_25_ );
   nand U27081 ( n27209,n16572,n19193 );
   not U27082 ( n19193,p1_datao_reg_25_ );
   nand U27083 ( n27083,n27211,n27212 );
   or U27084 ( n27212,n16572,p2_datao_reg_26_ );
   nand U27085 ( n27211,n16572,n19189 );
   not U27086 ( n19189,p1_datao_reg_26_ );
   nand U27087 ( n26556,n27213,n27214 );
   or U27088 ( n27214,n16572,p2_datao_reg_27_ );
   nand U27089 ( n27213,n16572,n18763 );
   not U27090 ( n18763,p1_datao_reg_27_ );
   nand U27091 ( n27100,n26140,p2_datao_reg_27_ );
   nand U27092 ( n27098,n26542,n23384 );
   nand U27093 ( n23384,n27215,n27216,n27217,n27218 );
   nand U27094 ( n27218,n26563,n27219 );
   not U27095 ( n27219,n25067 );
   xor U27096 ( n25067,p1_reg3_reg_27_,n26565 );
   nand U27097 ( n27217,p1_reg0_reg_27_,n26178 );
   nand U27098 ( n27216,p1_reg1_reg_27_,n26179 );
   nand U27099 ( n27215,p1_reg2_reg_27_,n26177 );
   nand U27100 ( n26637,n26299,n23381 );
   nand U27101 ( n23381,n27220,n27221,n27222,n27223 );
   nand U27102 ( n27223,n26563,n27224 );
   not U27103 ( n27224,n25111 );
   xor U27104 ( n25111,n27225,n26524 );
   not U27105 ( n26524,p1_reg3_reg_28_ );
   nor U27106 ( n27225,n26565,n26564 );
   not U27107 ( n26564,p1_reg3_reg_27_ );
   or U27108 ( n26565,n26241,n27092 );
   nand U27109 ( n27092,p1_reg3_reg_25_,n27226 );
   not U27110 ( n27226,n27054 );
   nand U27111 ( n27054,p1_reg3_reg_23_,n27056,p1_reg3_reg_24_ );
   not U27112 ( n27056,n27019 );
   nand U27113 ( n27019,p1_reg3_reg_21_,n26991,p1_reg3_reg_22_ );
   nor U27114 ( n26991,n26572,n26957,n26348 );
   not U27115 ( n26348,p1_reg3_reg_20_ );
   nand U27116 ( n26957,p1_reg3_reg_17_,n26959,p1_reg3_reg_18_ );
   not U27117 ( n26959,n26698 );
   nand U27118 ( n26698,p1_reg3_reg_15_,n26725,p1_reg3_reg_16_ );
   nor U27119 ( n26725,n26332,n26763,n26630 );
   not U27120 ( n26630,p1_reg3_reg_14_ );
   nand U27121 ( n26763,p1_reg3_reg_11_,n26835,p1_reg3_reg_12_ );
   nor U27122 ( n26835,n26605,n26817,n26372 );
   not U27123 ( n26372,p1_reg3_reg_9_ );
   not U27124 ( n26605,p1_reg3_reg_10_ );
   not U27125 ( n26332,p1_reg3_reg_13_ );
   not U27126 ( n26572,p1_reg3_reg_19_ );
   not U27127 ( n26241,p1_reg3_reg_26_ );
   nand U27128 ( n27222,p1_reg0_reg_28_,n26178 );
   nand U27129 ( n27221,p1_reg1_reg_28_,n26179 );
   nand U27130 ( n27220,p1_reg2_reg_28_,n26177 );
   nand U27131 ( p1_u3213,n27227,n27228,n27229,n27230 );
   nor U27132 ( n27230,n25589,n27231,n27232 );
   nor U27133 ( n27232,n24471,n26261 );
   not U27134 ( n26261,n26232 );
   nor U27135 ( n26232,n26214,n25264,n27233 );
   nor U27136 ( n27231,n23857,n26222 );
   nor U27137 ( n26299,n25106,n26214,n27233 );
   not U27138 ( n23857,n23441 );
   nand U27139 ( n23441,n27234,n27235,n27236,n27237 );
   nand U27140 ( n27237,n27238,n26563 );
   not U27141 ( n27238,n24499 );
   nand U27142 ( n24499,n27239,n26817 );
   nand U27143 ( n26817,p1_reg3_reg_7_,n27240,p1_reg3_reg_8_ );
   nand U27144 ( n27239,n26511,n27241 );
   nand U27145 ( n27241,p1_reg3_reg_7_,n27240 );
   not U27146 ( n27240,n27242 );
   not U27147 ( n26511,p1_reg3_reg_8_ );
   nand U27148 ( n27236,p1_reg0_reg_8_,n26178 );
   nand U27149 ( n27235,p1_reg1_reg_8_,n26179 );
   nand U27150 ( n27234,p1_reg2_reg_8_,n26177 );
   nor U27151 ( n25589,p1_state_reg,n27243 );
   nand U27152 ( n27229,n24459,n26223 );
   nand U27153 ( n26223,n27244,n27245,n25779,n23371 );
   not U27154 ( n25779,n25794 );
   nor U27155 ( n25794,n25791,p1_u3086 );
   nand U27156 ( n27245,n27246,n27233 );
   nand U27157 ( n27246,n26214,n27247 );
   nand U27158 ( n27247,n23566,n27248 );
   or U27159 ( n27248,n27249,n25267 );
   nand U27160 ( n26214,n23566,n25787,n25805 );
   nand U27161 ( n27244,n27250,n23566 );
   not U27162 ( n27250,n25272 );
   nand U27163 ( n25272,n25105,n23984 );
   nand U27164 ( n27228,n27251,n27252,n26244 );
   not U27165 ( n26244,n26227 );
   nand U27166 ( n26227,n23566,n27249,n27253 );
   nand U27167 ( n27249,n27254,n27255,n25116,n27256 );
   nor U27168 ( n27256,n27257,n25266,n27258 );
   not U27169 ( n27258,n26170 );
   nand U27170 ( n26170,n25814,n25787 );
   nor U27171 ( n25266,n26171,n25809 );
   nor U27172 ( n27257,n27259,n25787 );
   nor U27173 ( n27259,n24348,n25104 );
   not U27174 ( n24348,n24400 );
   nor U27175 ( n25116,n24517,n24523 );
   not U27176 ( n24523,n24401 );
   nand U27177 ( n24401,n25805,n23987 );
   not U27178 ( n24517,n24394 );
   nand U27179 ( n27255,n23990,n25012 );
   not U27180 ( n25012,n24395 );
   nand U27181 ( n27254,n27260,n25806 );
   nand U27182 ( n27252,n26789,n27261 );
   nand U27183 ( n27261,n26790,n26788 );
   not U27184 ( n26789,n27262 );
   nand U27185 ( n27251,n26790,n26788,n27262 );
   nand U27186 ( n27262,n27263,n27264 );
   nand U27187 ( n27264,n27265,n27266 );
   or U27188 ( n27266,n26267,n26266 );
   not U27189 ( n27265,n26268 );
   nand U27190 ( n26268,n27267,n27268 );
   nand U27191 ( n27268,n26428,n27269 );
   nand U27192 ( n27269,n27270,n26429 );
   xor U27193 ( n26428,n26652,n27271 );
   nand U27194 ( n27271,n27272,n27273 );
   nand U27195 ( n27273,n26547,n24412 );
   nand U27196 ( n27272,n26542,n23450 );
   or U27197 ( n27267,n26429,n27270 );
   not U27198 ( n27270,n26430 );
   nand U27199 ( n26430,n27274,n27275 );
   nand U27200 ( n27275,n27276,n26391 );
   nand U27201 ( n26391,n27277,n26594 );
   nand U27202 ( n26594,n27278,n27279 );
   not U27203 ( n27279,n27280 );
   xor U27204 ( n27278,n26652,n27281 );
   nand U27205 ( n27277,n26596,n26593 );
   nand U27206 ( n26593,n27282,n27280 );
   nand U27207 ( n27280,n27283,n27284 );
   nand U27208 ( n27284,n26542,n23934 );
   nand U27209 ( n27283,n26543,n23456 );
   xor U27210 ( n27282,n27281,n26364 );
   nand U27211 ( n27281,n27285,n27286 );
   nand U27212 ( n27286,n26547,n23934 );
   nand U27213 ( n23934,n27287,n27288,n27289 );
   nand U27214 ( n27289,n26140,p2_datao_reg_3_ );
   nand U27215 ( n27288,n26136,n20645 );
   xor U27216 ( n20645,n27290,n27291 );
   and U27217 ( n27290,n27292,n27293 );
   nand U27218 ( n27287,n25696,n25265 );
   not U27219 ( n25696,n25715 );
   nand U27220 ( n25715,n27294,n27295 );
   or U27221 ( n27295,p1_ir_reg_31_,p1_ir_reg_3_ );
   or U27222 ( n27294,n24061,n24254 );
   xor U27223 ( n24061,p1_ir_reg_3_,n24056 );
   nand U27224 ( n27285,n26542,n23456 );
   nand U27225 ( n23456,n27296,n27297,n27298,n27299 );
   nand U27226 ( n27299,p1_reg0_reg_3_,n26178 );
   nand U27227 ( n27298,p1_reg1_reg_3_,n26179 );
   nand U27228 ( n27297,p1_reg2_reg_3_,n26177 );
   nand U27229 ( n27296,n26563,n26589 );
   and U27230 ( n26596,n26294,n27300 );
   nand U27231 ( n27300,n26292,n26293 );
   or U27232 ( n26293,n26297,n26296 );
   not U27233 ( n26292,n26595 );
   nand U27234 ( n26595,n27301,n27302 );
   nand U27235 ( n27302,n26502,n27303 );
   nand U27236 ( n27303,n26503,n26504 );
   xor U27237 ( n26502,n26652,n27304 );
   nand U27238 ( n27304,n27305,n27306 );
   nand U27239 ( n27306,n26547,n24296 );
   nand U27240 ( n27305,n26542,n23462 );
   or U27241 ( n27301,n26504,n26503 );
   nand U27242 ( n26503,n27307,n27308 );
   nand U27243 ( n27308,n27309,n26364 );
   nand U27244 ( n27309,n26362,n26365 );
   or U27245 ( n27307,n26362,n26365 );
   and U27246 ( n26365,n27310,n27311,n27312 );
   nand U27247 ( n27312,p1_ir_reg_0_,n25790 );
   nand U27248 ( n27311,n26543,n23465 );
   nand U27249 ( n27310,n26542,n23974 );
   xor U27250 ( n26362,n26652,n27313 );
   nand U27251 ( n27313,n27314,n27315,n27316 );
   nand U27252 ( n27316,p1_reg1_reg_0_,n25790 );
   nand U27253 ( n27315,n26542,n23465 );
   nand U27254 ( n23465,n27317,n27318,n27319,n27320 );
   nand U27255 ( n27320,p1_reg0_reg_0_,n26178 );
   nand U27256 ( n27319,p1_reg1_reg_0_,n26179 );
   nand U27257 ( n27318,p1_reg2_reg_0_,n26177 );
   nand U27258 ( n27317,p1_reg3_reg_0_,n26563 );
   nand U27259 ( n27314,n26547,n23974 );
   nand U27260 ( n23974,n27321,n27322,n27323 );
   nand U27261 ( n27323,p1_ir_reg_0_,n25265 );
   nand U27262 ( n27322,n26136,n20618 );
   and U27263 ( n20618,n27324,n27325 );
   nand U27264 ( n27324,n27326,n27327 );
   nand U27265 ( n27321,n26140,p2_datao_reg_0_ );
   nand U27266 ( n26504,n27328,n27329 );
   nand U27267 ( n27329,n26543,n23462 );
   nand U27268 ( n23462,n27330,n27331,n27332,n27333 );
   nand U27269 ( n27333,p1_reg0_reg_1_,n26178 );
   nand U27270 ( n27332,p1_reg1_reg_1_,n26179 );
   nand U27271 ( n27331,p1_reg2_reg_1_,n26177 );
   nand U27272 ( n27330,p1_reg3_reg_1_,n26563 );
   nand U27273 ( n27328,n26542,n24296 );
   nand U27274 ( n24296,n27334,n27335,n27336 );
   nand U27275 ( n27336,n26140,p2_datao_reg_1_ );
   nand U27276 ( n27335,n25761,n25265 );
   and U27277 ( n25761,n27337,n27338 );
   nand U27278 ( n27338,n27339,n24254 );
   or U27279 ( n27337,n24050,n24254 );
   xor U27280 ( n24050,n25746,n27339 );
   nand U27281 ( n27334,n26136,n20628 );
   nand U27282 ( n20628,n27340,n27341,n27342 );
   nand U27283 ( n27342,n27343,n27344 );
   nand U27284 ( n27341,n27345,n27325,si_1_ );
   nand U27285 ( n27340,n27346,n27347 );
   xor U27286 ( n27346,n27325,n27345 );
   nand U27287 ( n26294,n26296,n26297 );
   nand U27288 ( n26297,n27348,n27349 );
   nand U27289 ( n27349,n26542,n24321 );
   nand U27290 ( n27348,n26543,n23459 );
   xor U27291 ( n26296,n26364,n27350 );
   nand U27292 ( n27350,n27351,n27352 );
   nand U27293 ( n27352,n26547,n24321 );
   nand U27294 ( n24321,n27353,n27354,n27355 );
   nand U27295 ( n27355,n26140,p2_datao_reg_2_ );
   nand U27296 ( n27354,n26136,n20635 );
   xor U27297 ( n20635,n27356,n27357 );
   and U27298 ( n27356,n27358,n27359 );
   nand U27299 ( n27353,n25730,n25265 );
   not U27300 ( n25730,n25726 );
   nand U27301 ( n25726,n27360,n27361 );
   or U27302 ( n27361,p1_ir_reg_2_,p1_ir_reg_31_ );
   nand U27303 ( n27360,p1_ir_reg_31_,n27362 );
   nand U27304 ( n27362,n24055,n24056 );
   nand U27305 ( n24055,p1_ir_reg_2_,n27363 );
   nand U27306 ( n27363,n25746,n27339 );
   not U27307 ( n27339,p1_ir_reg_1_ );
   not U27308 ( n25746,p1_ir_reg_0_ );
   nand U27309 ( n27351,n26542,n23459 );
   nand U27310 ( n23459,n27364,n27365,n27366,n27367 );
   nand U27311 ( n27367,p1_reg0_reg_2_,n26178 );
   nand U27312 ( n27366,p1_reg1_reg_2_,n26179 );
   nand U27313 ( n27365,p1_reg2_reg_2_,n26177 );
   nand U27314 ( n27364,p1_reg3_reg_2_,n26563 );
   nand U27315 ( n27276,n26389,n26390 );
   or U27316 ( n27274,n26390,n26389 );
   xor U27317 ( n26389,n27368,n26652 );
   nor U27318 ( n27368,n27369,n27370 );
   nor U27319 ( n27370,n23933,n27371 );
   not U27320 ( n23933,n23453 );
   nor U27321 ( n27369,n23919,n27372 );
   not U27322 ( n23919,n24372 );
   nand U27323 ( n26390,n27373,n27374 );
   nand U27324 ( n27374,n26542,n24372 );
   nand U27325 ( n24372,n27375,n27376,n27377 );
   nand U27326 ( n27377,n26140,p2_datao_reg_4_ );
   nand U27327 ( n27376,n25681,n25265 );
   and U27328 ( n25681,n27378,n27379 );
   or U27329 ( n27379,p1_ir_reg_31_,p1_ir_reg_4_ );
   nand U27330 ( n27378,p1_ir_reg_31_,n27380 );
   nand U27331 ( n27380,n24067,n24066 );
   nand U27332 ( n24066,p1_ir_reg_4_,n27381 );
   nand U27333 ( n27375,n26136,n20652 );
   xor U27334 ( n20652,n27382,n27383 );
   and U27335 ( n27382,n27384,n27385 );
   nand U27336 ( n27373,n26543,n23453 );
   nand U27337 ( n23453,n27386,n27387,n27388,n27389 );
   nand U27338 ( n27389,n26386,n26563 );
   not U27339 ( n26386,n24368 );
   nand U27340 ( n24368,n27390,n27391 );
   nand U27341 ( n27390,n26385,n26589 );
   not U27342 ( n26589,p1_reg3_reg_3_ );
   not U27343 ( n26385,p1_reg3_reg_4_ );
   nand U27344 ( n27388,p1_reg0_reg_4_,n26178 );
   nand U27345 ( n27387,p1_reg1_reg_4_,n26179 );
   nand U27346 ( n27386,p1_reg2_reg_4_,n26177 );
   nand U27347 ( n26429,n27392,n27393 );
   nand U27348 ( n27393,n26542,n24412 );
   nand U27349 ( n24412,n27394,n27395,n27396 );
   nand U27350 ( n27396,n26140,p2_datao_reg_5_ );
   nand U27351 ( n27395,n26136,n20661 );
   xor U27352 ( n20661,n27397,n27398 );
   and U27353 ( n27397,n27399,n27400 );
   nand U27354 ( n27394,n25265,n25631 );
   not U27355 ( n25631,n25630 );
   xor U27356 ( n25630,p1_ir_reg_5_,n27401 );
   nand U27357 ( n27401,p1_ir_reg_31_,n24067 );
   nand U27358 ( n27392,n26543,n23450 );
   nand U27359 ( n23450,n27402,n27403,n27404,n27405 );
   nand U27360 ( n27405,n26563,n24385 );
   xor U27361 ( n24385,n26425,n27391 );
   not U27362 ( n26425,p1_reg3_reg_5_ );
   nand U27363 ( n27404,p1_reg0_reg_5_,n26178 );
   nand U27364 ( n27403,p1_reg1_reg_5_,n26179 );
   nand U27365 ( n27402,p1_reg2_reg_5_,n26177 );
   nand U27366 ( n27263,n26266,n26267 );
   nand U27367 ( n26267,n27406,n27407 );
   nand U27368 ( n27407,n26542,n24446 );
   nand U27369 ( n27406,n26543,n23447 );
   xor U27370 ( n26266,n27408,n26652 );
   nor U27371 ( n27408,n27409,n27410 );
   nor U27372 ( n27410,n24471,n27371 );
   not U27373 ( n27371,n26542 );
   not U27374 ( n24471,n23447 );
   nand U27375 ( n23447,n27411,n27412,n27413,n27414 );
   nand U27376 ( n27414,p1_reg0_reg_6_,n26178 );
   nand U27377 ( n27413,p1_reg1_reg_6_,n26179 );
   nand U27378 ( n27412,p1_reg2_reg_6_,n26177 );
   nand U27379 ( n27411,n26263,n26563 );
   not U27380 ( n26263,n24425 );
   nand U27381 ( n24425,n27415,n27242 );
   nand U27382 ( n27415,n26262,n27416 );
   nand U27383 ( n27416,p1_reg3_reg_5_,n27417 );
   not U27384 ( n26262,p1_reg3_reg_6_ );
   nor U27385 ( n27409,n23897,n27372 );
   not U27386 ( n27372,n26547 );
   not U27387 ( n23897,n24446 );
   nand U27388 ( n24446,n27418,n27419,n27420 );
   nand U27389 ( n27420,n26140,p2_datao_reg_6_ );
   nand U27390 ( n27419,n25618,n25265 );
   not U27391 ( n25618,n25635 );
   nand U27392 ( n25635,n27421,n27422 );
   or U27393 ( n27422,p1_ir_reg_31_,p1_ir_reg_6_ );
   nand U27394 ( n27421,p1_ir_reg_31_,n27423 );
   nand U27395 ( n27423,n24081,n24082 );
   nand U27396 ( n24081,p1_ir_reg_6_,n27424 );
   nand U27397 ( n27424,n24075,n24076 );
   not U27398 ( n24076,p1_ir_reg_5_ );
   nand U27399 ( n27418,n26136,n20668 );
   xor U27400 ( n20668,n27425,n27426 );
   xor U27401 ( n27425,n27427,si_6_ );
   nand U27402 ( n26788,n27428,n27429 );
   not U27403 ( n27429,n27430 );
   xor U27404 ( n27428,n26652,n27431 );
   nand U27405 ( n26790,n27432,n27430 );
   nand U27406 ( n27430,n27433,n27434 );
   nand U27407 ( n27434,n26543,n23444 );
   nand U27408 ( n27433,n26542,n24482 );
   xor U27409 ( n27432,n27431,n26364 );
   nand U27410 ( n27438,n25809,n25806 );
   nand U27411 ( n27431,n27439,n27440 );
   nand U27412 ( n27440,n26542,n23444 );
   nand U27413 ( n23444,n27441,n27442,n27443,n27444 );
   nand U27414 ( n27444,n26563,n24459 );
   xor U27415 ( n24459,n27243,n27242 );
   nand U27416 ( n27242,p1_reg3_reg_5_,n27417,p1_reg3_reg_6_ );
   not U27417 ( n27417,n27391 );
   nand U27418 ( n27391,p1_reg3_reg_4_,p1_reg3_reg_3_ );
   not U27419 ( n27243,p1_reg3_reg_7_ );
   nand U27420 ( n27443,p1_reg0_reg_7_,n26178 );
   not U27421 ( n27445,n27447 );
   nand U27422 ( n27442,p1_reg1_reg_7_,n26179 );
   nand U27423 ( n27441,p1_reg2_reg_7_,n26177 );
   xor U27424 ( n27446,n24254,n24249 );
   not U27425 ( n24249,p1_ir_reg_30_ );
   xor U27426 ( n27447,p1_ir_reg_31_,n24240 );
   not U27427 ( n24240,p1_ir_reg_29_ );
   nor U27428 ( n25783,n25805,n25104 );
   not U27429 ( n25104,n25802 );
   nand U27430 ( n25802,n23979,n25806,n23989 );
   nor U27431 ( n25805,n23984,n23990 );
   nand U27432 ( n27439,n26547,n24482 );
   nand U27433 ( n27436,n23990,n27448,n23987 );
   nand U27434 ( n27435,n27449,n27448 );
   nand U27435 ( n27449,n24403,n27450,n26187 );
   nor U27436 ( n26187,n25814,n26133 );
   not U27437 ( n26133,n25807 );
   nand U27438 ( n25807,n25291,n25809 );
   not U27439 ( n27450,n25785 );
   nor U27440 ( n25785,n23984,n23987 );
   nand U27441 ( n23984,n23989,n25291 );
   nand U27442 ( n24403,n26188,n25806 );
   not U27443 ( n25806,n23990 );
   nand U27444 ( n27227,n26225,n24482 );
   nand U27445 ( n24482,n27451,n27452,n27453 );
   nand U27446 ( n27453,n26140,p2_datao_reg_7_ );
   nand U27447 ( n27452,n25265,n25574 );
   not U27448 ( n25574,n25573 );
   xor U27449 ( n25573,p1_ir_reg_7_,n27454 );
   nand U27450 ( n27454,p1_ir_reg_31_,n24082 );
   nand U27451 ( n27451,n26136,n20677 );
   xor U27452 ( n20677,n27455,n26807 );
   nand U27453 ( n26807,n27456,n27457 );
   nand U27454 ( n27457,si_6_,n27458 );
   nand U27455 ( n27458,n27427,n27426 );
   or U27456 ( n27456,n27426,n27427 );
   and U27457 ( n27427,n27400,n27459 );
   nand U27458 ( n27459,n27398,n27399 );
   nand U27459 ( n27399,n27460,n27461,n27462 );
   not U27460 ( n27462,si_5_ );
   nand U27461 ( n27461,n16572,p1_datao_reg_5_ );
   nand U27462 ( n27460,n16576,p2_datao_reg_5_ );
   nand U27463 ( n27398,n27384,n27463 );
   nand U27464 ( n27463,n27383,n27385 );
   or U27465 ( n27385,n27464,si_4_ );
   nand U27466 ( n27383,n27292,n27465 );
   nand U27467 ( n27465,n27291,n27293 );
   nand U27468 ( n27293,n27466,n27467,n27468 );
   not U27469 ( n27468,si_3_ );
   nand U27470 ( n27467,n16572,p1_datao_reg_3_ );
   nand U27471 ( n27466,n16576,p2_datao_reg_3_ );
   nand U27472 ( n27291,n27358,n27469 );
   nand U27473 ( n27469,n27359,n27357 );
   nand U27474 ( n27357,n27470,n27471,n27472 );
   nand U27475 ( n27472,n27344,si_1_ );
   not U27476 ( n27471,n27343 );
   nor U27477 ( n27343,n27345,n27347 );
   not U27478 ( n27347,si_1_ );
   or U27479 ( n27470,n27325,n27345 );
   nand U27480 ( n27345,n27473,n27474 );
   nand U27481 ( n27474,n16576,n19468 );
   not U27482 ( n19468,p2_datao_reg_1_ );
   nand U27483 ( n27473,n16572,n19469 );
   not U27484 ( n19469,p1_datao_reg_1_ );
   not U27485 ( n27325,n27344 );
   nor U27486 ( n27344,n27327,n27326 );
   and U27487 ( n27326,n27475,n27476 );
   nand U27488 ( n27476,n16572,p1_datao_reg_0_ );
   nand U27489 ( n27475,n16576,p2_datao_reg_0_ );
   not U27490 ( n27327,si_0_ );
   nand U27491 ( n27359,n27477,n27478 );
   or U27492 ( n27358,n27477,n27478 );
   not U27493 ( n27478,si_2_ );
   nand U27494 ( n27477,n27479,n27480 );
   or U27495 ( n27480,n16572,p2_datao_reg_2_ );
   nand U27496 ( n27479,n16572,n19464 );
   not U27497 ( n19464,p1_datao_reg_2_ );
   nand U27498 ( n27292,n27481,n27482,si_3_ );
   nand U27499 ( n27482,n16576,n19358 );
   not U27500 ( n19358,p2_datao_reg_3_ );
   nand U27501 ( n27481,n16572,n19357 );
   not U27502 ( n19357,p1_datao_reg_3_ );
   nand U27503 ( n27384,si_4_,n27464 );
   nand U27504 ( n27464,n27483,n27484 );
   nand U27505 ( n27484,n16572,p1_datao_reg_4_ );
   nand U27506 ( n27483,n16576,p2_datao_reg_4_ );
   nand U27507 ( n27400,n27485,n27486,si_5_ );
   nand U27508 ( n27486,n16576,n19329 );
   not U27509 ( n19329,p2_datao_reg_5_ );
   nand U27510 ( n27485,n16572,n19331 );
   not U27511 ( n19331,p1_datao_reg_5_ );
   nand U27512 ( n27426,n27487,n27488 );
   nand U27513 ( n27488,n16576,n19325 );
   not U27514 ( n19325,p2_datao_reg_6_ );
   or U27515 ( n27487,n16576,p1_datao_reg_6_ );
   nor U27516 ( n27455,n27160,n27166 );
   nor U27517 ( n27166,n27489,si_7_ );
   not U27518 ( n27160,n26805 );
   nand U27519 ( n26805,si_7_,n27489 );
   nand U27520 ( n27489,n27490,n27491 );
   nand U27521 ( n27491,n16572,p1_datao_reg_7_ );
   nand U27522 ( n27490,n16576,p2_datao_reg_7_ );
   nand U27523 ( n27494,p1_addr_reg_19_,n14939,p2_addr_reg_19_,n17703 );
   not U27524 ( n14939,p2_rd_reg );
   or U27525 ( n27493,p1_rd_reg,p2_addr_reg_19_,p1_addr_reg_19_,n17703 );
   not U27526 ( n17703,p3_addr_reg_19_ );
   nand U27527 ( n26298,n23566,n27495 );
   nand U27528 ( n27495,n25269,n27496 );
   nand U27529 ( n27496,n27253,n25267 );
   nand U27530 ( n25267,n27497,n23976 );
   nand U27531 ( n23976,n27498,n25809 );
   not U27532 ( n27498,n26171 );
   nand U27533 ( n26171,n25291,n23990,n23987 );
   nand U27534 ( n27497,n27260,n23990 );
   not U27535 ( n27260,n26127 );
   nand U27536 ( n26127,n26188,n23987 );
   nor U27537 ( n26188,n25291,n23989 );
   not U27538 ( n23989,n25809 );
   not U27539 ( n25291,n23979 );
   not U27540 ( n27253,n27233 );
   nand U27541 ( n27233,n23565,n23983,n25271 );
   not U27542 ( n25271,n23982 );
   nand U27543 ( n23982,n23995,n27499 );
   or U27544 ( n27499,n24265,p1_d_reg_1_ );
   nand U27545 ( n23995,n27500,n27501 );
   and U27546 ( n23983,n27502,n27503,n27504,n27505 );
   nor U27547 ( n27505,n27506,n27507,n27508,n27509 );
   nor U27548 ( n27509,n24265,n24256 );
   not U27549 ( n24256,p1_d_reg_6_ );
   nor U27550 ( n27508,n24265,n24258 );
   not U27551 ( n24258,p1_d_reg_13_ );
   nor U27552 ( n27507,n24265,n24260 );
   not U27553 ( n24260,p1_d_reg_17_ );
   nor U27554 ( n27506,n27510,n24265 );
   nor U27555 ( n27510,p1_d_reg_22_,p1_d_reg_24_,p1_d_reg_23_ );
   nor U27556 ( n27504,n27511,n27512,n27513,n27514 );
   nor U27557 ( n27514,n24265,n24262 );
   not U27558 ( n24262,p1_d_reg_19_ );
   nor U27559 ( n27513,n24265,n24259 );
   not U27560 ( n24259,p1_d_reg_16_ );
   nor U27561 ( n27512,n27515,n24265 );
   nor U27562 ( n27515,p1_d_reg_7_,p1_d_reg_9_,p1_d_reg_8_ );
   nor U27563 ( n27511,n24265,n24257 );
   not U27564 ( n24257,p1_d_reg_10_ );
   nor U27565 ( n27503,n27516,n27517,n27518,n27519 );
   nor U27566 ( n27519,n24265,n24264 );
   not U27567 ( n24264,p1_d_reg_29_ );
   nor U27568 ( n27518,n24265,n24255 );
   not U27569 ( n24255,p1_d_reg_2_ );
   nor U27570 ( n27517,n24265,n24263 );
   not U27571 ( n24263,p1_d_reg_27_ );
   nor U27572 ( n27516,n24265,n24261 );
   not U27573 ( n24261,p1_d_reg_18_ );
   nor U27574 ( n27502,n27520,n27521,n27522,n27523 );
   nor U27575 ( n27523,n27524,n24265 );
   nor U27576 ( n27524,p1_d_reg_5_,p1_d_reg_4_,p1_d_reg_3_,p1_d_reg_30_ );
   nor U27577 ( n27522,n27525,n24265 );
   nor U27578 ( n27525,p1_d_reg_20_,p1_d_reg_26_,p1_d_reg_25_ );
   nor U27579 ( n27521,n27526,n24265 );
   nor U27580 ( n27526,p1_d_reg_15_,p1_d_reg_14_,p1_d_reg_12_,p1_d_reg_11_ );
   nor U27581 ( n27520,n27527,n24265 );
   nor U27582 ( n27527,p1_d_reg_21_,p1_d_reg_31_,p1_d_reg_28_ );
   not U27583 ( n23565,n23980 );
   nand U27584 ( n23980,n23998,n27528 );
   or U27585 ( n27528,n24265,p1_d_reg_0_ );
   nand U27586 ( n27530,n27532,n25263 );
   not U27587 ( n25263,p1_b_reg );
   nand U27588 ( n27529,n27533,n27501,p1_b_reg );
   nand U27589 ( n23998,n27500,n27533 );
   nand U27590 ( n25269,n25814,n23978 );
   nor U27591 ( n23978,n25787,n25809 );
   nand U27592 ( n25809,n27534,n27535 );
   nand U27593 ( n27535,p1_ir_reg_20_,n24254 );
   nand U27594 ( n27534,n24175,n24176,p1_ir_reg_31_ );
   nand U27595 ( n24175,p1_ir_reg_20_,n24170 );
   not U27596 ( n25814,n27437 );
   nand U27597 ( n27437,n23990,n23979 );
   nand U27598 ( n23979,n27536,n27537 );
   nand U27599 ( n27537,p1_ir_reg_19_,n24254 );
   nand U27600 ( n27536,n24169,n24170,p1_ir_reg_31_ );
   nand U27601 ( n24169,p1_ir_reg_19_,n26947 );
   and U27602 ( n23566,n27448,p1_state_reg,n25791 );
   not U27603 ( n27448,n25790 );
   not U27604 ( p1_u3086,p1_state_reg );
   not U27605 ( p1_u3085,n25789 );
   nand U27606 ( n25789,n27538,n23371 );
   nor U27607 ( n25790,n27501,n27533,n27500 );
   not U27608 ( n27500,n27531 );
   nand U27609 ( n27531,n27539,n27540 );
   nand U27610 ( n27540,p1_ir_reg_26_,n24254 );
   nand U27611 ( n27539,n24217,n24218,p1_ir_reg_31_ );
   nand U27612 ( n24217,p1_ir_reg_26_,n27541 );
   nand U27613 ( n27541,n24211,n24212 );
   not U27614 ( n27533,n27532 );
   nand U27615 ( n27532,n27542,n27543 );
   nand U27616 ( n27543,p1_ir_reg_24_,n24254 );
   nand U27617 ( n27542,n24203,n24204,p1_ir_reg_31_ );
   nand U27618 ( n24203,p1_ir_reg_24_,n27544 );
   nand U27619 ( n27544,n24197,n24198 );
   not U27620 ( n24198,p1_ir_reg_23_ );
   xor U27621 ( n27501,n27545,n24212 );
   not U27622 ( n24212,p1_ir_reg_25_ );
   nor U27623 ( n27545,n24211,n24254 );
   nand U27624 ( n27538,n27546,p1_state_reg );
   nand U27625 ( n27546,n27547,n27492 );
   nand U27626 ( n27492,n25743,n25264 );
   not U27627 ( n25264,n25106 );
   nand U27628 ( n25106,n27548,n27549 );
   nand U27629 ( n27549,p1_ir_reg_28_,n24254 );
   nand U27630 ( n27548,n24231,n24232,p1_ir_reg_31_ );
   not U27631 ( n24232,n24239 );
   nor U27632 ( n24239,p1_ir_reg_27_,p1_ir_reg_28_,n24218 );
   nand U27633 ( n24231,p1_ir_reg_28_,n27550 );
   nand U27634 ( n27550,n24225,n24226 );
   not U27635 ( n24226,p1_ir_reg_27_ );
   xor U27636 ( n25743,p1_ir_reg_27_,n27551 );
   nand U27637 ( n27551,p1_ir_reg_31_,n24218 );
   not U27638 ( n24218,n24225 );
   nor U27639 ( n24225,p1_ir_reg_25_,p1_ir_reg_26_,n24204 );
   not U27640 ( n24204,n24211 );
   nor U27641 ( n24211,p1_ir_reg_23_,p1_ir_reg_24_,n24190 );
   nand U27642 ( n27547,n25105,n25791 );
   xor U27643 ( n25791,p1_ir_reg_23_,n27552 );
   nand U27644 ( n27552,p1_ir_reg_31_,n24190 );
   nor U27645 ( n25105,n23987,n23990 );
   xor U27646 ( n23990,n27553,n24184 );
   nor U27647 ( n27553,n24183,n24254 );
   not U27648 ( n23987,n25787 );
   nand U27649 ( n25787,n27554,n27555 );
   nand U27650 ( n27555,p1_ir_reg_22_,n24254 );
   nand U27651 ( n27554,n24189,n24190,p1_ir_reg_31_ );
   not U27652 ( n24190,n24197 );
   nor U27653 ( n24197,p1_ir_reg_21_,p1_ir_reg_22_,n24176 );
   not U27654 ( n24176,n24183 );
   nand U27655 ( n24189,p1_ir_reg_22_,n27556 );
   nand U27656 ( n27556,n24183,n24184 );
   not U27657 ( n24184,p1_ir_reg_21_ );
   nor U27658 ( n24183,n24170,p1_ir_reg_20_ );
   or U27659 ( n24170,n26947,p1_ir_reg_19_ );
   nand U27660 ( n26947,n24162,n24164 );
   not U27661 ( n24164,p1_ir_reg_18_ );
   not U27662 ( n24162,n24163 );
   nand U27663 ( n24163,n24154,n24155 );
   not U27664 ( n24155,p1_ir_reg_17_ );
   nor U27665 ( n24154,p1_ir_reg_15_,p1_ir_reg_16_,n24140 );
   not U27666 ( n24140,n24139 );
   nor U27667 ( n24139,n26750,p1_ir_reg_14_ );
   nand U27668 ( n26750,n24125,n24126 );
   not U27669 ( n24126,p1_ir_reg_13_ );
   nor U27670 ( n24125,p1_ir_reg_11_,p1_ir_reg_12_,n26843 );
   not U27671 ( n26843,n26879 );
   nor U27672 ( n26879,p1_ir_reg_10_,p1_ir_reg_9_,n24096 );
   not U27673 ( n24096,n26846 );
   nor U27674 ( n26846,p1_ir_reg_7_,p1_ir_reg_8_,n24082 );
   not U27675 ( n24082,n24089 );
   nor U27676 ( n24089,p1_ir_reg_5_,p1_ir_reg_6_,n24067 );
   not U27677 ( n24067,n24075 );
   nor U27678 ( n24075,n27381,p1_ir_reg_4_ );
   or U27679 ( n27381,n24056,p1_ir_reg_3_ );
   or U27680 ( n24056,p1_ir_reg_1_,p1_ir_reg_2_,p1_ir_reg_0_ );
endmodule
